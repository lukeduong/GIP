PK   �EX�&:  �n    cirkitFile.json�}]s丱�_q辊
$ ~��}wᇻ�Xoxf&*��Ql�ԫV{의�~VU��H�ʓ�x�t�G�&HH�|���}x�u�O�������Ǉ������<�?5�5�7��vϏ��=5�~���s�={��!k���oC�]Q�vh\����3o�1��3یm�*W������|���~���Ǉ��yW�ei�ό]��eU��,o�</���~go��}��i����HB�	铘�=�����){j�?���>=~l����=>�?�K���mF2�y�m�;��iȬu}A�	�w�����������yq�O��Ed�.OX�s*��ʪP0�YETe�<�l_UT�'�Y"��BB_�
��~)D 1��U	�����̍��|Q�Yc}��a���]o�A�*1�ZB_�D��[Ku�,��H�~9�1� �>��g&ioHr��"գ�P��tU��3_U>�ﲮ�Zk�ޔ��HޥR�OM5�z}jg�б�]֚���j(��{�:qC��.|�TW�z qK�����Y Ur���$���E�Cd�Q,h�����!�$I��C��������CR�'9D`!Uj�CR�%9D`!�L�Cr�CR�#9D`!�N1��9�v�!�v�!�v�!�v�!�v�!�v�!�v�!�v�!�v�!�v�!��˵SXȵSXȵSXȵSXȵSXȵSXȵSXȵSXȵSXȵSav�\;���\;���\;���\;���\;���\;���\;���\;���\;���\;�fWȵSXȵSXȵs!^'q:���E02q����h�l089; ��߸p��f��{5#bBs���o�"��V�I������>͟Mf*�i+�uiR�r���b����&08��7�Z�&Ӕ3&�7�b"mc3���o,Ǫ[��ˡ��.�尶+����#,;�+9J�Z''U���,&N�3���o��z{��v(;²3�k�k;(;²�ˀ��#p���G`~q2�~������/.�fuU=c-���8�r���P��ЂUpx�����O��c���	M�x�� ��Ȱ��j{�ఖ\K��4��^ME:8�[�yk�h��� ����`�A��#0��7l?p���G`~qk�~� ˏ����wp���G`~q;�~�0ˏ���F"���	���_��4� 0?󋛷��G=X~��������G`~q��~��ˏ���V?��������M�`���,?��+���X~�7�b��������-�`���,?�q���X~�����?���/n��`��_ܺ�8���#0���l?p���G`~q�<�~��ˏ���F��������`���,?�������ˏ��bZ�������ń`���,?�8���X~������?���/�?�`��_L��8���#0��rl?p���G`~1Y�~��ˏ��b���������EX����ˏ��bj%�������ŤP`���,?�����X~�q���?���/���
 � ���#�X~�Ӷ���?���/&��`��_L��8���#0���k�`��_LO�8���#0��Xl?p���G+�6f%�̮���eZ̍�/�Yn�~��wsn8ٙ�q��I�cry��s\ey	�����Nr�˜��_&��ڐ�1���)dx�JB@��T���I�CR�#�Icp�H3ѫ�
�0��m"u#���zf���۾�:��m`໡��.o��ý�J�ʠ�U=-U���A�zz���~��c��\��_&��X�2�����.�U=�E��F�vB��h�����f��n�/���a�[��ov
���B�������T���7;�tk}�����Z_���8�����̭���f�Nn�/�x��7;�qk}���NF�Z_�������������7;uosbyY��9��I�̼��Ic,&�(����o�Kn��V��������U=-$��i�yZGx�����8�W?ݏ1��/'�t���&�nnK>�`[d�j|\��!����F��0�S��)R��;[ɝ�r�4��;[؛�2��y
�nRj�u�\zw��H?oT��K?oԩ9;�p�N����wN�S��L��2#��Mܙ��y��eY��ecS��o�>�G�d��we.����.�����r�c�^��)�a�Y��RNú3�^]�a=��I�Yw�/)�g�]ڿP*"b�]��P��=S<`��7�>,=���.�sJ,�'�s�W͍w��+��ɼ�1k��e�m�f������?V�t�ƪ��X�ӱ�zz
�U==k����5`UO����gX�ӳ<���������=���?^}��]��ǫ/��+_�x���w����T���w�������|����ߕ���B������q	����?^}i�+��+_�x�'��e�=?�Ǐ�O7~����+����V]=�F_[�hd��i�d�ƺ�1"#����/cdQ�\�Ǧ����C1�h��{�	��3�#PQ�޵2F9�F��F�o��Q�bTb�g�P�V��Q�bTOom�j)����ֶ}W�B�&�jOj[�޷$��m�-�������Ǳ�BN0�Is���?y�|/�-��L�� �}[BN0'�������T����>Sq�/����c8����8���0G!�i.�	����C2Ӝ	�L�-H}	�d��'��[���LsP N0w0G!�i��	����($3��8�t��t�d��G'��;����̴C�	����($3�� q�鸇�8
�L;N@�`:�a:�B��a�ps�0G!���0N0�0G!��0N0�0G!�L�0N0�a:�B��a�`:��t�3��8�t<��8
)f��q��x�qR̤
�����(����	��L�QH13%�L������oƸLX���C�:��Dp��`T�Y�/�]/ә.-w�n�9W�]�\v�Lp
G�U�+-pEX�����^����+®s��^Ȁ����ι"�:犰��ApT`����T��1��]/�q�X@�+�p�e� �����sE�u�a���@��J*\��� 8*Ю\I�k\�bX҉�Tؒ۸�YǶ��%��ߨ�V'�Z`��N�E�<O>ʶ:��[�4��sX�&�`*l�9xP�0�l ~��-���V'#�HL�-鰍{1tl��[�a����V'"SaK:l����De*lI�m���aA'.SaK:l�^%���e*lI�m�s�c[�H�tؒ۸wLǶ��%�q��mu�2���6��ӱ���1���6�IԱ�N\�t�ƽ�:�Չ�Tؒ۸GTǶ:q�
[�a����V'.SaK:l�]�:��L�-鰍{�ul����%�q��mu�2���6�ױ�N\�t��=�:�Չ�Tؒ۸7_Ƕ:q�
[�as��V'.SaK:lc����e*lI�m���c[��L�-鰍�+tl����%�1��m�N\�t��\":�Չ�TؒۘEǶ:q�
[�as���V'.SaK:lc����e*lI�m̵�c[��L�-鰍9�tl����%�1���mu�2���6�pұ�N\�t��\T:�Չ�TؒۘSKŶ�N\�t���`:�Չ�Tؒۘ�LǶ:q�
[�as���V'.SaK:lc�9���e*lI�m̝�c[�,Ji>t�\'.�u�2���6�2Ա�N\�t�Ɯ�:�Չ�Tؒۘ[RǶ:q�
[�asd�ضЉ�Tؒۘ�SǶ:q�
[�as���V'.SaK<�/�D7m3�i��[o3�QD�!����&��N�ü%��v#J"��F�D�(�s�7�L���Y#6�Α�<,y#ʔ�z~�F�D�(���[�伫�kB#lz����y��gu�]��]kMћ�<�~�]�P�2�����Q�Z������gƌ.�C鲪�m�7C��Po[�� \&�̏�߈rP��#�_P��}�u&�� 廡��.o��ـ�֕����,�U�e��*/%q��F��)Q�
lDI��eUyY(����:��b�7u��V�����
������[a0>�:�y+ƋS� o�i0ƋS�o��xq�ޭ0/N�u��ũe���/N�ۺ4��xq�@ӭ0/N��ũ�9��`�8u�V���|��Ɯʦ
T՚���f�x�#������Z��BY}$�]�X(n?Q��	P�VYT�w� e�Q�PV�$e�I�PV[$e�A�n�A�`0޻>����v+���h�2s��P�}�X�fv��y��rXo�,��T�И(�a�x�".nuډ�2���11��B��u�{ߒ ej�m[U"�L�z�:ٝ8c��l(�!�|�N�"3U���X�F?�BY��j?�Bqk^7�jt� :[gގ]֚���j(��{ߺu��P
��P&���/�Ĕ)e��P���m�((S;���֒':||�ۢ�L�͍I)CY�}(O���c曪���6Y3�]Y��j�����:��BY��[���x��P���&��,�:������+����d�jO�BY�Y(��4e5�c���3Y(��L��8���:�d���3y^r^����3y0�]�J��`<x}*������dƋק�y0 �x��T2���S�<��O%�`0^�>���u1^�>�̃%0^�>�̃9��_&������s�<�|��w�����=_��������/f�0��@����l �@@f5C���4�0�i4a2Sd a2S�a2S�a2��#�8���6L�	&�($��0�`�M0�F!�}����o�	8
��c'��L�QHf�c8�t��t�d��	N��7n �q�q��ϙ`8�t��t�d��9N0�0G!��<�L�-L�QHf?�	�a:�`:�B2��9'�L
n*����($����p�鸃�8
����b8�t��t�d�+�1�`:�a:�B2���N0�0G!�D�0N�9qܤ8L�=L�QH1!.�L�=L�QH1+�L�=L�QH1�'��L�s����b�I'���0G!ń�0N����ϛ0�a:�B���`�`:��t���8�t���8
)&ւq��x����$Y�$lh�}.+ *�p%�f7K��F�U�+�p5�Y�54*Ю\I����b�Q�v��J*\Cܥb�Y.l�4��
�0R��,6�\I�k���u�b�����f	�Ѩ@�jp%�f7K~�F�U�+�p5�Y�k4*Ю\I�k\��D\*lI�m\۬c[��K)�҉�H'�"��K�-鰍k�ul�}��%�qͼ�mu"0���6��ױ�N�t��=:�Չ�Tؒ۸CǶ:ј
[�a����V'"SaK:l����De*lI�m���aA'.SaK:l�^%���e*lI�m�s�c[�/bJ��t�2��Y��L�-鰍{�tl����%�q/��mu�2���6�IԱ�N\�t�ƽ�:�Չ�Tؒ۸GTǶ:q�
[�a����V'.SaK:l�]��I:q�
[�a���V'.SaK:l�j���e*lI�m��c[�ՊJ�u�2��9��L�-鰍{�ul����%�1ǀ�mu�2���6�Jб�N\�t�Ɯ:�Չ�Tؒۘ�BǶ:q�
[�asp�����e*lI�m�%�c[��L�-鰍9Qtl����%�1���mu�2���6�ѱ��N2��d:q�׉˼N\�t�ƜA:�Չ�Tؒۘ�HǶ:q�
[�as8��V'.SaK:lc.*���e*lI�m̩�b�\'.SaK:lcn0���e*lI�m�q�c[��L�-鰍��tl����%�1眎mu�2���6��ӱ�R��4:qY���:q�
[�as��V'.SaK:lcNF���e*lI�m�-�c[��L�-鰍92Ul[��e*lI�m���c[��L�-鰍9Kul����%ۗ����ɴC歷��(�ҐY���Z�R��aވ��M�%�Mv#J"��F�D��(�\�Q٭7�$�QoDId�ވ������@λ�&4¦�*�L�g��|V7�e]ݵ��)����Q0\V[e�%�}Y�z�3cF���tY��6˛!ϋa(Ʀ_�e�.,�U��PV�����3Y�(�]Vwy���@�l�nʪ]X(�va�`첪�,�U�e��*/eUyY(���BYU^�ׁ�㽩㶷�`�7u��V�����
�����[a0^�:y+H�1^�:x+ƋS��n��xq�ۭ0/N�(����xq��֭0��ƋS�n��xq��Э0/Nι�ũ#0��`�8u��L7�T6U���d�6�(�S�<�l_UT��Y(���B�<�j�d���J�j�d���I�j�d���H�j��y�y1޻>������i�*ڡ���<u�5ַ�F*|���S=�����Tc��v�BYm�,��v�BY�j�1��M6�ݐyC>t'm����}k���`��wm���e�_FS��@g��۱�Z3�Xe�Vc�[�e�.,�U��P0vYmG,��v�BYmG,��vT�u�S66�����z�M�}WVႩ�ua���e�_X(����z�U�d�ј����6U3tyEu�nʪ]X(�va�`�ڎX(�툅�ڎX(�툅�:�d���3y^r^����3y0�]�J��`<x}*������dƋק�y0 �x��T2���S�<��O%�`0^�>���u1^�>�̃%0^�>�̃9��_n�����{�������q���7?�?�w�>6����v�O��t���o_�}��Ś��'�M㪦)���mx����.w�뇺̝�\g�p���o�j�j(�&�yQu�v_gm�jj}Wؒڲ+��n��CUx��:��<ڮvYmG���#���k�-�;{��eϜ��3uk�W��*���CV��e����ZCaԙ���/��}�2ܿ��"k�n����ѹ��	s��L�;1|��m�֬�q�ݢ6��&��28U�U�6��S�f,���6EЙ&�me�U�W5&�!�͏U�9��Y7E�UM^�8�#�s��YwN:;��6�s�[_4q���E*E���	N�B����`����u�������-����hIs�eT���af�d��M.��'�0Wf���0�w��U�+pET.7�H���rk���3�m���o����%�٢�����`�w{�����ء0�=�n���N|wY3�&S[ɐ�{��$o!��kd����&V�I�b69�X�n��h$�y2�`��<9�fn�y�c���5�+퀹�K�B�3/��j�����-���:D�+��\	#Yu%���9)I�u;�5b�;'&[���R��b"�+y1�kPL����d"1JP̥y�A��1��g�'�=z���t�&Y�b:���,��1%��U[f�@���M�|Rr�D��\�(�s�+f.Ӕ�9�!2��&�̴���r��1�F�0���d �1���M�kewO'������.���J����ǿ��y�V-|x�¿����o?�����~���W��W�������V`�	b�	H�cN�������`e���p����t�����p�	�c��UBo�lVN@�zVN@��6�o�����M<@L@���o��bҾAL@,͠�5tMy�&���珲ځ��b���ޥ?����+�g����
x�Q�|I�ܫ�{޳�/5�kn�>Z��w�N!g��Uq�ѻl��3Bﱐ�b��`��e+�m<�>��Bl�X`���@ $��A�{�����������w��0�zk�]���������񷟿�����5��p�o�L����Z�*��i�8{�z��}�����	�Ō�a�����u��_��~SN��LDH�[�A��*�7ڕ-� ߜ-� ޣ-'ު��o9�Fo9�~o9!�o�H�mw��	7��	���	��_%�;��������� ���$��� �ϯ�x�=�rF��rF��r��W���t9�6u9�nu9����eﺜz��`'��`C��`_��b{;(�������oo��|�x�}~n���_ǽ��w_���?�f?ܘ���L�N:�8#%jV4!
I�9)##e�ܜ�HiB��sR�N�����|�H·��W�I��T!'UJ!Ha���.@��*9�z��*� �sI?��
�Dh�\ԭй	��$a`���}�v��r�+���	RJk.�N�L ����;Q?E{H)-���1�����>��RJK,��0���<�f��b��f9��F)��b+N`��q�R ��bi$ ���)��W+�B`����R =u =�c����R =u =�c����R =u =�c����R =u =�c =�c =�c =�c���#� �#� �#� �#� �#� �#� �#� �#� �#� ���r���1���1���1���1���1���1���1���1���1�< �� =�c =�c�ݣ 3�~��O F�{�"���,�o�QqfN��K���4g/�к�o��`fN�zRӥ9]��g�a��֭d֘�ZwFWh]ݺ$�ݺ$n��ZwFWh�,9����#0�0� ۯ �ˏ��f��f�O�}�\i���3�B���
�[���{'����]�_�����e�`:3$4ø�mCl8Ah��f8��z�X��٥~�
G�s�R�c �Ͷ3�
�n0aZ ,� 6v8�4|ttf8ߊ:���襥� ��gNXjatD�̐���u�����a\w��!:�3$4øI mCt�fHh�q�zr��aܜ��!:�3$4ø�mCl�@h��f7Šm��͐����Q�!���Hh�?Ӏ�a�H��!:N3$4ø	mCt�fHh�qچ�8̐���;��q
�!�ƍ�`:t�fHh�q�#چ�8̐��M��q
�!��ͦh��0CB3�e�6D�)`��f7��m��S�	�0nPF����a�\��!:N3$4ø1mCt�fHh�qS;چ�8̐��|�=:N3$4ØL mCt�fHh�1چ�8̐�c��q
�!��h��0CB3��3�6D�)`��f�m��S�	�0&-A����aL���!:N3$4Ø,mCt�fHh�1�؆9:N3$4Ø�mCt�fHh�1�چ�8̐�cr$��q
�!���Nh��0CB3�I��6�oχ��G�)9:N��q
�!��d`h��0CB3����6D�)`��f���m��S�	�0&�۰@�)`��f�ߡm��S�	�0&�C����×3X��ɴC歷��(�ѐY���Z�RϏ��X�|qc�Y�č�g�c7�_8.����:O��n~H�����9\!��%D�X��t����2���4�yB��p��%6g�͏a=?'o#���%N=������gƌ.�C鲪�m�7C��P�M�t�n�y��A�vG�&lǂ���$�y��]g��������6�1��7q�T�U��߳�_QmV�+�ͪ?Kս��,���������RZo�EyY��(/��(���A�[�>8?�s+���^n����Lɭ RO���@��RO�x�@��#�H=q~��V �'Ώ��ڧI=q~p�V q�,���o[��8?Um+����m�z��䰭 RO����Ѝ9�Mb��5����*
�GG6�;�WU�%F�,�+�ê?�(����� %B�|�� �Jdտ�Y��4@V�+�U�J��9ە������1�JG`Z��v(37�  E�g��mf��
�w�-�����z��̓{JL\���sbZ��МS�@��朘�d�ͧ$mBlXp�)I��|J��΅k}�dC��:���L���5��a��H���w,��K�q��.�ƣ�FW��u���e��l���o����[��L<,na23��,���̄���&3%���Y�hd,�y�u��n�f]b���Y������P������7U�գm�f軲
L�n�;܂�%�,��w,��K���x�� RTe�yGc֎���T����ݵ�`V�+#V�+V�+�V�+�&����.����.����.����.����.��(��kc]���M� �^xm"� ��k�< �'^����P��&�y RO�6��zⵉ`���M��4�'^����e�'^���=�ۛ������q?�|�������÷7qh��q��1�QWcƁa��!�4g���oo8�!�С"g-�bEά�k&�'�&O�Hx
8� v��`{�^���if`Zs2-혖�L+Z��4��F�Әu�Oa�ML��5\��bk�X��>�𱆷�9sQ���/�1�~���1����U,�c����+���A����ax�j���˾��m?Zx���J�9?+�G;ṆK������^"r�f<'!':�yv������;s��^k��>NƇ�	>�u�">n�O)�S���>����P��Q�sr���P��J�#� ���*z�����2���|����C�+�E)Mg.@�[����3��J�j��\{�T����)� �z�ewJ�2̏��s2�.���O�{N&տ0?ڊT�^���R�_�e㓅�Mu#̏�"B��T7�\ 3Ђ;�T?���"~�EV6Ց0w���-
�M�$�m=���0�����Jf���M�8��dI����5GH�	�/ݒ��'[~g����]�PdN&ջ0?�K��ȸT��\{!k���Ku-̕/2B!�Ku-��.2B1�K�&��<2B��t������Ǧ>�YOs�������e��=\��Kt�D�K�p��/��%?��.��K��R1�T.��K��R5�T.ճKt���A_�y��t4�mEG���"t��MBG���&t�	͍BG���*t�
��BG���.�h;��=����b����.�h;��=����b�v�s�أ]��.�h;��=����b�v�s���]��.�h7��;�����6 ?e6?�N��a|�}���Յ�E��v���K��vn�q�㇙�˻���\�͙�*�1sm�Q�4�'53�q�ev_>�/:m��2ϳ�A��͚�W�����USYo�1�v�������w����/r�u�=�*(b>�Y՘��}�b��xzցG��|_���*��S��)�1����c����˓�d���P7h5ڢߟ|s��ߚ�&��<�雧�O����0}����C�e=����O������Woo��|�sUt�/���M��x����0o>�Ѱ��������ۏ�׿=�������|x���<|������t���^X��oƧ/�Ͽ��C�%�	"gh������c�Ƿ��w��{��w[��.������`�H�O!xo9�u�0\Y�l��eC�:B�1��P����������y����?|~n�=����cx��f����)������8���֖w�mQ��o��d���8��_C��S]�~�Ku^ҔӅ�'��s����/���W�7t��LP�k��(���Vfm��*/�����҇�p�O�h��)}��j̊*�qU�T����5˟X�KX��Q���*�w���wUEE^��r���cә���9��T/\Ә����Y[QU��Xsp���$3]�vj�u~��^94����_���:Uu���:�w�0ya�(\�����t�g�\ ������s�.��.�T�"���:��~3�˿�zݽwC����O������}s��+ܷ�����2:Vy��h���8a0`L:��jSV���Xe���<w崰c�9�VH]6���9z���ۋ�L�%o�_���f�X�}1{�%ʕ8��_{�ԇ����;�+���J\�]}>[`g�L��8t���jc�c��R�Ts�=��^�n�\��#����8T����V�P,g���.���@��oy�\yN/����
?�~�J9��wY���6?+W%�\n�����׶\���	z�m�����ͼj�؋s._�;�e��\n4�x/mo���&��=��^�`��\R���%j�܋�]{��\,�U���"~�������a��_�)ve�r��˩/��̯`p�&�|z$o��c�F��mJ�7}�P>�Mhݘu��c=4e��F�d�(?8����~�MG'����G�� N/C�|_�;{�P�k|��վF~�ï5�:���E���ݕU^�adS��1�����X=�u��<�������T��:B�	r!��]q`_��x�})���6��)
:c}� �F�!Np�;��5u�M���y�D!�>V#{��luLd��s�S�!V̫4�e���|�4TgU���o�z\tN{9��Y��rNrq�[��D�1�;�+�Ly~�8\����Ʌ 2V:	,�t���V��X�R������b�w����zMu�"^r$&6{����B�~WM�5?>��k6e��|�,�G�u�gm7���LU��6y�m8._����~��6��8(Z����+y��껨D���ǂa�R����.�9��C�w֐NۑJb�`5 �_�s�����������i��r�KgnʩXu��&�b�����C�oq+��":��:�!�M.�����5]��U�Q�����L��������aY����s��{	-0����a ?]��_��>S�Ӌ�����gl�	�K��\Pв
�����I�������f�|ӴY�6MV]���kB�'aǡ�|��-�<�oM1H~[��i��(�8�u���0�+q�:�} T݅g��P��zM�����N��������r�����"o]Z�Y?ݺ|��]�!����j�׽����DW,�b�t����_q�~;���_
s�Kyz�>���ɕ�h'���+����Juz�>����=�i�T��k�߀O��K����y����Kyz�>�rx��/��;���^)N�T�W�+��=�����k��{������1�w�I3f��BW�pmr�D����z������)N����塟����S������������<~����!"X����I\�_���8s/B�����3����~�?|��������Ͽ�?�� ����������w7���7�����ws�]P�������?��%��	ox�ФB'�槿���>i��w�}����Q��x���M��Ä��w�}w�^�y�&^���|���m��4��2 ۅ����!c�ۥb��I�����n~	.s������:����C_��~[��Xx_��ͯ??{���|��׿����Xa��i��w�ز31�d�nh�'�&!yU��,���<�P��=���)6���ś�h�nu-�a�Ы��8ϫ��k薟xE��_�e�*!)��+���ǘŘ:�٪�G�蚔m�t�72k:�*��u�Xc��bubh����[,�/W���ج�,��1�Xw`׻&�[�Z��]�!�̤�]+�ȝ	�XRj�sae�زO��~ ��c�/1��O9�Om���'-Y>uQ�8�����*Rn��x}�8[�`g�n���,�,"�K:�y��XV�����b\g����@������1�ۭ�s�*}�=�.+�|)-H�b/I���l
�6P�q��|���s^��y��3D+*׻�M]��)������Mm�����1�g����zՆR�M�v��*�!Uv�ׅT��F4��
�<�=[��,�2��~�vI���T�]�������d�t^*9#s1bf����i�Φ���:����Y�`�.�����uxŘc�M��K���xY�����C��n�kL˺_^S�<2�,��Q,.�\jZ���i�̷��7�Z�k��ʷx^�R���~�z5����Um�Q��b�X��[R��/��i��O l��oR#�KAa�p)Țo����,��:v����b�����`�?�٧m^��N�g,�(�V*1ӎ#v,s-�ޚ(�?+����m����(7�n[���q�b�j�
�@�����z�s5?�@u�Śɽ(��>9��R�|_j�Qھ+F��,�ʼ��z�B�em��U
�L�E��
r�٢V���W������R�|Eq��tܫ�nv���*5gR6�yw[K��O�J�{�ZWx�[�9���a�����%�uA9��y�r^�<�*|f� �i�f�WqE.S�o�:�5�zݗ���c�m�,��w憚�l���sUr��N�V�!�����ŘӾM>��Ewf��_�9,��نվ��f�3�w9ɘ����Aߪ3��{���\�z$_�i-g8|Y�.9��0f1�Όw�KexG�}e5��l`��5����)�΂o\�O��憇�IA�ʡ�6w�I�]��N��^�J�溜/H�b*ߚy�t�`���j()x���yƮ�!��7.��?��)KŸ²�76�LCX6�1�9����r���"_w�c���q�e���z4���<��lXĲ�JX^��g�K�E��b�o�f�
K��C;^��;���N�m���lu@�7.��^��u:�U�N��?�v���T�ٰ�uW�f��,�����Kq�+�cKE�v�^2�a��βa3�����׬)��QD���weV)�w�q�ۢ@;o7� WEgٰ�l���R���X���e����rmƶ�O��V!��Ut��6p��,��,��,��e��T��r�z�����h��������>O���������K���?��y��s|�����?PK   �EX ���  �  /   images/23edf803-1010-42bc-b391-ef0e69fabd63.png�^�PNG

   IHDR   d      ��{�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  .IDATx��Y	TTg��jg-�b�whA��-D���t4�Q�����tt����̨�9mgr8��q��h�v�%qk�p�MQ6�}(���*���ﭢ��$�?�yū����w��woɛ��G:; �J12b����ɳ1ѰZ-��l��I����;_���pU���;v���.�P�ȍV�Y"�$����~��E������7nH0�y�=���/=�0�w'~t�����N>�:$�XG�P�Z,6+<|���R�������b��?E�3x�v��\�׋[��⟂8�81���v�7���澺�#f8ɝ&^�E�l���R�'�!^!|�`6�o��a�S��ʤpW��<��A[�ak�X-O�)�J����'2t&����I��8�پ&rq���0YMz���_��;���#��1�.��v�C����}:���fti���b�����^_�
C�;ˑ�I�L&��0���z�'dW~�pu������������.W;&q��D`d���ZTvWbY���H,bF��m��Q����q��.f��B}o=+����ξ�T�T�>c+�]�ˈ]�.(�J6L���#��=d���/��a�Z�AQ�������6t��].�^ð�bs�f\����rx�C:��t���F�Q*���5����!$O�!!��fo�G�m�P�	���())�e�,[�=���}j7���n(+�LI���?��W�p�����N�u���?�f[�T�U��7��6���ư�ޡ^��6�w����w`e�JV�J�B�{�z�ثI����*1hDs3z=���cr�d�n�� � V`��
���#�"��^^���7|]|y�d�~S?t�:�E]o�k`cz�Y�6^���	�l�]G��)d�]ʄr\H�S���b6�&�T�V#""OF���&6�GȐ�8�x�8U�H�z�	��&���K�7b���3hT^h̯AN�wP��<��h¢�xg���r�5�{t��֋oI�k���r���t[����>�>�NR�_k�ʑAF#���m�eݔu�6������}D{E��Ș�Ĵ�44�W�k�:!Z���`���Iel(���9-�3wZ� 5 �����=�=����<`p��s�Z��$񞐳B�"^�������� ���8�`6������ ��MC��op����p��u|v�R�E�\Q�_LZ�4�$�/T�TP*G���M��<�pL��d�$6Ʊ�0=d:�=^�؏������0�8n1z{l�#�0�0����h6�*��R�ā%8:~}���%���S6������Y����T�)�u��]��h�e���!{}b@""=#�����GQKs�����W	�`2�p��F�M��8N�Zw�I��g�ل#�	'[!޵B\�r�.U�B��j��8�d�@�P⁹
*��nKѨ����_�Q05p�X�Tx������e�$����.< �~2�_¯��DÖ�gC������{s/�7_Ǻ��0z!C%[��0u�u���v����t��}b���3*=���!Fm����)?�=��������2PΡ5RQ�z�7q��<~��Y0��Ϯh��	6\�sYG�-��C��U�
�J�z!�%Fv&1ol�k��/�l�c�!^n21�id}R�6�-�=�S����M)�W�l�����f�(,�|���Hx��oh͓�
��'�?a�Y���s��a�mlC��V��r�e��C>�F�E��n�)2f��:����d�I�=�C][V�����
`K�l���a�"�7�=��aֵ,`�6���6OیMy�������3�f�����ވ��e&Fq��iN�z�p�@�w窊�
~�D&A�&��A-E�3c��&�:�A��+"B��m�P	/*�ӝ�
Ŝ�ټ����ם�Iy..�9�|��/�����,�L���%�K�?1�jd���G�GQ�����W�fc��Y�#%G���p�p��αiEyEqB^��U���f}1���B�fnŮ�]���G���GlbhDH�Y�p�+ȭ��d<5h*�<����o#�+GMvy6j���
�'��������E�Cuw5�9�^�������I�4�7�H �h�L�ʎ�W�7�c�a����W�by�2�<v)>���`9Z\[pBwh����[����/o�`��Ӡ`,"��}�!�9�|r���U�c٢��K��e�n
7�IY��?8��L��h���EL�����F6rd�s�x~�y��z>Sd2�ˇ^f���P�V��mi�Rd�ec㩍8��+��W��D�C��
��<a9��M�9�(�S�d]�BT`#�N�q�&G����)�	9�����k������%�"b¬R����$���ނ�Swb@�ărV����F�t�9\�pr����C�쀗W 㲅��r/�D������Õ2%G��,����VD���ه��<�d�I��q�ġ�q5.�_��/��FD!{t�Q�{g���.�E�p��[�A���bȜd�3���Q&r\��l�y��ʭg�bZ�4["r9L����3��'�䟄y1�p��&�^� M}Ml�ڮZ��
V�B�A�ҖR<�?ƌ���I���3���̢H������##7&�qH2D�����
��/�mBk�}�[�ɂm�HK��ۏ���o��+^]0[`�5U�HH���
��o�~���B{i�ҧ�*ʿ����%eJ�f�Y�yyW9Bաl�42.1)���~�ơ�[����ј���������L��:������N�����ը��ȡ�#G����ɘO������(4�w_ލm3�!K�ŵ	��H�� �����B�'�&�"X'��}�b��!1�M�<Q!D5�ءD�����^�[�%�j��o>�N#���%��|���{�WQ^�Z��(�-�G/E�O�~���ٴ��ab��V�6����z�j�w��� 닒/uUأ\��������F��ކ�;j>.�x�6������R�O�R~bp"����{G.A����yT-2q5O���)��,ğ��̹���ʶ�oo8ɜ8Fk%23X���"lm���u�6��ڊ���q����HL���p��$���>�1k�D��3S��}���F���48�����d�?Ǭ��عb�RL򛄯J��������X�����I8�/���D"q`4��h�D&��h�d8�D`�8(JV�.ۋ��7���>7�Ehͤ z��'�{��L&[�*�7�!��!�Jɝ>�&�L(m/�"�*w"^B?n*7�\�,P����О�KH.��"�5�'G�!c�����������Cs_+�jQ�f`�PZ��Hפ :)1�	��`��x����IMFX��~���X�BB�����$�4��a}�z�)$���m0�&�7@ᾧ`��܎wμÌ�DJ&��	H��?���?]������A�p���T���a=�7]g�9080�~�6��z��P�U��
fZ���W�ƈe99�>���MFe����x�	�
y�::v	�4ו�[mB�c+bb�X�[��Q\=]�]܅"�B$��Qp��ҋ�1-U�%�R���{����(E\\B#���4,�������1=a:J�Kh�j����[��ex˩��������}t�(#4�i/y7%G�k�r��9�<K�Jm�[a���Z�T��h��r��	�h�Gă"��`20Q!�r�Z��ی�=ǟx���G}��R��k����l�i���]�v��0���4�����������eX��p���!����6+��g!<�V�=4,�=�xyv:C�X���}x�[?� �Œ�����a#�%(������m��ʘ2�!��R2�4H��X2=�	\<�e�4���:�n��ĊF?,
�#��ߑ��Eu{{�����<":�n^?����\��d·F|���+gg����Ȩ4ȔJlH���0�x?eP�@(�����u�uO66ڦ����4�aإC�0��J�z���R<��FY����.�=�|#�3ؒ�c�?�G�����n=��    IEND�B`�PK   �EXR+`�p �y /   images/29dd1623-773d-459f-838c-8b03343154c4.pngL�XT]�?�4��Hw7(݈4H�tww�����ݩ�t��tw�{�����8��ٱ�'�^'�4*22����G((�e((hlDx�S_��,&���� �F��#9�h;CA�uCн�j��IBI-U��.�FNfP���,�v��&Ff,�N���BDPPo�d%ޫyd��k��]�����˄���Ag۞˞��f�; Q���i�C3ɅK�x8�!O���-*���F?����1��e*�ʓ�|#���	'��~:r�1�����#GЂ1�)B�\�w1C���{�.d� ���O��D���CO��`n�x��#�£A����Kr�o�%ׄ��%�WP��U�Ď0P7���m(A���RH�wu�5m"~�<4D�8�Vs�
����|syE����GO̎NL�*-#-!:���w:%e(�l)FA����o�A�U��ը;#ha�������l���)��#h!��W��wl'v����œH�)2�1�$�J�d�����ɄK�b���\�(�.)	zA���U���=��!�r?j-�4�_��:��g
�8BQQB��ęp�$��P��-*@��0+H*0\'�qd�"j!rWw��ߋ"r/a�\����?�#�8���}�?ܛf.B����o$���v��=�X ��,�1EGhGM0eW,d�T��إޔrȻ05�iDbb�o=��OB�` kT�S-;HɰdМ�(-��]�Z���b��UI���~�OR��Eōes�()�7l5<�v�\��$R(�#�_�KC��Vn	͂q���sZ���0f���S�pd�����u��:C��x=�-.Ul�d���=�)-�	�����Ή�Ҋe0C��1Gr�WSK��L��W�M�u}��K�Ɛ�Oz����j�c\�x�Wy�7!U��٤}�❯�G;�/N�д�x�����\�P~��	gV��x��a@�2�N�Kؔ���,>z��ɴ��'3|���E�Z4�XR��8�����ˡ|�9�p������\�^k����A�GK�����O@_b坆�ǧ�y~nW�y���)F<���/b8CS��\�p~dT:�7�|I�Mt=��ܮb8ɧ�OU�=���]�0#h�Q��8<+����H"r��.��d��P�����_N�1��?�m{*�2��F�%�2	R��:�[��q<ğ6=��������4���-�/ɏ(������P�Q�`���)�����>)|r�:��a��F��s|s�t݇��W���+�|�F8�	��h%�p�*w�U>R|��mH���'gD�����ѣ��۪G�Lڊ��H3.-!1$v�݆�`{�c��e��2,�fI����o25�g�@v���t@t�O\VE>QN����������x����_�\{������~���g���S[�)��Ka�P��m�'^�<v�J���K�~i����Nn��t�)�O9�� 2ڎW6�v�t�����$�kj�Hu�߃���O��Q�c�ଃ��v:��AYad�Cmh�oַ��4����ϱ�6�gS�!&�Қ�26b����ߙҢ	�0G��c㣜�����a�v�'|L:��V���GT(w��)?�*ژ}G��������K`I�-3��[w�m�~Ca�Q\I��:/��烶����|�� 3����T�4�	�A���F3{W�(/}���\��W�=�M�f)8$@F��\��5S�p��_�[�>=�z�_��B���jޘ��r�Nf?2���0�uo��]�
�X�����a�l3BN~���z� S��=�}�5�s@c,�UwS��K덨ĎeQ��N�Y�-���<�> 8x�e�OU�6ӎ U����|zL�B0<���qߓ�g��x*{���x-��`䪡v�$C!�\���G��?���>�s�|)����Y�}"��#��S�y�g=Y�Ʃ*�=��7r��m�vuU$��fTh�2`�<��䱵~���F�g�XO�|�p/ 7X��o�nbfB���$;�xN=7�̞ڕ:�1��)&9���{������"��4�;$��)&��Yp3j�t�V�rgFD�L$��:Im��EC,(-�;�O�Z(8;�<��L���u��Sd�/d[��/����fG��&�>�G�'�(�ū�c�.�z,B�B��Ǎ�BV(L��~WX^ٸ��pnN�ģ��_8���k��b�x�@�〚����tW�'�^n}I���U
_)��V������J?�M�͢| L-��hy~BA�*�7�2_��GW�bˈ�<�+?���(�����0�G"6���;7�tb�-�����ϳ�0O���u��eJA*���1�����arlM?�n�hi7�cLjy�%��^��r��,d���l`Ԯ"�"V�*�eyo�׺�{[���s������	�tbv�ƿ�R�堉W/�s�M�N�'W�_O�^{SK����	��ŨI�<��W����O
m��<o�������L�������x_����y�Ǵ��Ԇ�fP%|��Q�|ut$�#H4�����"��������̀Y�c�b&K�ﵮ����!�]�As��?)��:��$�!�k(Ho h`�4��ܻk��G&W���ka��% <a�׊��!3��s	 ���6�e���tK�w�uQ����z]���/�k~�\ۄ+ki@.p-A��p�X�.~�x�tF��W���wºn��ùܨ��S�s�a,�\��ef(0�0��]j�8���l�<��p1��6�Lr�_53Å�X6H�
VĄ;�e�TxX�Y!3qoi�P<�n�[��dA��,�J�Kn�ssF�d�������6A�����
go��#��F�g�4��3�cw�{�S������H�"�is��C�3��\����K,-�r�����)�t��%�k�ty]]��Θbx&�&M�M��_��4G�s�S5QPPA��`Tf��� �C�Y���N�)�	w�y��Y�{�dl/�qɁ[W��t-OW�Qu7����4)��.����yJ�:E�]��M�ݰ7�7"~EK��犲��P�n`�� A
{�	���=�am�(�!��V�+1���G

���o����o�(����m)�
�C�hrKڏ#ٞ�]2�]�����;�͆���PLlM�Dޣa6({�B}5�J��F��9"�oe�z���m�2"� 6���Vh�?�4á����!,��Z��,�vt�0M4�f�V��"H�"��P0;����K�{�p�Uӵ8��� ĵT#�K>mk��,~�I)�$+�dY#���[���1?a�������KE�jh홹#1U1��om�s;^����9�<s`g�h�P[���2�<��2I[�g�{|l�M�u�YM�}���r������2���'~BÞ�@2��(q�S�[���˱���o�{h{�߶�ñ:���m�������.t�HBe�H����F��yA��wk�A�Y���I5b(�놪3</!�y<�/"/D'���Ug�>?��E?$
	?W��/��CE)�j�R�3��0*ä&�\�#;�t-RX��X�B�i� 6X{"z�>��1%a|�,Bn�q\�m��~�{�kv�v�u��QL��䷐ee�׏�z���m��II����g�g�<�Ø�=�ZE���=�2���h��?wd|³+X��h�[ğ��;�'7~�B��*�*M)���Ǜ~�� �P���?�H���m�V=�8�6�P�;P?�:쇘*:�m���[�m����E�g�s��Iq	�@��&��Xs+�cظ��'3_j��5���;^�A��l.�,���e�C�P�)����F�#>z%=c��@�wV�#�>dqD�-���?
�%����_`*H� !���g2�����Ъ��#��Y���9?��M�0@k!G�ֹ����k4������*�<qs���v-�y�7���S+u��v>s�Bt�^l�q݅E��գ��*�3�C��ԇ��M#�4g4��MA}��6���@%�$�nu�׏�����[n�����ToE$
��p����
�#�rȁP�{p���� �@����� �cDh�8�"�������Hc��y=)��mWr�n)���%4ӫ*DbLh�k����+`�"� I@��I����V�V�?U�U�p~b;��lh�;�}���??`�Z�c0�a���^�hEgc����k����M�q[����7�x�b�j��vi�2`sy�.��Z�Ə�	!.z�ki)�ɵj�t8�zv?�y��9�f�c���,��������.��a���H���%�q���|��x�p��9d��a_=�V0��t��otr/��%�"�mT��H��C���Ut�S�-�`�%~!A����ר��(\���f��?�{'�0A�g�' ��oJo���F����0����E�@�og�p�uJ&N���~�5<����@ q�3� � ϥ�i�:��A�!�<(cZ�N�(tmN����(���"�7�� %�?R�FF+�����kla��]ͻ�4��;�9M?�Z聬^_zX3��R�AT����k�� g�m���8�Y%���FR�e($v���.�Y�ɩ��eud�Ю=�n?��.VKyr���hXT�A��-�9�_��Bb�ɕ��z�E�5����"���a������gZPi е^ڗA)�)E�W�8�f�!�@yY��:l1�qRqU�U��_Q�&~�Cd���Z�'@\�0(�̠\tH�74ҝ������n�KC�n��-��G�a�x��G�X2���I���s��[��jӚ2��e`���R �b�E�5�4@,�#��O���Lt��R���H��B�i���- 1�='�p1������9�l�1��z&��Zr��ӆ39�6�_¯�i�~�����h��t����2���~��R�f���V�я�����9=�b�.�3P�6��]��#�&�ܘ5�:�����b4�����B��o!A��]��=/��ژ�'��K��f0e�B���	��;4|7>�̆YȰ�+u��(��g��/.?��)[)pC�����\E�V����5/�	CKn����о�|盈o����p�P��/�D�	J{�3��՜�4�9C`�TIU�֋���]z���@ ���!	/O`b��A��EQ�A�- ,Ϸ��hp�eb9�!� �jZ���*FTR�E�������by��?��b��>8gb������Vz����$lU�k�ԏ�f�����M+R�MІ/SO`'<�K�]	�:���23�)dt�5%d`@s����	���
!ZY�����������u�:\�B��71 U&L�+l�������� ��j�)�u��!����x�h��ҹ
ăT@#��0����n?R<�\�pK��<#V��M�q:Պ�P��tn~��(����b�����w���'���4)>d��>�����{������8T�5CQ-тvDh0$-aK�Du��K���0S�����u)�W��t)qM�r���;# ����nt�5���@QV�:e׈S�_y����� ����]���TW���=6 ���zm�lR�(�,���|`5�	{�~����-�������	���RIc����in6+�e�3�}x���Fi� P�fjed�w~������M��/~N .��4��1�����B���1&��~��[�-�ԕ���C�ґ"���j���U��������A:�k*����ZB>I�8v�rW6{��<��@]�;�wN�=�i$Q����X;=���p��,Y�C�s�dע+��y��Qr ���W�pM/��y�F�w�T�K�z���%�ݻ=������_<Эf�3�06�R���t�$<�V��R�Q#��>�p�c� 쿸�}�;iš�Ĺ3�u��mOW�;{���	��v��95�'�ME�/��>��@���;̬�w��m���L��\��Iy
+d�����t@b-E=S�����(���kF��]�ӻOI)x?
sZd4�0�h���K��"D��#a�"�B��w���9+N�UF7
���cCj��)�/����j�%E5v4+l9��1'"d��2�l�A� rq��C���2�[�}dse[]�����4k{9�ڟ��/��b�}�������yv}��K
oG_��D���u��'Y}?G�7.�r��ƛ��1Z�j�!��lW���1�Ԅ�.�ץ�Mv[pvccMW�̐�J+\S.��oyE��(1��EI��K��Kɪ��;$��?���x�\��㳹�up=V7����9��0ꤢ=�T��B���m����2�;q/Ng�,����_��������o�Ը�:��;�N����-���3�k	Y�i._Ϟ�$~ȥ�䚚�X���>	v��S_\9��d�i+�**���� ����i��F#p��E�F��C�"���J5$�ȹbUh@��� z �B��_K��XR~�˴������.L�������(�rFI+m�h$�Mר�'P6s+��9�L%5N^�4T�eY����/>nq�l��e���f406>�.��y��i�
��׭w�|ܧ�3��:_��B*��=�L=���>����!�~"�W����yH���
�̐Od��r��k�)ߊ��o�S�)������Ik�U�Ŝ���w�ߖ}\iv�>��#N3z�;1�H���]N���|bS��Ax�`���r+���v�p������6�8#
�¢eSʹ���qD}�)�2��5Zr��dd�xEV�P���k8�.�AfX���Y6����%@��3
3�D�!�]�h������eƵ?�\�ɯ�$Z((Z�_.ّon�\V�O�=��}(�W���/\�S�;̈��׏��'K<�5,4�=��
�XF��1ߣe_�J������n���R�1��Ӝ��
3rtNms�#~���@G�é���Qn;Jb7�>We����+��hf�)�)-����V�����-]15X�v�o�f��0�f^�� ��/�'x���7�H���y�$�A�T���ָ�cI���+�m4v�\0|������B
b�����E4i�V����	\ؿ(��$��DX7قW�d�.$��ƙ�0u�J�k��������1Z�?s���5�13���ve	#Ǖl�9���]t�q�f?���KssZQh1jYrQpN~�m�g�F7{7�{Z���w�k�S�����(lU����'7@V��qv�y���ß�M���8����y�
	��<i�nq���;�q��q���V`S����{�}�o�4�8�F�d|��ǎW�9�M��؅A��18�V �9�ہZvUnTf�PUOmV37C/��(��Ջ��U�j^�>�B�$���9�X_���չ9��8D8���E\b��B��b;�s����բ��?㿫~&'{����?�2;���x/N<z�;Q��$�~+&��q������A^�<�H���
�じ�Q�ǐ0L E]�(������`�����Tz��Úz��n�a#X��K�l��o��� `����(�̍�E�
�U_�t�t�嚳L1����5h�a�y�����VOj����6�36��M�I7�8�)�ڤbw�fpy�-���?|t8��t+�N�/+ �_U���N���_ph��B���@Eb5m�ﴛ��7���F���^��\�Y(6�����?�+��CX����v!���{�{�M6X�P?:m�A�v���i��������)(���0��aqqbjB���$�:�C�K�"{Sv��u�;Ȯ��b�3ߩ�F��;	�*ٽO�SD����L׽[Y� [z�H���<*�B2�Q�w�?JV6��ݶ{.>Ly�ٵ0@�CBAu���Gk��@��Γ��ʊ�*̜���N*V�#�3�o�vn69ց�[/�b��+�Fߍ��4h�.�dE_$(Y�+��9�zp��Ab����l@���y���`���QV�>Se�\!Řj���Uq����'f N.�˫����a<X�K�K�X|���41��J�b�bY1cYJ,y��,Won�"��>#�w������tY�ȭ����EpƱ���]߿��]�͍��<�5�� y�]�l�����
F(x:L^�?J:�Ψ]�]��̑�")Z��M�K"�:O}�������q8������~Y�Js�"J�y3�^�1^ �J04<�'�y�� :��V��������H����Ľ�r��.��?�MĄ:O8��=-��˸�A��P!�v��ݮ`��=�����,W��k���h11���iN��4Xy.QWG*���*)�o�g?UR��! S�mR�QFǫ�,�;炔����'�'��>\r,���e�=��%�ZVL-
�]#,�W��sA8b��РVJ�����Vbܠ�\�dyn��S��rfl&{�i�a���/ё��O�1Cm2��m��H��5��s��'FsS����ps��#���fꌊ͑���S�z5����{f�q���V':�/ػ n����F�O��$��z���S4��9J:F�F�hs;��@������Y�c��Y��'�氼I�:���-ɧ����������� Ud�����K�z.�v�*~i8�՘��Ʒ��	��v����͊2��,$ML��(��w�!��V:��nn���>:��1'��Q����r�;5�CH�������vO�,|*�f�G�%k�Q�?_�'�R�N��h���ӆ��Ofa�N��Akޞb��B������ �F���h*�"�/^�h��I58�I�'?
1��U�� �e��Mf*�fTs�HU�E�,��9#�>g��&k[�r�8��c��t�����*9p���޽Y�k+�3�&"Z���pˈ�Us����=	 �o]���w�j��Z�@��w�#�!n��x�P��s�s��ݷq�>?D ��Y�-lD��dы�܃2�����LW[	c9�~����K�$� <���Ra���o�i������3ƍ,vr,��E}��.��$�L�Q�&�&6��x�LY���<�$'-�i���613
2�f�F���$��W�L�$�5*7j�)[�q���7D�?,� 5��|ŀO����ţ��+[onb�G,h�ss��%�����	����v�Ī,m�H�Tꤢ�5r/7y�yd�v���+�*�g�ϑ�����,D�o�c����=��4������4���Y7��G��4�^, @7�nBj���u� GU�l��䆩��o�1m��A9$�$V���#0�}����C��U�>ԛܪ�E�k����G�������a�g��3��g6����Ce�i�����x��^<!~w�1���O)b����"����:4|�D�z��nȝ�2u�h~�r��	����q��d�V�sN�n8p��R.��Ȑ�{��N��*�o|��oS��v���ט������8?ɵ�>[���'G��ez1��#O�ы/߉�R�D	�+�k�-[Q�����<�&�J�k��F�$g�.�ƃi�U]X&�1�kY�I:j�TN_	A�/|[Hu2Ff��V�O'G�&��AA�&�ܢ�5�M#�b��,��YT,��	� ���M�?�2�?���P�/�Ƕ��jM,�*=�[��+������܆C��4o�ݞ�"�J�;U�}W��l(l3Eֵ�sN��������@]gD�s:�QK�N���sZ�{v ��3�sNg_g3��d<���Kh���
W�b�#X"4`�cyw���-R&����++Դ���;�^U���9ߒ��$�8�@�'����X�]@�T!��������>:�d0�������j�!��wtP��I�����Q+o��}��?�O��T�Sw�:\Y�[��J���,uk�˽��5���;�A�������(A�[���|QY%��l���+��$A8�s/��0>�ߦ�/ɦ�|xCe��%l����)���.]��#��������c�������$�=��E\���-c�0�ߐ�����	>6>}G���~zY .� ���:�ҝ$><_�[{���f��*�Zh�ܲj�gx�g��~�$�,�7�3nfo�=�3�63�)?�$[�/ML*J��Rn�?�� ��e��nW%vq��Hk���� ӷ�ws¨V��� b�c��!=D=ڰ�FtW��[�WtPg����ܷ�R�R�d��U\U@_�,��~�]\�ú�i�iJp�IIdٲ��G��j��}�`��M��j��cW�cLp�����$�x�q���Z���l�	R.yO�8E�y�,�>��>閼բV�c4����j�f���x�!���&I�JT@���tk�5��&l��nc� Mr�^� h+��X+�~��	�$U�0�(��]��oU1���D����F�!����8P��mӎj~0��9%��I���Wx�Z�;.,4,�%�ok����W���{��� ����<��SƵ�i��T�������V���@ntt�b�~���YZ	GR
/�{3�T6�����[o%<���J�yڍ9��]�t���7{���x��U�B��ؿ��}��ѵ�m�����3z`��S�<'Qqycd��T ���,���sߟ�D~o�P�9ܢ ��l��'��k���p���3�@۾�w��Z�3� 0i��OSlb !~k�u�����:3��/�܅6q����1�M�hg��r����i|�!�ģI<��!�>�{�&3�Fh͚��y[���3�dvQ[�Օ�yI�lZ��cXb5vF�ˉ=��g{���wt�䴑��V{g�J����{����p�����,Y��AN|��S��{>La�Y�UMׇ�%��>$h��6���NE����Wܤʇ�-�S.	�H�y�gtF�qt�K����3=1���]�}�}�P!�l(Cvv��Q����]����$���L�(��"����R6�C�]�����L�O�U��Qj�Cj!�!��`��[�����p}pR��?j:� �h%t��6$(AȼC��$l!>X��/�|�m�1����d���Q�Iʱ1�u��h n�|���۰���W~��Y�/��QFmX#��>�?,h�tv+n��,�[y����+��t��Q� �_����ͽz�¥��آ)�����5�˺=������8"�-�|�y~G�L�?T������f�_����8ڛ�h҃�g���׭�$���}q���(ʕ�M^2V"���R�٬z��\��/��⣧�rv��$���
���L.�'�[������Z��ʽg�������ߙ����1ZAG�{�� �Q�]�^��|[%���:�17��7��]�&W��=U��63{�t���� ��H-� �����Z��/lQR�c����� |�]�K(C��U�hNW�����#ܧ����#��ss	TV�ʁx�O�$����l������:l�,>�`�AK5r�\`G�����cZs��n��>K� ���#�`n<�O��ÞZ(x��@���r ���nz����;4|�mۆ�V���O��CF�p$��	�	���'����
��q�m������<i���G�-w!Q��0þ�s��`5�M)V��N/?a?�GN?�sF����~�S-B�r
���<�m���z�c�/�$����$�X��.�˷��n|���
�[
63h��ݥ�0�c�y�=�4ތ!��W�_]��@�:]�(�����|D�D隆�c͓�ڕ�b�8Ͳ��xB��e��8Ӊ��L�>�����'��n����[�!�dL%*S|KR_T_>B�z�K�~���v.i��kT~P��Ѷ��4x���,&}q�K[�;[�u1>����yԒ��nPE�,Ҋ��(��$l�������Uk�Mx|�5���rĊ�%��MŐ��g�t���Tm*uz'��c6�vC_m��+'���I���O�8����Fi;�i�q��o���k��4oYl;�8�?CY)��z$-�B�D�q���l���K&DBZ���fj��P磅EkB��J���!�!VjLhh���QKДޕ0�� �yJ^�jh�=���!�ڌfNS�d�$]���-����5ݐ��oV�U��{F������@����ܑ���B�fW>����P�Lm]�f��h��3L	�z��0�58�����^K�=�c��76��ۊ6�3G).B��_}K��7۪�%�73��:�?��0�������em"����m���/1����]aTa�=h�e�D��!�p�gL/��ڿh'D.�,�5�K�mFo�,@�嶝>�O"�#��:m]Q�bEnI�N^�44TG�=��@���PIY��?�W�����-&��{!�V..f��@�$�Z�x��(��Ͳ�mԕ�4����ۉkH�����dP��IM�'��(է�Y$�x���I��KՓ��˴�tGM㞧�)�rF8(�}���o ��ſR��<�؎����\���������2�z�ެhupw����q�~�4���D?��^	���O!2�5�ԟ��"!�{?�^1��� �A+����Fq��Jtk�A��]f��d��{�
���M����XVj���A�H^�>��Ÿ~C���7������i���zlk��A�l�Qe�[�:G�jFPϩ�P�i��˪f\�.�[M�}9��G�ܕ���QbR��r�z��
�C�

ۺ��kH�%y=)�x9Åp�y#b$�gt3EQ� �"�kt����C�$X>��wSP�������n�;��ĪT��_v�;��AZ�Ʃ4����s��xɯ�5�^�������A�U�Q��Ŕk��,g���7v��Ҍ���Y���$%�����,7^�@N�.�׳���Α��ێ�X��n�z	oy�+�M��3�5I�����fW>L՟� ��GJ϶�ȿ�ŗ8��v�C�~�̃2�`v�Ge��A]�@[����ikA҉R|�S�ւ%*|/����!����.��kcV�{�7��_��̩�1��,r����
�)p��N��ot��L��}�Doɴq��&껸-S���n�o��j�U5�/���|��7��w�u�r/2�"�Ą;0<Z;�X���sjN�weWe�V�5\�\ɺѐ�Q�8:��M1�2'$ [�%��4Tgҋ�{QxlH�wZd-m*3����~P�ض��V1/1�?��:j$ZQ�i��`nă���m�A
l}_%��5a��4��\.s>�:�p���5�;�	)9:{m�i�ey�S�Y;��,�_!d����C7�av0�O��[3�?�u Ͼ�@�8
����'���#������x_^I`M�54M���P�Z�V-Y-!�
����6�a�2��Ī��v1�B�u�����o�ix�>�o��,�PVɩ�)A#9���h���!��	��H�E�&Y�T�B��PGP���`������ܽSm��f6,��>�e�1�3/�=6�U�)���
i���z@'��Z P�� ӹ>,<DR�������C:�R����_ېw
=�-�4��v��!�H�bH*M�7�C���N�^yn#��'���o�Z�@"B�&��4�� ��G,�
oV����|Wh ��k9VoU��-�$ۿ9��Xʗ4��7KI�n���/Ƣ>�00�����.Ww�瞇��	Vd��Rc�Y1�,G�my2&M�i`
��'��ٮ���0�0#�m��8�r'[؈svB�4'DqR�F,D�Tw��O�G_�5�nV��o�G �S��^;���n'?Dy~�-./d��F��P:��i���Ў����9�|��GE�����(a.`��7����;l�l��j`���1�7{{���G�E����$��4R��C�����ն�}��y�&��\���@�+;e�;��@�s�J��U�+Ee_�,n��&T#g�+5��Z���n��� ��{�>�.�ג3����XO^��=w5}���_�G�s�]�g7LN�%EE�7�ףK>�{�#��cG�m(��<�z5����2��7�\ٮ�xjɻ���͓��G��-ٖ�م�}�̺��3�&�%�J#Q��z��H�xsW�E�n�%W��i��i|1�w����/f��R�̈�]�)��c��N�����꬙O�����>	d�sWIw�D�����ݹ�Ӌ�ۍ�ָ�O�[�F���DT7��ij���0��b�#�E�ns�4��֞�y$`�&-~�@hH����\���tV�?K�<�:*>kI����v\Z��O=�@���D0@}H��p�����z?�ZD��nH�m
��P4�<v�t�Rm;��"M�UG��bu>Ч����,*��@àL�o��iO��1�a𭃱�g�i�*�>;
>58S�D��F�5%j0������Yz�Y�a�m��������,Rj��5Ӭ��gn�;��M~ ���rc�ۦ����Z��bI����v*��_>~����6�_���>bA�W�Ze2����jV�?��$V$J��gayKGy=@�jf�D[�g��Y�� �קw]�F�s�Y�����Ăd�?�k��tJn�ۭM�9�8i�Ha�p$�>�������9�Ύ��>g�����L0�J������(4��7�)��v���rH�"�y�����*�K�F�C��5��Q;�2�M��m�F��/�bȿ����!�ZuI���J�vrl�j��(:<�e���a�9�5��r6�VB�(���F�DS���/��
6*=O�f}�H`���I=%.������Y^;::�(+#��\ޘCn��9v�:�4�8؋����r���E�Ѭ�@�����l��@���eQ1fe=S�8��ϧO�"!���Δ_�b��k��!���n���,(����nj�^:vՋ�f5�Oo����0�˕~Ci�r.��}-��}����-����.d�H�ܸ�7#��Z_�@�x�`m*?�GA�"3�Dh���	���6�ԋ��m�wd�w�}ά������qE�w��'l3<�.��̏�ۼ�:rop� ���j�l���{�w�A$�"a��<�h-}�I:=�'	�KG�#���Aj�_�@B�Bv��DnY�!S��x4�y�g�������!)�-\M�~r�Yq��L��ʇ���m\i~�������Pm��*f�T�������[��QS����&̛����*iA]���^[f"��R���O�{'!�����՗�G7�������9�S߼������p�/�y���8H��"�ػ}r1���F�]�{쏩������kH����;Õc)-_!EE���`e�(ȭ?�R�O�Y��f���������rV,񑤺�ۼ��o%�RRGm�BJpEs��ݽ��HLj~1��b�R�\a�3P3:Z�w�'���f�S����y������J��<�]�^��r�_�\�r����Y�e0��Ӌ�͈��-��פT�E��9!��ܞ��Uy�G�!6��F�G�Ү� �V�\�Ẽ�1���+�n�8\ǽ����ꎞ�cۣ,�����	Sˆ}�����x�/���5�0�/����p�f���d\����_yw��^m���䎗�U�5�;�L,��T�e�΋ِ��8���'��]S�=v�����ܒop�%� �s�`y��'��4O�MX���cn4N���ϔg�U���q�3xF�n�M*�Z�iz��.k����TLr3�[���k�P?�*/_%h�X���r(q���Xx�@g�%���z2N�W��KE�Wu��=���_��bVcΌ���;��O��=}�Y�]h�x6Р���~�-�7+:k_��GG癶������z4��T��hL>t���Y�4�d�$4����q!�m������
C��&�w�;q��~F���}]��[h$~�������W�ť��Y��s�,|>hdf�br�����@8U��Y�Z_����c�o��z`����z�\��;C�l	ug}����y��޸nl0<���%��m��҅��$Lmyf���������/�U�wVw��KV�	9��@z��g�-N<�iE���0��c�>��U�^�����9��4D,�3�^���������e�Wɸ������.����<�=7�;ޔo�Y����D�c_
��wĠX�)��A�Dr�"��U3� �}ʗ�Cз,��f%l�u3�ϑ"x_��(mSUƧ�3�"y@�s�M�%�
b�׏�D��p8�<�cO�OS�?�s�֫�J�s,zr��	,��<=�^������J�6`h9¥���\?�Ǫ�<R�q�	��?�R��{�#�a�ٻ3;�#Ҏ؉���U/|��g����l��ȉ�m����
��u{6Me���"Zx�]~�K+�^��}��H��[O��x^��E*�d�;�	T�gְ!O+�Zh
���w77�L%K��?37����,��P�������P*�X�&Qk��O/�z,�H��(���(��'���IL�a`E~��7��� g{��yD#EJ��Z`*�0$)��O��5��_���p�!����Z�����ǂ1�?��;� �6e��"B�"�)xJṻ���[B�]F�� ��˺7�t��=���U���ދ0�|��_I������H �z��"yC�_��'�FH�T^�����'S�,C�u�<;�	?Z?
��˝L���w&�ۖ�"�O��<�Ә��}���\�>�!�'���k2��]��,���=~�׼�D_����"�1��繫$K=�T,iB �p�Q�3�!�(�r�9�o�K��W?m�������Y[;�����h�NC� �-��@�K;�Oਨ��N����>+�2Jc��7�'�A�m)C�u��K=$=W=���b��p�?Iqq�I��K+�?:�Eͭ5���K�D�cMz��l�*�íz�;�l0�KP���x��P�"��X�\(����!�>�Sz7���L����q����P��`�G`_�)ɥX=޲�6J�S���+u�Y�b�oV�#fq���W�uS�����M5
.~��f`�  $9��Ϣj�O��92� \�0�@��9}Yh=�*�@__S��Y����s��Y�i��*��"�-u��"X���(в�H�VwJG7��8O�+d�)x���4�ѿ�9�<��G�W�E�|��-H��")-�%�t���t�H7Hww��������3��}~�va�ޙs�q��,����Ֆq��ӶX��f|�rx�	l����?d<�"N�$=;߭s�y�c�R��d��>�=1ЕuR���e=�-F"HT�x[�t����t�]ā�47L�����?�~ҳ���f���,U/f�����;�n[`�#��e?�en��M.�
^�^O�G��T��������zE@���ܩ4�%Ey5�%��Ҫ�5>�\�Hq_Sx7-�~ �N��'���+8��;����+��;�1n�N�p�5�L��0��v3U^�	>��ͽn{]�U�g��������X�c�+��RI�p�q�UB�F��*�.��F>�t�T��������5�\�U<��X��dgi��&H�������d��Y���m��/�N�QD7�&.++��q	5�Ks�L���	��]�M-/9F;��%�5�)�Cüp�e��(]�O��(,��������o/?`(�(�R�?2z*����w@0���Y�����J����³���;��{H�;�e�D	��)��g��#f��!���)��I#���Pᘳ���ΰ��e��@��H"o�Ǌi�`�r��4/߻�D![H)�R����Gۅ�Ȝ�!�w�I���B����kD"��G�!����i"g��N?�����i�XNn�;X�%�-GU�m��ٮ(N�ST�	��ѿl������֙u��|^�Z�Gėkm�c��Ã�o(����K[����ۚ��,�lpk����Q�-��d�.�#�-��a7���ʉ����SC㒚�U�_���{��Qu�5��������H����ug�}�\����%��2�n�&wo�7���x�N��(� =�BU�~��d�A��"�g�JBO��@�uz�T���̥ԥ��G�b�ʷ��{�Eٜ�-^~>��G�����q"��Re��~�8ㆩ?s��}��^�l1T !����ST��ip[���'[K=i{|��`��0j�s�O�E��U��nmg�V�{�1C8����j`�M�M�1XL~�@ݾ���_�3����Q'��bƸ�p-z��܎��u���Y���4[�qH�%�w��/��|��V��?7��e�PyG-I�3b�IA0�Pr�`(�H�W,�`�C�"X�
VO�;v,��t�����Z�¹ӝ������Gҭ���H�2+��@w��vБI�����c�@)��y�[sj�)ls9�5<�5�
*�;����M��ZRK�x�)[��:���r�P��Z�i��P��f��;2M�����%I�iަ=��)z���v%&�$� �#5���n��{�c^��4aG�O���ʣ�?��~³3��m�1OM6�2IX��K���Jߗ�n�ZMo{���g+��>��L���)Jo���8/�"�u��ի�=pW�K͡9�������ʒ� v�S�r�JYj6�(�3[��V�ɖ ڮe&!qm�t���@��%Ó.�Ү���j��Z��䊺k�7�.�v�}ӛi�� U���gY�3�f:����"��ف���^��{>.py�E�F'J":��!!)��@�!�V����A������6��1���\k��2	��&�	WChD���~��aMa!לu���G��l���d��>�ӥQ����ĭ�x8"m���/�P�h�����_m$�f�(���[�9��G��(2�2�p��N�n���sIq�l�Z� ��_[�B��א2a��Zvr����]}�4�J�̙.#:㳖�J[�0\|��nޞ�{�iX�g݌��Ｖ nL�Q��[_Ż����~3�#4���ϟ?���_�Ϊ�販���~��-
&��\
���x�Y��|� ��ku�^{�"~T��i�3��!v�������񪑆al�lgh�܅S��+�����M�@�K�Q��3d� 6������N��#�ڇ�U��$�( ������$Ze�6ĂHUq'��7@����=�'�>�B'
���NHYzj�~�� O�U5��8:+"�$T������;*��G�<-_li�sE1~CM��,*C\�>��E��ۖ�q;>z�7}�[6B�� OŤF#����!��E���Z���~�g��}E89F=����!M���RO����bbb�a��\7�S��ҋ��"����?�D&)$�w�#��-��cg�)ȡ�m��J�Wj$<�=�/�e!��i��07�{I��5���(�׍�H����"`��m�+M�n�[B�&jUa��OtAbN����aO�+��{jb;"������9���h�"��E\	kji���ﷳ�M�b=Gl����2�����:�{]�>�S����}����J�� m����J����wR�Ӊ(J�9�9?��j��	O����(��u��#�:�+w�A*2�F�$4|��J�L�ue�_�3#2�'9jV��2���8�&�VUǪ�RE�Ms$�H���AS���+R�^=A�9A��=�G���s����c���k��H
xϯ�ׄ�4���������Z��̀����G�C2�s��9�oP�d���Z������~r5W�[�O@z	EFL����*I?wы�h�֗w��?�K? ��䞮Q6
pm"=�yZ@U�������6H��R=�)�@%#*��;P�En��W@>
\��]����I���U	����K��.]����e?<��cί�)��(˘5������Z[�Yt*ކ�O��W����e
�����[�8��v���2��-���r���XS���_Oa�\�	�B�j�������&�{�(s�:��~Ŗ[�{׽���wC���,�?�"���F�PN�83��Ƚ�>v#7�����Y��0ű�U��u�Gyr�ҍkĞ���}��K�`�`��E]@L��(EZ���m��ޑ颂��1�Tr�8#;��FKJyމQ�+p&�Kt�V��sKl���-;�䗰T�N�[��X�Ň��������D�Ҽ6���&��ʹ�]p�HEf]�!M��<�;�=-Go���"z=���R���L�O�ۤt�72��5��V�Г4���Ǆ���Z4/�{����X̤��o�"�.�j�k�<&G�bc����1Ҧ�ZF�4;s9[����&A���x�y����w����%Z@�Dr8��F��F��X�1���pw}7JR��g�k�ӪIa4D�&�&��װ��1�{xc��NR`d���"	&��HBD?N��&�l1�0�g�r@��Țj����������H��'�u!x��^av�H$e�`j����{��i�t���w��p���?�=�ii"j�ǻ���Mnu�M�j�Z����~���2E^ *�|���m���]����@�jE��Ex�/7��K-A�W���MoX:�9�1��a)����6���o3�m�<�#��ݮ��,��ߜ�~��Q�:�sG�9͉ ��k���Fs�>TX+8��հ����+�6�]*�!�tk�Q���L��ST��T�+�6>1D��X�e�b�܇��k)L�
o��C���ST[�� _xj�%�o_��V藀;���/͕/���}�������+����3�3Y�F���ͻ!��" �ߚ~���}ONr�6X<6�kkvQ�GȉD�4�3wv=`-^�L�����w��ڰZ�������ܣyZ�gPJ�\x�9��ҋ	��b�bl�o�Ŝ�|�P���<���-m��@��b֢�:I�Q��42�����֪62�2f��1 ����8+*LZ�<�ۑ�!Nq�\�H�6M�u�\��	�{V�c�n�P�p'p��x���ܭk�T�c��ƹ]ϩ?$��aQ����L,��q�Oa���O�wX�梁mHqy�(�)-���WAt��2{���5q��7�I���f��n�!����VL�K�'�`2����k�K$	����������Q�r�C��N1i�T�������?:�ނ��k�>�f6*����'������d��X4z��'Yx��\}����W<
�5���V�S��0�e��_���L���z�a�PN�CA�K���YQ��T	��D�/ˬa?���� ����p ��a�ˌ��}���@j���ߥEV�K>��5$�t@�kv�B��="�H��[	���@&�8�i)"6D&�gt
�E�q���/�kCd8�v��B�B�).�r�\�鶨���q [���f-�9_�ȒA�\sb.�aH�N��o�E��p��#'��l�!�Aݦ��w{���{�Y�3���rW��Wj=EI|���Z~/�_�߾�W׮��Ѹ�ͳ+����J�e�j���cXcӍ�g-;q6&�L,1V1;��H5�q������ͬ���F�y�����47���v��b��-k]�m|�f�heӭ��r�"�]B���nGx`��U���7�H�p�[s��^�|&0�:���굞��Ñi��A6O����-���(S���:����\�:��1Bs&�_���� ��[#V�7�:���7��LPi�h������}�+��$˒}q�{~�n�3���Z\%S�=i&U�݁/��T�.�.ݔQ.U.�!?ɿG11h����Sy���內�l����$���� NXDa�E?�&�fn}�y��_������؅�縱�k񘐭9�O�)�w�%����ȴ�g�'��X�9AV_6_��ؒ�g��+�0��8 SGq�q�Of����#����m�l��wI�����1#�To-?�A����Ƶ�p����+"��@�B��@oH?u~�:�"藹���h�5�:@Ƌ���d�_��� � �N��-�u��`)�UL~u"���c��1?#�Y}C�>�\uKI|\��Xx?��<�D�D2�v����H��h����Rk��sQ�V>�&�R$��E�g�������r��D�F�7��a�՘ �6���x2��c�{[k���p��Q�݅����c�OX��ND���X�0`�Mss���o0�d�J{�j����j�=�*:�ȏ�2���K<"Ga6�JD�>y�rAߛ�7W=��Q(�3�395%�1J1,k$4U�q����Oh�3�e?�zR�r�q"-�|�ύ������Լz�t�����/*�m���;Y�o��Y^�&Nr�Y���! {�"J-���� �VZ�p�vD4��mp�o_����A����խ�{�7y�ٴk���)ccs�+�g�)M1��x{�Wu�/L�zQ�S]A�5�`qԴY�/ȭ�j�^��L�cfʇ��x�hZ�"K/���Pipl���'�O�Fås��������� �)n���$>�W8���ۧ�j+��ƾ/�|#�3l�H���U�	��?d<���TnX�(M�������Q1�?���@���rD�&�9��	�1���p�4p5����Z8Fbp9�Ly�9%$�6�?��,'��Y��o�+���mGK?E����b��ɭ�u�����:���gJ��`$��1��!2T�|�=�7�қ���N{�T\�]-��\�O0+�x���u����r������U	� ��s)+a6���=���9�!9�������}5�CNG\�S:��~_�
�0~���;���t�<��_����!��<N�J�oK�z���zy�w�#��L������P	Ċ���TB��g��m�f�fz����y�R�WŽ,��@�}���@��������E���4@ǻ5��p}q�{ӽث_؂YlWܟ5�s���wv���\5�����OG�8ˆ؂��{��׋�/�ђm�"�����T�H�p�.��j����Xb�áR0�㔯T��-�'�S���B�p9��~��5b�(0$�*�I�لxt�1k���������a#\IEŧ�wB��S3��2�`MP���T�	@�w=��i�	�xz���dݤ���e�C�>��	a��LQd����0�鵏J����#��9�hw�(���ܮ��ڷ�6� Ne�(�՛�dBr"{���bz���/��Б�V����	�(��n�F�f<�s��u߳�gb�����R��=��ty�:��fK��R����F�O,VX,���'�Yƭj�'�,��kszk_�OD*K�<T7��;>���53����A�p��,�9Vb��1�Y�`:M �?o�X��2vf�;װ�LKto�*]�0e�q�`j�{������R�֮~�>㇑�J�[�&���'���H�eb�b7�����I5ou0�i��i_P;�N<ͷ���>l}��!̋�p��(F|�d ݶ�r���!W�+?���<����m	�c�ݸC��d�!m7?��4�^�E�  Z�}e@��4������Ns��_�0%�䮇9�����
1�G�侬���3ET�#�A�4�b�?�t�����{M3��',=n9������͡�C�c��_���e�N��8���2<c	�j������R����k�_x�\ƍYG��t�B���l��gN��~Q�� �	Va�����,��H�k
>��}U���z(M��ٰؤ�π_�������Fą�;�(�\�-��F�i
eg��2U����<UB���.(ۜ�Ɗ2��)d܌\�/��Ʃ�?*H���Sc?�۬#�ÎEDc��Qɭ��?)	qT&L��r���|T��l���	���j�D�=�_p�cŖ3��d17d�j�S;j��9�.ᘁRs��3��˫c��f1�6�����~�ϵZ��2��4#�j�T�Tu(7"v��;��O>�>��لշ��J��[C��f��5?�{9�dI1X���~��7�.r؈lXm�H�\,|	F��&J�P�����NV�ei�TH�S�&_E���qtv���9� ;`��K?��qg����gr1Ѧ��׀������z�1�dW�4��Y����ʧQ5�چ�ى��u���Y�^|�O�u��}�Ȟ�'6B�}#K�
�If����~���I���ג$��j VMFR#h.��7+�5�ꉦ���W?�GMGkC�jx@�n�� ��yOj��(1ua�̸�\��tt��~v�~;�J�#�L��.T���j2��ٌ��ع���(|V���G��6l<���l��=Ό�S�8�{t����NM[]T���m�L4�@��#2V�D_�E�tg���&3��d;2��DP���ȕ�i�䬫�9 �k��Kn겫�7��9��N��ح8h� �v��)c���kH��*K~��K�f容=w8�o��4pg7C�+?�):��Zٍv��a;" ��gԋBQԲ�q��6�"�g�&�X��K�'��c�#�m6"�*�9�M_G:7��g�8#�n��HOaܶN^W�_�/�ګa�/��	֡�pW���E�3=��p�7����>�I�U��Q{WJ�/E6����`���WQ����S/?���{�sZn�zYe����B�g�K$~�1�z�R�XdC���׉���R�*	r2�6R�;���~�m���F0��c���<�!��E�L�$�P-�W�ڬ����og�KA���@�W����g�Y����<��"e�ÙA%6���lꤿi�˯�fO41���F��P��nX����i��1yMc��^)�c�������%�/��g���~7�y(��hj�y8�Љl�k�2�[�{a�~��pvX4\��g]�cw�Rp�p���Ny�� �J���k(����Gd���F8C���3ѧ7���L�M������ѐ!W�Fu�;0e���%�J�Ը���G�#�I,��=Q�HA��ѢՒ�����_\�V�P ���a������<���%�\�]u��s�����ZDv�Uc�WMߤ������]���<�9÷o��~�<j�k�26��n�aiKk�l������g ���@ I1I��\r��!
3� ���T�9�l�|7���%d�	Z+ΚY����v�>����a"�g����P1��/�w:��啊W�
E�zfL�Vbo? ��6��ݲ@O.���A�%H�w�os��V��n�����@�`�R���R+6�5�N�G��@��v��Kd�Y�����V�e]l�Hh�֕E�wո�� �\��]G�~S�~���[�'������Y�<�C�S���*��111#�ݦ���W7�V����<v�����<�.���`U�v.�C�����	�j�����1�+��M�/�ؘ0�����,%М���F�o���f�dִ>ڰK�X��w�.��y��Q�q�;��D7^�����V��7�VV�5�-�M��������>#<�0d5�!�:�J�"�}�e>(�ܬFq�%�E��>��ը	{�l2d���Q��Q
8�7��W�nuf���uf��m�Q����TH�q{-��|���!�!W��O�B���χx�J������Wݐ"�W��T��h�g�P1*]���RU^]��`D�3</�z������l�[�2�1�τ0�I2����|���O::�,��ӝ���xf��V��D&�J=�81�� ��.�(Uէ�⡥�l;�&9���{���pq��,26$�é�~q:-��e`ZҐ��K$q>٬�K���x�p���]�N-,zo�8 \ ���&~j���쾿_/ɟ(3U�J�w[�G�!@.��yqe�Ƒ_-��G�@�����JJi�S��2�x����+\R���>{X��1O�s�'tn �B�
u�z�y��%�*0��}��E���JL��[fjI�[b���ʥ����_���f��C��z):��Bnnma-���x������B�2ʒ�[rQMol�g�p�sT��p;�YP����y�ԡ�>���m�YQ�O����n��Sy�V+p^2������[Sho'W�#��,��۹�8�e�>>���ͳ�Ep�mTf�G��*D���0fd�����v����i�,"�TT��JV4���g�- �<Z�nE�_r�W��F� C1�[���s�yn�#��4�]}�ډ�<Y#w*���nX�$��p[�3ާx��$+:}7��}�4�I�\#�2o�2=�~CF�H_��t��<s�?s�'�p/,(~�$g��ь�Y��xQ��hw���Z~E��ݜ�I��g;�/(# 3	�!�6���+ߔ���A���گ[��`߭�"1���<$ M(y)�<���q'f+_�[��$&����8o�ſ��+�H���|l��篂��I>�#����v�Lp�8��D��	���s�
|�u5ŧ��"?}X�u-􇅣:"���E�l&$�z�$��cz��Eܲ�gL���
N�m60]�<�n����bK ��+�G�SS?��N����`Z�X�M����?�H�!D+��}%'���K��%�L ӯ���qs���F�u��k�����������?�1�a@湚�ҼH%��퇦u�����C���Q�O/����F[%�r�����H�/ޑ���X,l��n?���׉o�9Վ���.F.2�ǯ�7G�ィ�i�n���*������,)�v���Qz����R�B�K-�����Q4��Z��t@��Nn!m��u�7��c����޸C��_ÿ��#�*���*�0�
�ҭ+0:�>ю�'��_��͊1MK�L䖭��f��xߩG��F�J�3f]��Xs<��%c��Y��x޶���N�������P�O�[�bg�GMZ��������K��8��r=?{Rr�j ø��u�-��Ÿ���ӣ�¦��/���=�cU47:_8��^.��p?#(������f.�h1Fc��_��%H���woч4�c�ʿ���NNEw��y�c.�:B}=f��r�c�ϗd���k�"V�p��c������L����Wz ?x�<犫0TsW���.���5J�Q���3�&9G����7o-+#�g����L8V\�lS��q/`:'���
�Q�u�uD`��Ӥ���啵p<VV#>��i�2-��$v�IQ�Awk��h���Ѝ�ͮ	����_ѕ��d�pE7k���D!��2#�R�İ8��c��]C�~0-u�`<�̧1�Y���6�Z��F�Ƹ�9��Rr�D�xh����z��v	b�\K]�￭E��?Ţ��*kN_�1E�u??~ĥa�{/?H,��g�N��PLR��'�g�[�:Y~QR�/��	��x� Z4�iSo�GxS�����Xr:{���%�.��s\de�*$�0�`'����xj?tN:������fo�	�<F��� I��T	��!aԏ�_�<&1}O�&�zx���v88HHA��yJK�%��EΥ�+��t�1�o��t�[�F
��v���Y�Xe����:��a|n�c�� VR�t�������Ŭ�HkV1Ak���T���)�˓��Ò��q�m�sQ��J�J~�m���@�!:�E�=�A��C�hGxy�A �W^�SZq+ðoftO	��v���	q��}�a�n�"�Q��G:3���*���a|��N�����o�eJJJ,,,V5��i*�;�f�����n֬ZB���?KNr��
a�t�J���g8Yu�����3R|\G�ٕDȗ��C�����+�w�n��,Y����<L��r��H�9�#& ~�ydڹgd���Ż��@�6�:Жq+,�z����a��mQ�e�kn�_]�� �#gn��������s�GkDĈ��*�/*�h��� �VL���F�d�2 Oޭ� �,��1�1 ���@q��R��`A0``��11Ԉ�`��oE��C���S�$�F��;��x��`��t҇08ϥ̅�q���G?"j�;�S#_�!�O{���UH�s��$i�:��Hn���ɤx��&��B]R�q�����Q��Z�.9_!���Y����O��oύ���P��s,!>��j�m�5��qb+��6锭��c���JY��l6h��ǝ���YPo��.!�qPn,-��H���26j���J�_�xl�l�W�>���	ц���4�ز3P�(-F�pEy�ӛU-�P�����0@&gїX�`�a�p���v�@��v��p��*_a6:2�ضj��L��B�Rn�x��P����_�V@����b�'f��}�eL}��^�b$�"�kyC64��CB�c�8�y����.�z/i1u~i4�C�(?�P� ��MG�1'Z^�m2�`	���On�NU�OL��Ԥ��n:�wY#+���+��s#���l���n��d�}��$#�O�N>�GGnD�^I'�Qm$׌��ㄳI���d��-l3��Z��@��Т���� ���
�sY�K�S��Y�$�[�x����N,�-�����]�g����>���wɆ�{)}��'%��qϟ��6'�t�8��U�����F�� \\����U���6ֽ�[�}N�@�6���/��K�#�"�$�{�B�� P/���P�k�q>��{ڎ$3���':�,����<R��ޅd�D
�/zВ�!��?h'���`�E�5aJcy;6Ph�)��UcC�q��'Cmj��y�Nh�h��Z��o�#���O��c|w�����5`���[��Y_�:{ݧl�I�a���>�-y%Q�=}˸ԛ�}j����ϋLdBC�*;��<`��]Vc���- ���V�y�H@�1G��`��E�tZϓ1����!+���^^����C��>-0��� ��X��Q�M����Gv�Wۈt��9}�3Ҽ0H���40�qc��J~����?��l�?��h	!{�u�ȍޛ����+��PA����x�Օu�xy؊'}�K�/,\ܢ{���ʒ��{XX*j��6��b�0<�S�WZ�X�9^��{��b8�G���[��w,�@�� x^fh����	jx~x�)[|��H9-x%�XX䈃��xh� �	:`W3޶�$	!�~�g�M�٨�/�6A����ґ*�����A�0�c�8���-��
�0$Ž��>�/��o���dF��P
%x]�5�$�������"����Ll�H'��ι��k����9�F�7),wsp����?XэÕ'���P/*��ul����	�����2T��6��`]�����U��ɅR��t?�����k6m[H��א��`gF����m��-���6��[��U��I����po���p�dO\��ڥ�?�E�*�I����F��Z[k��q��~x�Ibo4��Hc����9_g�=_��b�`�E���
����^jG5D��J�@թ����B�%@2KB����T�E^}�����a�W3W��װ׀� �L������_<����Y4��؀��A���^\\?+���TC�)B�˫1��5��m�J�%�PC��דZ�e��s6$|���'Ȼ��L%Z�>�RM��I^J����Ǣ��K��a�A���Lzu�Dr!>
$�H�V��0ͤ��B�{�8����j~-���2�n�d#>���i��5�\#V����DGt����lURڑ(`L+,Se��1J1`ms�w��U
T3��D�g��kDu/�4B^\N��Zd_�́�_e7K��K�o�ޟ�<|i�hZ�u}�u�~t�6j΅�"d
���R����W���U_�r�"P���ݷy7Ԝ����aC��&��5#�'4���6�E��u������a��ĩߣG�����4�2�a��og� ������3J�7�xt(��h�E�-�`tж����$�a
"��9�' em�f��.1� �L��ܖ�b{�G	-�0}P�]�c��QrKT�ԕ�N��Ǭb��3�>$���n�.y5$^�wi�&�ɴ�:�����4s�F��kU�m�'�gRU�:D�l�G>�7��{������=ԐU�]!D�)�Ihe�dB� -����"O>˻Y�<��Mm&��O_������=��=�M�s�4g����Y��+h[�>^�ܝn�����TN��)��g޾\w�w�G/���@�������;�1��O��I�%�E�?��S�34@�160�]�a��L���a��`Dɏ5,�9K�PlWl�2X&i!i���7B0�"���_'Y�)�
F���_GX��hi�70KH�i2���?�ډ��H�?k�����p�å��¬�"��b��#ۇ�4�Wu��X�'�gkE��^q�t��& �I%H�b�+D"0&��S�x0�JJK�3����q��RƷ�h����+�(�(�hX���[�ʙ��~+-��~������co�pY+>Mq��������ZvȀ������琼ԥ5^��O�[.e��[�0:cW�h�)k���J����nMdw[�g�`L�L<��������g<*��k �'�SQ�+�N�d�~��^L�?p�
x��<�#lC�{]��\��$5��3$a'�ȓx}l�9;����~��ܷ/���pL�Q��������_���f�ϟ�ê��F9��p���aܣ��~zgØ'�[�t!P�"���@_�\X���o�T1�n��gܯ_6Ґ���_s������?8�&R��+�'�Qʪ�pRV��X]�"��o����-�D�m�Yֹ���X�G����U��~�n�x��!��u:Q.�D��ѷ�CCIF	���1ʂ*�Ç����b,�8F(�<��ø{(��x�^�a=1-o|",.ח���HJ��g�d��z�c�"�V�..�BR��2|%(���Z���u��vh�Y��@Z1l�K8|
46��� `P0 !�;�>�����LE����e�R5�V8�vd�|P?CrE��o�Y M8��֪���C��u�!Ag@�Ѱ]A�odm/��@4_j��'��	�_��ߞ5\�_�<[�X�r�V3�6A!�f{��W�H#��6h��(qs�"�dۍ���`�� {�s��_Q#�#.*�9��]�3�O5R[~��/u�q0�������G�m�14�����'x�=�z�^�3w�Ĉ,_t�֯w�+b����y�X�
�}�.�:L�L�z	���߇�@�6�������"c�cpiԟG�0ۨ��xw��J�5�ıy�@���<���~��%F�zK�R6��>41���R,{��hX2 'd�bB�
^�ʟ��n!r�����d�&)t9��[��}���ȕ�I�"	}�m�R+�O� ��ݲ<`jh�8���|�8M������|�����Nu�7-g����Q[���� ��i�ٷ�і�nF��p�s�7Z
Kɒ�yj��^03=s��$o���G6�.�.�տ��"������ʡ���~c2h���!��G��9�mlX]�_/�Ĭ����~�G�|���\�cS�.�2�b��cp�CI>�X�rX|����MyP��*A��%�����o�o�]ؠO��B��h�F_��P��$G9�R��ErB�;��4'� %�t�A�hEV����| �|j)i�a�k����2G�����ć���?�w3����I*DѴ�����7�+{�%�-u�uQz	M	������/�f9~����`R�k{Q�6��4���9�l�����@��ۺU+���OF�G*?m?c�]�JH����7�z�ir{��0m;��bdz�E�`?�j
g��*��_�ē�`!ڝ�����3t����0f�j�����9f�`6���7_p���B!��?C^0d��@���i�*B�I���h#5@?a�Ug)C����ԛ��t��YɞI���o'	X@���*S�I�<�,�NM"N�o|k f�_Ǽ�+�%2��cFi%�Mڳ�%I�H�f�e�HQ�i�՝������C�-�`3m���/+
[�/ �l���
%����L�J�4c�y��>�>X�j���&%ǒ!>^��/����fI�Ɠ��r��2�q�mZ��
��ٰ?�Ӡ7�Gyr����I�!#0:����w3a��v൛o���������p�5U�}�&���Q�7βFbrX���ى?%��?�$�ߎ���(��n.G�ʋ�8�B��N��?N$�G��.V��K�f�ц��{��O�<OB�p���i g�΢0G�Ɓ�ޣ]��.�xڲf4���DG�AU�;bA&+ss����.���䬫��xZ�	)@��F��ϣP+���v�vܪ�G&/�/��˻/ņ�]�ϕ���l���}?Q���o���,�t���1�G�Pҷ�t����K]�ߛp[�;b�a�N{k�ƴ�d:�!��)I'�4���KͨN@AV�"]TK2�1�g��%���@��d��2�E�Y�@����
�ǲ�
�|p�{��pg����%�v�����p+ ���L�FfG�.����y]=%	- Ox���ZJ)-�� �2D�~�|�!�sҖx]�8���
�w����d�2���()e��t�W�RҮ�M�f�p2���d�ͧKà���EB�f���Jn��a��J�o��!���v����j�3�̻�01�͵��ݗ��U���Q�_��\}����Y�ף��/c�.��F�Ŗ�'C=9��G�y���~W��ҍ˹f�%[�S��9��1T�i��u��������FZT.�.R�{u�u� s@.W�a����� n	H�ݜ��IK��n�Cgc�o0��#�g�32����Q"��@�3}b����IL
2��"E9t?��B���������# ?\3�l��u\;�d�L�Bl��pag�V7da�-p�cț�J��}GH��:�۫6$��b�:�Χ猟�q���y�~�Bv��SUA����j�7�Q�*KՋ0��,�ȶ1zb{\��i�? �?c`Dفv����M��%��V�>�3�*=�/�h����,m��ߧ@�_����6yE�����������'!���
��#�;�h�CrW��x�cB%g|b���́.��y�I���"uް)K�;%���)��wA���e�WV%��>�
�C�X���C��)ό88.g�=�t�u{C���Wy�w=��l�� 
	��:4Y��ﾾco�KkQ�:�(�����	fki����i�'`��������O^��l��'`c� 䪆�y�|��_\X<��,�{u���������/w�"(#@�R�҉ M6����Ij%A�7Su��fg��gJ�ފ�o��>�!j�1,I"��̠i9�Y$>����9��~{��VTII����>y�>{�B�T#�@����\M�ߺ&S�(h��^�SH�����Y(eˈO*���vg͵��*�����S�k�����ʝ+ؔ�{+�`��?�+>�5�+�$��Е�LHzҦ�.(GY$����	b <�Ȧ�`��H���ȗ�7,򯅙��3>0�0�^��ß���s�����)/���6��L�����ymN�zL��#£[Sn2ZʾHT��b�p7��n]���I��UO���\�ӧ��k$"
j]�_��}|�E�d��7Wm�%xj3��(&J	��&2�M��@��̲�%@&_6�o$ȾD�$��� ��J&�( *4��FP��|=�ʻ��c�}y���B»��� �Y�=���F���us�ά�n��YÕ��S[�ʐ��g3RU����&�bo���X�\Mx#߼���q�T��1�!��������Q���Ə{B���c!���Vb�mm>���R�JnE�/�K"�M q��E��7u����/�.���V�:q���%/CŠ����ΐ)s�5��[R���4C�3�BT���4+��}�_��d�̘Ѽ�}Y}J{k4��&�M�ċ,bQI0������M拦�9.�CU}��[�:����ߝ񘼕���#���� i��ӳKϊV����uK�#���i���SMb�@��͆Ŗ#�{�㻽���֪���$�L�������_/�s�����km ���ӄ�2v=�M5�gE�y�	�"_���|�ڛima]��:A���7~)�i�%���/E�L��9O,W�����~��7w�5.�`s\��Q:���]팊i�6�����bHW�V�b�F)����S��G�L�C\���o5i"����ÑΔ[���Ư>E[Eܖ�p:\���x�{�=����O'��n�C"�;H�7)�����|�9H��
���`}c����YM�2� s���3�+\4!�KnMI�aH�(�8T+:R��h:�8�f���!Xpw�`�5���Cpwww	�]��C�ܝ����M�*@�]��>����]'Q? (�/.E<���ӖӸ>o�L-^NsO_KT���>�lԜ�mlfW�����{��eE7$6L��_b�{ �9�5.��;ËNj�����p��a1����|N'���@1�+�Ę+�.FE�N���<���p_AE�=�̒�/�Z;����������<$��L�qG��@��:��vdt'���������`Ycvve�0QcAĺ(�B���j+n^���IOcFa�h��vR� ��U���pWn[ո.iklB>F��3��5&��b�]���A��>�y]��?l�4�M�:�9rV�EI�ΎL.�,N+��[G�N]��S-)���d�]��	q��){�,�K�{�����BL� ~���l¥���(��6GL��g��=b�v��.?W4����¬�'K�)�	���4�\��h�]�RA?"����N���И<f�LZ_Df��@�����l�C~]y��8�xt�pT{ʄ���m��^�1I3��-�h0�ܻ��?��
�^���0�6|l��{ڹ���lϵϺ��+�!o{�u]�'c��'^?!�c�-�PW�����ߚ�kD���i�<I2s�"�`�/a��-�v���������ohD81���g
I"3���������fC��-�!�?�U%QT9i�ax}N`m�^XUՒ߽���),ڂ�����{P#���7��&�q>�wI�N������ I���zv�ǩ"�\Dᮜ��X��r8��2e�S�v��O�GvQ޷Q(�>��;�9������0��L2Y#pหD��RǮq��i?��Ç5A����ҨϬ�Uհ"����bHNQ��z(�gI���P2��:	!9K.h����\aLti�cNT���۬�twWb��m��Ӡzr���S�Y�ux88|�M�N� ���9�9fz7l���i8|2�zB!C<NV�s0x+��@��OJG�?q�kMw=>Dӆ��gj�.�� ������*9"�̞\E��oU;A�����j��Fՙ]�x��Hf��<��۸�e�jt R��SB����M�|E��m��l��8��ӿ��S���� e��K��񶜸�u$����$lQ$\� �F����+ܠ�"�sW�5�uG]E�7�@\m�S�M�y������vh6�II-�q�	�ݏ��6S���6��^��H +�G,\���2�=H�� ty�����[͗Z���,���Я�=L�ſC[\��Dh��}1�Ă���>Ϳ��v޴%�mii�c+G*i���`�� ݔ��7�����*��4Nd��!x�+$-D�� Te���p��:Sg�ܗ�~�-�����yjEDb3b#�����p����b߶d��:5��i�rZ���7&��м*jj��uzl�'#�k�6�)	*�{�2"��Wۥ�#Y{U'T�*!����n�{�����2g�e>	�������p9��+J������@;�mJc��'�K HF�+�|*��@=�I�]��0��@�J����_&x�A�00�+�5#rW<�o>PPPN�C5{K]���8a&z��5X8;��AmS��qm_�qt`�#�uI*�J��<3ć���.���}3�;ib�'�j����TqVf�;��W���@�������~�[���<q\#��l14�{��DW���a����x�p��w�F�BPFe��P���c�
ʓ�����f��Sw�сBPCfq���h'��4�`���7�f�hЋ���E>��H��������숅_G��$�+eإ�����O"a�Bh�L+%��B�(�m���j���΁�-�&�a4��F�g0���O6]�>�\!���9�*���/x�f�g�+4�\y�����_�{h�zc�ok�ې�� ������+)����[��M�P��~-�f�2����j�5,�(�Ekl��uJr�咿e�6�T�T�fΠ:#��M���±f�puʴ|GM�I�����SteI�<�����@N�B�b�6zY��{(<���ujr_�o0��?��y+�����5�}c -x�=�,�P42[=��Ҧ~�ՔA#<�A8\\�	�:�
959̙�Z��m����9X�����Q�_	�D;t縻7(���+SU��cPP�[�+2H�I^�>���j���^�@�]���&$�JN��]�(����5��t�=P:��&�h���J��PW�T����
>`��xo��%9C�fģN#{��aH�� L
��<��a�8+ST՛ձ�:,%�S���B����arn�N*��Q�y�zt��˥��l���P�jF�#����Ч����-�%�UF����(4��c������<�Bۈ�2"��wᗞ�xD0�H�OV��C�S^��w׋�ol�7�>���%U�����p���=�UuS�d�7l��)n�W��S�q���i(�Xl��������G�X�ᆳ���X�2�[�m���^L���<�}��]w�S����Rik5���� �,����$h���h�OG����WRi�w���ȉ#N�LY3v��'|�*L׭�N&3�e~�����m+���)^H�5*L�i(V0Z�B�X\kk���$�"2:Z��!�Ů�R+�u"4�������F��l���t�Z����o�q�t4.����b�B�������\���U�Z���4Y��y�s��R'4TO����RDF�󚹸I��S�d���3F�6q�3/P��@���ݛe͝}8�8*���a!�a�Z҄����5=֩�f�pv ��q����xQ�/��L���|�c]��,�4��������Xu���	-��������;p9�����?uR�w�w�mk7���m�WUATJ�Ƿ�/����pd��:��KN��«�b�Kd��T"�9���Q(�Ic���TIc3��j+>פ'�����B�6�Y"P4>���,��)�⹙��~"�7��I��Y���vzٷ<�8W�t�r��z?�$/��,��ٞ��������G��*���q�`���� �$���l��Hޫ�(�?N�<�|~�5�䎅�ݲ�fN���d7�zF��%r�x�z1�D�φ�Oc��&�[�_�>�5�[����cMNq5��X��7wF A����U�)�3wۣ��㥙����(YX�����Գ5Te�d�Fq�ӎ�'�+�-M'`�j�@��;\��w�+.�OWnB�V=��]h1Z�Փ�|+W��j��<�"����
�����m�}�%[��zq=�\9����pN\p
V��+��̆�����x�G8���?��������?�#���1�OY]�����	��Q;hVvCG�y��ʔ7L��q�Q֖ �N�ۻ���+s�S0(���@�*���]Jt��S�"?���ߘ>��^>zJ��@�,����K6pd��Pr����%��@ԫ^�)��B�M�g��V��ʹ���>z�J���N����ӥ��S�6�Q7���ѽ�.@ z �O�� �~ѝ�X��X�raG@���`��|j��TS�������x��?����
�#�7Y�P'�g�aa���u�4�p �QHo��U��ŋ�
�n{�A� lGi���1'U@h��:}If���P#m��aOUfY�[��l�;�e�K���A�ʫI�( Y���d,�m��𯑻��B�P0��ɨ�Z��*��{�������}}����Nl��!��f���U�%���ׇ�����lɧ�=ǳ�N�_o]N*98���Bn]L��H;�	�'����S��y��	�
��[�#�*+�ߒ\�~��m�FE�eYz�l?d����S��}XScK���"�,n��Q3ؽ������������7z=M=v��	�d�` ��6eI_H�:���DnC)`Im�q�5U����*��� l8�au�8I�`5FuCހ7>���¡.���'A�pe!�=�@F�/�n�2�ڗ.�!�����LR����N��sٓ�[�Ө� �Z���M�i�^����ӟ����_Ŧ��`�|I���e���K��oI#�:���,Q|�9n׷���E�8��"�J(��O��D���@�Y�����D<�����*��y�1٭�V�r�X,��s�!�)��.����� ��]����oq�a�	iV��XN�<�4S�f�Ԭ2l����>�fZw!W��H!L;���WZW��19,��íxqf�Sɍ�(~B��*�ѼlC� 6%>z�0˫b���@��q����?G�(��T���Bu��\/ۻא��꼮Xj>8�6C�\�o������G���0�O_ �t�<�1=�vgs����_ԪV%o��Z�S4ڷ����V8�* ��ڻvH�'�yxn�������.�/�bR��
_���3�����������o�^��|���;�?���>��yL��FIZ9V��[RY���a��<ꔺ��2��ȌD�����E�����S�bi�4!ǭ( ���yʗ������S ��`Hu�ђ�/���OY(�Ǔ�K�a���ÝC2�Ȩ�� �:ޖ�WfZ&b����|�؛��^�3z����
n�>W?�#��pR��_:ǎ>S�3kQ	�4�1�!���`�axl�e�)�Ӄ#sq}w�s�1c�o 
N���,����@��j^-��o]X_�H�|oZ�x+�����)=*B=�_R��21P.���D7Eg���b��W�L`͆W?hE)���R�^6\��;ýھt�9����tn��79�vEy�u�e	��=� �{ݙł*��hv��ҧs�����>��~�l9AZ�%c�6B��w�?=빃�.~�I=���`B`�W�pm�4�AA܅(�>�{��O>�����be�v��r�aj�*p�����FK `��Y<�;�sg��H6	�0F��{T�@�Z$ �������8����	�z?����d��'#����>�{������p��̉B�G�}�IF���Y�a�7�~�����[opL7���zI��7�BpMA��6���7.|=�0�P��ʇiPe���KFoow4���Y�0@t�Oŕa���a����m�`�x^�~�Z�40�AeF����t�^�����\^<C#-b/�~<7��ت(�$N���w��T1n�=B�uw�1���ßJ�t�
�
1Ų (7N�����7.��ĳd­Fx��ٙ{.Z�N����R+B�T�lA��v+�PA�5�_1��Jb�?4)g1MO9@1L!eR,|�4$6<6ږ����.b�L�J|��j�=QL����?���;z8]����{K��@ao���~��{n�G���~�Ұ�(<U����h�n��@�� W�D�Ub��eF}���f��.S~��^�>mv��W�:[e��zEk%�^^>5�aI5L}� OQY9���~��`��]�"����F&J���hC��69�.>''f|\&���|=�,���ʊ��p�>//�ŒU�>�'+z�a�r�����d�D��ʥ����Ov`pg����Qm���� Q��pj���4=\��C��
,F28*꓋���E߁SBb"���뵦�_BR7Fckܬr�����Is��O�e��������*��71�>��f�9��_����D'e$]���Omӏc�Y�:�����W��:Jɺ72Rd���(�}{��k�N:;Hy�e�P1�$+֓����c1��*���:s�?㿚(���W�k��h++4�ːe�!�!��*[<���-�x�*��G�uJUx�&o? B�h��/�UAK�h�z����f��)��(5x̴0��g����ä���>�'� �&B^ޔ��X��bIz��D�P�	�n��W+w6i�V܀7�sF�f��z���g�+?�(s�������q�	���q��{��͂�ֶ<O��{�ė_�c���	�;\�v�vNSJô�m��wrVt���D!5#������EZ�Ѿ�*���*�I���S��80}���-/%�E��K�\$F�S}�F����O�ց��jaN`�$~*��L����_�pw"�jD���>Wk[LXM�f�b�۟�i�"�rK�9�omu���#��qs��h5Amo�+�֨���кL"eӫwA��w������C�7hln���O�����I�F�Z;�L�������a��T8�tGO���N���f�}V@�;(�Z!V5P��б?��M����!�3�eɀ��{�7GV�6+ k#�qd{?�a6��0��t&c��'�@e�s�W���W�����ԯ����a�t�_��J�Ψ=�'��t���Rd��T?q㾺�#�Sq���"�8���9��sD�a�<���N��rw��P���0��+�.�����)���3�1x`�J�L�x��װ���B��f@/�����k�n�7��G
;�.�4�h��HAF_��;�vz(|�az>�o�,��sig���1 j�;֌D@���}����o}^KFiǞ����ULIFQ��r"N���`r%�8H���?t>7'���)˥���i�~���Qe(Ɣk�M��C305T_�a��LB�j?��C���l_[����q��Ρ����)Q64 �����A����¢��4��`���N�U��z���m���RD.��	b[ֿ�}����u=K,����L/��[]��Nm���sf*`kKd4�ҿS1�˗k3�ظ	���vt���7AoLn�i��Y ��2������L{���B&�5�X%�������-B[��H���C%���ٜv��/�o�_uO;A`�����=zF�(��v��=d�3��W���!�t�%:�����&o�����E������$������,��[�����Re(�uR�W��m�<��!���ADA��E%���a���U�Y��[{v���� [�W�D�IOʋk;�G��T2�:�� �S��$a]�da�	��z�{��d���A���ӉR0���?���r���  V#S|��+�e����bۅ���,nC03�Q�У��(�~��:tE|�k�I��zJd�6�Tm�Q�@]u��WScXmm]T�;��Ɲ⃰z�:3;�#4�D<�.H��ϑ	�j���Pre���ꯑB/�d'��3��P��߯���c���[傉�\�w��D�mA=OɁ��-��E�V��-h� �2���+Pw�|Jt����P�.jkde���r͟,7��Z��аgz����-�ʻ�]��� ���'e�u������|h��E���b���e��O)�r���:�LF9%o��й	�g���W<����L�=!xxL�r��~2` P��xn/�S3f�T��_B�U��I�K��u�y�S�M��rH�/�>c��<үloC�8[*�x�hH��zn8��in@j�x���t_��:�k�w�~���ArF��e��f4���H����5�*��cZ~pVC��^	���4��y ɕi?IK�ԭ�(�_�=AԦ���z�¥��xvi��ƝIs�	��0�M��p)������e00�t�|=����IW�y��
Ry����P�@��%�36���A��mL���;W3s�`XpP�V���r�BH�4k�r�ܦ��ɧ���oC�xh�D&��e�|��\aXv���A������P��5�Q �2;��]m��|�?�g�Z��x�|F#���o�śC��R�
z��%~% 0��nW�!Q�T[��ÏPmN���t���o�����Qw������󹴊�B���`~��:���0���!3��Q��:.|���& ,�N��T.Չ��'Tr����@����"ArY�)��+���Cb� �x:Zb���`�C������4L�;P�A'���2�x|_}k�IzB^C��0@'���=��=��I���+K����U�i�aELq{N���݀s��D�No��<�f5���� �E�	Ԕe�1f�O~b� 
ZH���}����J����Q�C"\Շ��5���H>A 
X��Wx΀��������}�r�D��
ū���(����β�,4���\79�
��w{�rB몒i�g���x���fbb�;6_\gR����{���Ҷ�S��w��ؔ�	H/
��ރ���i'�ԹM��?����4���` ��_~o�ޙ���ѡȤ��Ԩ)c�MX���j�vj�0Kv�I��	�q�C{_�+V2ց�t�z�{��r����LW*}O��F������b�P�Y:���vv�1����]�\0e�פ���?Ay@��_��zo�VX��,(tɗ�a�8Mw{"�a����P��_M5���l9ȭ�F�
��\?�'�/�g�^�P�PS4scUU�2NK�l8aj`%��s���k.��K��K37p/7�uņ��e����o�AEp8"��C�2�zDUo�)�۝UA�� K����ƙ�I�[��8o:�#�-I��&_v�u���|6r�<���tu~Ç(ȉ�sʻ��׳���Z��ٖ�f0�@4����L�_c�髆f9�`�i5�:�[�>���ڰ��i&��)�B�m�Z3RkUc�à	!kAw�>5ѫ�g}�"��1I����������T/�4eFV�ԍa\:�>Q*P��(J� ��@l�=��ךK��Ҽ���<-c�@�b,99yg���b���ťw�!>++*1q��s���# �6S��5 C�%.�<%��n�>+��;lX�� IQ�w3:�k��ػ�n��r����R2hM�K�@�JH�Z��x����ۭ0F�8[v.�X��)�Rk�!2 ��G�zSqd��`��	V�D��1j����餜t�"���Մ�i�8
(|�u�vbOE$@q��ÁMin���ar��,O���z����3�o5�^`��^\����@���\�L�-�����vT7_*A�����9�FX-\�'UY}��j���)��K�Ǣ����A� ���4�̘A��_�)G�`�öFF}�k1��ӛDɎ[�	x���W�PA-�_��v�����&!�|$At����K��3�#�W�R�:���eBf.��o��|_y�Z��D{����Q?�?��H�ix�,:���m����)�`c�d[RI����Y[�'�%���"���@�0�ҖR��_��]�(x�O[�wƃb?c`s.G�[����p�, Fp��}k�֠HϖĨ�F���؜�\����^��c��[�.��N$�5�娷~Yk�ٚ��}����y*س�k���S��!�G����� �>Xèp{f�%���`:P�jZ�9�����rHD�%����H;���kx�\ˡ�m
�})���E4[���m��LTL7���0���A��#`��ю��#D�@��*ö@�=��v� �	��g�Y�)9�y�clk�p�A�y��'�\q�ͷ4��#{�o�����,��+�4p5���pi봆�e���܅Ԗ艭���p /��u�b ��f(]4��Ɂ_����$ǈ!k�8���cTc�*\i)@N�\G�Ⱥ_���+�,p"�"�6��0TI���֠��%�:��Hw�/�f1��[�h��]�eh����*v�$X5�::���K�3��L�(��%�
�UB��8����%�!ɒFWpZP�}�y����G�ғ~�Lr�PQQ��_ɇ�-���B�تYe��1��ft'��K#��f��r��Ҋ�����-q̎��}!��%�	���A�<��-O�HKK�jdx��+�$&����0�^������	F=~/�o�t��|�X�Re�l��_�!v��%�f+,���;��ң�\'�������,�y�)�l�X'��9�&������Ȫ��N�:����Hs��ÑN��+��ȞĶ�YM�˱�	"�	�2���4�;<S���(G���aZ�?U[��>�$��?�:���P%O�)g5�H@�R����T���:��C�za�,G�wg3CݟZ��a�9+����s�^�u走R�r�&��a��b^v�a�mR����s�[ه�'�{tv�
�]<�y�= �i�p�m� %ݥ��8�:�;�zi0����g_�1U�k�z��8�}��n��ȴ~Lk�)���g�1�𙎔�:�Z�WW��l�,��2:���y���Z��P��L��T��c����_��+ua%V433R�"�+)������Gu�#��3�K��L�%}G�^W���}�p=+XE �u�w�M����dC�Wj�6�W��>�`42�ᛐ��c��oIi^�+u��o�J���VZ�B��׆��PQ404"�MS�w{o W�lZexY�N�$p�d#ܶez����-�Nz����|�w���ﬣ�K��cJ'!aw��k� :��%x�yH�WYM4� ҦwvT���ރ�!ab��2��`[Y�Vf��C�T���aZ~�J�R>��)՜ue��ϔ��&�1���ξ���޼�>n�y��s��@ŀ�
F�A_Y�ZM~���|��s���w�@��,m�Hl��Q�?�T��<�7)`�p��J���(]VVE�n��)�A���OZe���d?h�i��$�2ځ8	-���x�
@V���7{�BGG�[��X��Pzg
<�x���a�A�+�N�A�8]�	'�^�S�N�.���D��_�Ք�����iO~ٞ�0)�2!Of�֡ݵ��a�u:�R��v���a���nV�$��O?!��(���%�&��Jxp:֤�Ȯ�_3��i!8�S%
Ac��/�g+�=Z��"���{?������s4�������0�^��ȑp�ƶ)sE_��w��*O��@u��5�D�ᕴ��Ԏu(~_G����[�V��Z��U�֎>Uµ�x2$c���o�ρ�+�j�KO�`4�!G���=���xk���#���%������)�ԋ�����5C?�m�9��3<��ޮ�u>07I3����THˈ�Az�����</~|l�eJ�Y�9��������Y����@�GH�(`�$-Ce�S���q�qXs�2���c*�
�Mp~���|��f�?��R:B�p�P�:�ԏ�e�� ���|�}Ay��Ӳ��bx2T���'�I/@os�S�/\򧨑��Vs��'��O�>�$@Y'�����2����^�ŞC�+���ڦ�B��&�ޕ(P�<���k��^qA�Jd�2H���,����0�����5~
J#e��n�މ״�x�\�c� V�h]YX�zZm�~��@�uuڎ������)�dǋ>
������{~��6�MП��k�\�PL
 ~�M^{WZ��:C&G��0!	�+�O�0?'~�:��V���sX�Ia�5+ЖaJ��Ֆu���.6�?K�%��||))���@T�;>��b;t�H��{�!��F:{��o���R���{4���o"Q5|^ד��}���Yz��Xw!���\� ^����z�:J7!j�E�8�xYq�4��\�xu5SjEQW�eLVB=}�K�¥D;Ղ$�\i�Wۋ�YxK�����@�i��#]���<���|_w�I����2#�joWD1c|=y	R�O�б!$b8/�@�uhga5F�#Ѱϋ�L��bc{���;Y~�]_d��v���CZ��تhs֊���y���bC�3re���k��<q��f��NL�q{O�x��<<%���kt�:�z��N�ʚUG���t�*��.K8��7��+e~7cd�`��P�t���chg`�����iz�pX�( B�WU&B�Dn��?7+L��$@��l�����w�ga��p�q�������sҷ���`'Y>�Ql���»�%V�T��$�ޜ|�qĶ8>6do�iS�Y{��gГ!�p#*`���|�B��}�s�X3�2�7��~��<��{�34!�v<,��.++���������;����g��m�h�<
�7�/��p���OC����טּ0���}G�Q��4Uff���R��/������ݐs�ݯk�~%�Ŏ�0��"�����C���r��p���9���p&�D�+�c�]1�)��O��������m�jʾ�TEsR�{��h��JE1���>�k��k8��r��)[���
�1h��$� ��wJ"���_}����kj�^7����8H��u���GB�^a1��%�}WW$����J!��c����R�o%�tR�g��k8`���t�y0���dL8����W	Ͳ*�
x����<���_<�<�G%��ʞ���j؆?7W�=��j�Y� ��3��M�C�Qtt�w1�j�*�ŝ��6Y�%�3�#`�I��������>۟Y�T_��Ć��(�@�zU���o��>6�]D���*�^m@J�N�@3c^���ꎆ��H1��[_K���z<�ѿHSH~	)H����#���c���~�l�.��_�ؿ<'���(��g?���Sd�U����l��C��;��~�N뿐���W=��8���W$]�F��F��KP.-���< � �2*��4�٭�������H�K��IĆ���o���3Ĺ�
UuիF[�'

+Ɏޡ@�Y_k�ENR���A�D%l�]즃�J���+�?!K]�}|�]�r_å19�+`]j>�b�19<�mAV�`9��T�[�؇؛�� VIM��ͭ-��^��o�}����d���dP|�tR@���^�j_�
�.y`�l�GH�&i|o�+��5Ml7/����s�]��c�q6��ǽ=��qc�����W\��;�q����PN�a�9<~�����/�*bg�z�[�re��?g�������t����^V�e�4��Z�P�����*�?��&�~��Es�d�m�8��MABM�T���J>t�d�Y������w���yQ��&��jL@�ίٰ����jH5\�J�\������2�W�����o��v��;ep�# 	�z$SiAX��	V#b#ab�&���kgk��<�M���CL8	Z[Q�c����]�H�����x?B�cDw��K2D<(�]_~���6�:3��
��M�H�����0w�)�G�M�Ç� ������<:n�;��vy.Z�9�Ilʕ�tk�����
����H'L�i�|���)��W^�!�&�&��}p[|Dwņ4�S��A�{��/�KA�'v1�!-Sk��yn�����??@4J��J@NS5�!2���D�L�q]�Z}����3�s�}`XF�(oH�X0J��od���Z�~��>��3�5��:k��>�J������G��гL��7/�Pv�&NL���V�)q��qL{�.7. ��z�O�����G �pj�:�����?�#O.g��|���%�n���*�%w��bBx}��2�s(��U�����uw3tX�N���&t���ՍA�d�|J[JmI��=�HG[�I�}fŶ��OSMYmn�������A�O�.��j�R��{���Ic�l�˿"CE �A�F�9����6`�:%9���Ǯaؔ�%ޖ�}�0/�v{�^<ؖs?Eӽ5�%ˀR�9}qIy�k"Է:"=)�:\[m:�q���![4�EM��� Y}ˎ� � �K6�+Ywbl7Z�v-�t� ��&�3xɬ=��$�i��Z���LU���>��᎘���?��4��~�{̗��
��%�4��]]�_Uvd����б���uH�+�K�ç���o�x��#�E�̹у������>�I;���)QU+�ff��ji[?X0�&]�.��-�98��D��Ȝ�<��h�n�K��]���ƻ�k��)KPˊ��+��5h��xfV��rf�R��������w?N�b�j?�nV��	����)�/����J�AOh�a�I҆���1h��䧐e�h����6�3��ذ��X-�k���eMw"�_ܔ{e�<�⺁u)u�K6��}
	�x'P<	����2Rxѡ�M�����he�$^99н��㔀��O�l^cMD����.��`d{��)��D�N\�a�6��H@�#�� v4�)�{��7{C�-��Jr�9r��iv=4_hVa�Fr���9D��V/v-Ni
1: i~��f1�t�꘠B��6�e2�����ș�,��%�k�ڱ�
��Z�P��L��C�qDi붴���?ɟ9i��Cu�N�f]��f�g�F�5t�>�V��?�$k������R*��]�Q1�yyi�x��ǲ�C@߳�����D��t�����\�ӏH�$Ĥ��T)���YlP�y@Y���VG,����0�#�ѝ�v7�@u����02�o?�[�
 Vmq�(��n�}�s����-v7�b�o���S����l8Q�P�gs�L> ���~38��4� �j&s�=�MZ�:���mɚ���� P�l��x�l;���ﾙYr�T*�Д��{���K��l�=����z�i�&�:��V��{�6ĥ�+e�H�w�3��2�0%��� ��LZ��$�Ql�B�Z��͂�ٞ�C�t�&\��l8?^��Fq���	�{�g�ёXp�S{��9�mY.N�㿚L�s���tf��^�<n��#��`���_�?8�r8��%���πB5�#�>ӍK4+�u۠��.@.+��ޅxd�i�CXYZ����f�\^΋mLt�̪|�e��;<0�.E�H�˷����Ǜ�<�+)5�v9���N��D���u�lOoI
�s�a@�@W!l g&�q���g[�t2�K�3�A�	���v��6dz$l�x����
��I������R��0�^��('�6;ܠ�L�
��Td|"����l�f��UN\�P��>����Y�а#:��q�wQf�	F���dи�>��x�c5G(�U����T}�P��J1�>��#p�<&�D"J�� ��(W%_�Z�Jt�
�!T�l�!	p� ���X������γڬЂxh+~�T�>�6'nV�t�̏�/�z5a����rv|x:-����q<�r��fa2B����o�m�6]����y�|!�{�gP�H��=쪺A=D�	�.Zz�Y���ٱ./�3F���~�����&�ZW�N[ݰ�V�P�_��|���#��
@r@NAz7�1���"��l0V,����S�AE��P`�1��@=�G�ׂYv���_�,5o�_��͈������]˹A���c3٩��H�����B�X��^S��Pi��kP�&�B�Ƃ��a.��o	�%47�Z�5O�R�������<^�i��u|@���|��.No^UE��FXC��v4��҆.�>����,��kǾI�Hьp�܉/�%@%m��.��A�VF�rSY����'�6ȡ�h��1V�:kE��o����J&���R��ҕf�_����
7�܌�;	���g����w*7�a���ÚL�dAAP�4F�&
�01)����_3@�k��B��AO��(��-��Bh[��U^3�{����5�p}2@0q�����K����9�I�Ԋ8Xx�j@�s\�5"���Ƙlg��z����.���wףC��b�s�l�~lx�BjR 1��nx��b�?ۿ1��#Xkq�7�9�V����l ���WאšЎ�h�h�	�������\��t2��2�ط˖����y>D~~T��j�oG��q����mo&�K:ž��	q�N\���J&ô�1�%º����h�d�Jz-~uy3/�N(�0�����%�nvƥ�9	�e?�
:P�d�<��*`-�q��$���g�;ܷ{�E�������7�U�)Ԑ��#�I���?_p��,@mF�CA�|�͸���a����@��^o���J��k�^c�;��c/kO)/�h�"%
n�=7�_YNu��� �p��H�'��Q�<%s�XC�f �/s/Ï5������/m���������7l����4����%
��-x7����t�LpH����-5�_�<�%���rr��G�PA'�"�Ƹ�f;N<)4�P�`�(�Hr�l,�Mu 8))*|3͋����֛t �3�_Fc�BoR;��☠���'H�+
.p�� �p�\t{mL���G[��A����*��za�BI��t!n�<yn	t���+�s͑���ֿ��Nu�3!�W����vUZ�Szg�,����A����_kF?�Hv@y��o����׍`G�a�բ��%{�֜�G�vX8
9�j�jl��Ʈv��.N�ے��6aT�*R����Ʌ�*��n��'B%�s'�=�����9���������c7����F�F�Q)h?xTR���J�J��5=�����~"�Ϙ�P" #�&�Ec��'��gV�",LJ`��D$b�����-I2-�xT��\����'����1��a��P(�׬��R�{\��Ɵ];)��?���a]dZ��7�,�3�2.�PR�|9(kk�49�9���� ���#�{Й!s������Cs���G�E�j^��]�-�����%�#^�?L�pg���D�����p�ٲ�+�YTY�>�+Hc�'�q�/��I�d��{���3f��`q�Cxe�9��[�йN/�$'-2���S ��%���+�_Z������K[:Uu'��7�moo^����C���Y�q�O�ؗ��A1�HwR�U�l�r��Å�g�9(`���d�qž*a�:�S�±�=C� �͝2@7��Yh4��UA��͏Q)(nȸϹ곒�$]F$d0�A��b�1�*�q{�yQ��"K��������yu�ޱm�j��F��Fc۶ͶI㤱��hl�F��;�{�o�d&�4��{��Z{_'4J��T[:p-�:E����9!4o*,@�лK����6l���� ��2G��뎲V&���}R
��������T�,�8������"��T}��8��?r�w�<���� ��Nq��DwN>����o�
��l�Fd�P<o�w��s[�fu�5�Z��Xa��Y��b��:�0�݋�D{-�W�ԃy��� �����q1I��gh\��6��LxV���
D�L~X��7�c�ĸ�S|��&	Q�K�9��
rh�ٔE�O�5��(I9��`x��4l�k- ��g�"iʿ����W%t���媛��Wk�Y��.�t�l}�r�MQ2�b��[��b�4

?�0w�)h`1� NL5:PR����u���]��X�ȇSs�[�s�POR�b`ݚ[S�*�sKI���I�}c�pr�$�ExnO $����_�NflZ�q��@��	:\������5�Tg9��r��!1�h�0�d��)�ѷc}O��!�+�i!!PP���ӟd!�Vj-M��c6�Q �n�k���x�zN�w]���t@���ǆ�|�^haΆJ�.9�<"�\���Y�r���x(�9�#��bR`2=R�"v(ȳ��p.��@|b�9��=�^�b�0C��D�ޔ(����n���kW��^�<�%6�l\��ٟ��
(�������0�<���m�ߡ�����r�l��yj���~�H� M�lE?������_l����g���+^�����z��t��Y#T%�����e�$�.aa��>�!���3��˵��tO�a�<|��@���dJ]�Q-t���D�q�7�8�0%�Oko�̤֙�p�+�����pZ�	�3���m��z�U�ëli�\ �1 �x1�[;C/�9b���)�@��Pntjr�U��;"߯c�8j����<���r���6_%���|p����~4G�6"G������G-�3��wW�%����<&���n?���,��,"vLT��f�w���6�dK|5e�E>q�V��Ȧy��h/|����'����t(�+�>
�p"bg�����˭�t^J0ebWa��DT0�2ᑿ�G��Le(oY77�F�@�����2F�vFM�j�g�Y:��{��{�l���'&�!K:����s7�mC80�N�8�#����e�&�[���³��]y�������\0��e����K_��p��=���u/����"{��ĭ���W�Ծ��`pXJ�%���#z��OnB(+�~-��i&�Y�-�~�.��
��2��y(8�>?�Wj��v�D!�,5E4���6K}�-�Ӆ6�a	Ye��jڮ˲m|�B�6I��?N..��$�TB�hҾ^/�-��w���m9s�^:P??_��ȯ����@�mla�A�p�`��֎@Hj�v�ը����L�CR5u{���k���3�� ��m����2K���C��c�h�#$$�����&�2���q���h	O)��!�o��ĝ�^Ӭ�R�Ʀ$���������2��f퐗�M?u��^��'d�g9�v��Y��T���7�s�\2V�b+�5�V5Ȼ��f�(&g�^R�~n�74LC9=Ԋz�t��� �úa�!��)�-@����D���\nT�ި��9�EG���{v;�d������яq�p%�dL�՝���-�$�*�����'���lI
�"4��b�G}�ӢVs�,9����%t���J�d���Z�P��Ű�s��=P)4aŠ�c�M�rV
���=(o�����ȧ�gMث���tP�H\��7':Trs�\)1b<_������8�X擂��?���I�a�ҭ��[��-ݞ��SI���y���׌˝�F��aN:3'�L1��l����5b���¦V��;�eҏ�wy�o�_�S�=Yw��Z�徛>ܮk5+�_Ƹ.�_ំ!�2��}DRQ 		����byo�feo��6��4'�	����)�U����fm>�����r�zm����S�#�U�i�C�������\��QY�����r�qޢ�B�.�w��h�7Q� LmI��+On2NQC�[h�){撠#�Ac��v�T�;���u.-`e37����~ ���\A�>��l�=B�3�;4�Xv<�� �/AA��WN6���_%�Im��ȃ>7DJ��k�fj/ۂ�z����u�úK�p��oi�����k#|ri��>���/55�E��uiڿ����6��G �֔oy?�%;j���cu^�y�p��`�4d;z�	eY�%�s����_I�<5ܠ��=�m�QC��o[�O����w��%�T��s���gτ�t+M8����ۂ��ꃜ�!���-�1��ۃ�1��}����g*tL�G����ῆ��j�&q8Y��[z9����r[�afB0��`�>ۖ9���jZ�
.�)��	�|h[Anl5!}�Byᔐ12Q��Z�'�滇 �,����a[o�Og���;P��<���0
0����p����		\��Ɏ��Lz��uR��Sã��w�����L쏪��׉�?�݊}ǘ�������1��K�Z��b@�����E��BKO�芥S~�>���OMC��t���",�#�y�V"�d|30rZ�=~7��3jWf�c�s�y�,�їK[~,ݓ�!n��܂�1O���!nn��r̪�<Y�!7�3$�'է�g�,�:8n��]]E�s�v�+[�w/Sf��T���	M�o�~bB+Lv
��c���l�=����Vj�P8!a%��Est>_�^�/y�%$-���5M����_=����86fаE�H�Qgu���C��*$��,��w��18U�C[�V��ƺm��x�J�I��č�S��e�M-(����v��ܲ̑���	q;z?nz^^;�Ż�Ƅ����s��"���n��$���/���	ٔ��q�=�,,b�_)M�}��ܖK�f�)�4�B�}���0^�ԅ���f �m��2d���,G�g�q�������˗�M[��RA�Uɭr�5{D�OoK�����ѳX�T�S1BY�ۦ�G���:}T�%Co&M��,d���lǉ%d�g]���+�0��z�=&��)�H��������a�P�ج�Ӻ��� 3���@zW�>z����&k��s�;#��>iEY�BY��Ġt����dy��F	+!�?��vJM���QW�LzE3:-��1 ��P1I(ȸE���1i�,V�3�&QSS_=<h�)@��Hx�5�g������i�sh�� �^�&lָt+ո��I(��@nۍp�^Bg�c��VD]K�Ж����W��DSd:J�{�p]�Y�k��)�6�6���g���ȩ!b�qÀ��7� �0;J#�Ǩ;�04��v?[I>Ƒ~��3�LD�%���]c3nwm�gzI��;OF+T��~�@���pN�`!�+�'����D6U���!����'�Z���Gnp�,cƢ��0�̎-�
��ߎ?�,�,�2.�&[�R�\�HTqBd���EU��7��()!Sw�:M�����4���:�b�+d8�l \���m�cm�Q��Y v �3�/������WN<�uz��T1���+�h�� �KP�0mȩ��c�8)�TL���%�R2��������&�yh��Kw���>	C����.��Z��hkQ�!�-" ���N�M��.����Ն_7��և�����(Svʸ���4���5Q��Z�!��c<�PZ�a�Ko6Ѯ:
<s?�I����j���f_��z>b	&3P�R����禜7�����v�#�-6}�9�`���?ڟCl.YcQ���"'�K;M��gd��Kkݍ	�%԰��s��Mҝ��&�]�9�3�&� ��}YF�*z�f����>�z��(�*S=�`�<��9oB�� ��^�-����߫�bEK{��key9z����ǔ��WCe�����+�?
�e{Gpm��

�������us��>x�z�����)=�?�=��{���?R�ȓ#����d������p����n����f�&�bV?���5�#��-���r�(�6�Ұ/rH��� PK�L��h�iL$��Z��6���`�ku�}��fT'��M���ֿ���+[�F���K��c�XJg5q�u"7�Ac��L.}�Ѧ�f���I���0�%�<l�t�p9��\&n�_�/^x�]� ��R4�i"6ʄ������J�t�H�^Lҏ�T�w�t�CrJj���8\	�L~�+-�G���N��Vh�~��[@��{UuQ� 䃑�X�z���5�ºn��t�:����r�	 ?A>봍�͋�!�-DP[���[�P������ʕVY�c�im��e�"7���r�������>.��X&;���n����Nm����7�?}V��u̓J��k�.=��*@z�U��M�����1�*��/`Y� ��&}��>w��$�ddz߄�a�[8���R�Z*�{'zN�psh5G~@���
3CLWO�֫c�\~'%��2� ��ܓ
����x>���ח��+����Y�� =\�� �wϋs��%�9.N�ȱ�O�/ۃ/�����P�RRq ��S��aV�P%�o��3;YD��oU��rP"׫�������D�D��s���t�ח��}<��<��		���"t	@B��
�#\BgS'��ӿ�,[�"���h��gi/�o+O��V� ���� ���Z��t�DWx[{�[Z#��o+C����4k��T�g'�W@�u���1�y&��v#D�H�2��7��:y�c�`������~�J��±/����� ��|ѳy%iM�~߽�d7� 6D��0p�E�Ǒm; �t����(_5,�g�[0�/��qiM�sy]��;̈mͪ��wGd02,��uY�l�{����	哐D�ᾓ���{ߌ�s���G1�+�!We�j'
zM�`�=��� ���&��yW�$4��)�$=�n�¦���`��߱��*�+� ˘C-(.b�qMu�6�Am���"�}�%o6� K:�v�2�9�� �����ܚH0x��~�����Ӷ	�K+�-D�aCT�ݗ!�<������ԉ[�[v'�L�b�L����m���5���PR �dM�k�olWkp�� q�)�q��Q��XT9����ݴ�YE[��Gg� P|F���G�3�U�b�h����v�}C��R�/�K�۸�����Z,�\ڬ�Y}�5|4��Y�	�����5*V.�'�;o�[�Wt��@����[��� &~L���z�.�K�������	BB��]}�ᖋVp���Y�kk�^���E�+S��&$
ب�����"��/��6������F:�8kYw���ޛ��я�����D��$H��=����Cvk�B�)�;��;5��֋�́�䕮oxAX!�X���Xr{qk���?�&"��O���sF��NI3�Q���~��K��UӀ6`6 @w�t4��z�;i�{�x0]��~����	֢\���{̯�?BQ*��cs��Z4D�&y��Q������i�9���t?�N����L�1=��<��+N���=�/�����m�m�/��CI��kA	PO�M���n(�e�#b��x�	�,��;��	��� :
�81�t�s E��V�&���'��@�*\&f �S��$(D�e���"�g R��T�t��kЂ��������qU�y��i���_�QGԢ�.�Ǡcv:���q��RVݚє�L(�Ť�����k�i�$~�P&��N�_�Y�F�5;�D��� �Ě���JHgF+jw\�Vp�nmc�XXX��Į�K�{�.<���3ܫ����nQ@��`��<�v��:_��9[�2�<+���~��\F.�{(�_��ʂ�[92QE�`�`�$���W* �(�r�z]�a�Y�]��������u���F���l�V��W�r̜��p��Ciz��)�t�yw�:7^�^FE�[(�	�V�7��|�Y�ur�(�%`BA��#J�����K���L��S�Ө;[���֜?�s�4$�Y�R�L�|����l�d�$�L��D�\��5ϹA��a9f:Ix��+H�]�Q�y'�[H��d�k�+��J���ŷ~�D_���Ue�B�J��J%�Q��S�!�X��� ��u|#䷸-��26�Ԁ���H��!�0;a.XTҩ���$}"M�V�wjuJmp��kh�GF�Am���D%D�Yb��`f�M��9_������k<��Oo=�Zח�RE����W�}�`��4[�K�ٔ��6F1�zf�1d%X7m���̾�ޅl~n�S.�A�e�����7Wʬ��2�C�PD����O��a<��H���nSbS�+�j/LA"�AKG.��^Y�Y�b*O���R�� O��cG�ph|�K���K���c�k��ܩ��\�[��ǇR�������T���� zwY�7�t��kM�IA�I�������gƓ⮼絫g�	F��k�k~&�^̟p� �+���cj�5.]=��W���]p��d3�<�|�V�L4�O��h�2+��r�?�����4z:�������m{�M����k����7PmY9�
�
�=��m��Ћb�<�%�ӹ�W�4I�J�"�4�X�ai?M����ގ��l�F2l�Gp!t!�\݅~��4�U"���4����\$���x��}�6�䛎Ç%A�f�����|+Ŀ�����5��\#����ߩ<��"m��<��A�htRTƋ�<xt"�y�t^9��ڬ�U���5���A9�ݧ��/���� hu=<#�2WԐ�<t|*���ύ��u`�h��ѷx�����	��L"$[^�����0��?��L��j[k#�#E$̡(�)�r��=�.�y�Rz$�Jr@y+�I��Y.� A3���v8�� J��[���z����wTff]<RR����?և/��?�Vi�+���Z�(cG����oN<�5��}#�'}E�Í"%�l$k\�.�-�bI�W�K=ɠ��av��m�o<p��A;ޥP��8+I��:�9�V}E�Ds�EC�m����:�lmΐ��9U��޽_q�x��j8_u���Br/��4Q�f�m��;"�z��͜1A �5�Cc�.� �
G/�պC�[h)2�JMD-z�� ��⋸(!�S��7y"�.�gh��j��#0We#ۿfC�Hw�\\�#;�VV�a_P��%����﷕�v�L���iwL]L�4�"�~������Q>�����A l6�8:@�?�ȸ?I9ߊ����61Y�xl �@��$����Q� �#�@�����������z�'����I�ǫX��L�;Ǔ��/R&Z�53�L%T���=���J������b�7DA���t�E��n�:RP���uq51=%m'}a�߼�w��'f����$d�]��ސ���2���Qƿ�Ŏ�{ܤ�����--E�M�q�n̦��������l����w�I���°-�)Q"?-f4�b{���rO�� ��5��G��|�������c�̏���J|�'�4�ߕOo�x �܈*��K�lb��A��s���r�ZwPt����g�	wL�d�f���"�8b�H����������f����ٿq��$6$�T�n�W#�����f殴�.�#�`"�����1`"TS� �Q�@��Z�<W[��?�� ���>�>��܋����&��4Ԟ�F���~
>am�S@uWV��Ř�nk�@n��Ҳ�˸�>�7��߹�S������~���Ε�
���>��Ս3L��+T���f�c�~oTE=:��S�PgH"*����Pb	�6v�Գ}M�3Yg�~;��@y�E1*q��ix�T �;��
T8�JW���I�Mm��FA=D�-k'�x
�s.r�e�u�ź�X�h����AqsV��s5Ӻ����ϸ�^�$];�ż1{f͖N7��M�M5��qA��B~�l5A��n^�����P ~u����>��KH��m�����6��ɩ����v�N"�?���U[;���#cB%Y��Q<H~1���'�>����B ����n�m� V���>�:ݧ��/�+D������M(���� fy��NRЛ���v!7���ˬS��'��Tp�ȃ�G� v"���\~h��-��K�����i��gIz�vv�b�[����i��:�m-Wz[&;��M��P�;.��@,���(�.$)y2�@�^iYm��h�B;(�&�ƻ����������ྌg��Y���ar[������,Vhv[l#���O�ol� ���>�s���uῲow|�0Y6����޹؇t4�f���]� ��r���@.C..��ϟ���u4�:����J��R5�#*��.C�ױ[Cн�>�i���:A�:������-��|�mD��QS�Y�h�"l��m�_���Y�y��w���^[Y'p��[�� 9� ���u���*�R*֖0`�9����ջ������V��k���n���E��l|�D�͉Y;�zي /��cehc=���!�⁗�X�U���G�6�/�/�-���^�c�,�{�I߰���J�� �Ƴ$����u}k'n�w��z��Ԁl����̣��E�*Egv�_[��HI�d���1�ނe�ܛǆ��[�p�/��ߕGu�ު�J��'���ڎ�Ss�ϐ�Gq�|x�o߾ f3�픋&^@���͸�2泯T@�}A�f��ujFl�?>N�!4��9|"-~}�^�m���Yu��콪��@�p�c-BKUS�ZH��،�N*E
{�v +���^Ж=��)c��1��g�ml����!>��2���I.�9�����I�yT��3�(�d-�+�Bvr
p4�9y��T�$�D�m�)/D���/�&HqD�G�������e���]�X>aM=p�5 a\��?���N;��p�n��r�tgda	���rA����2��^��=���Vѝ�"�uߋHHj[��ܦN^Ɋ�7�2Tx�R��=q3�P���)߁An�׼�xՕAX¼�C��ݥ�����|&"D����ŕ���H]x<� ʴ<�Wی�6���س��xm����)n�}��3��
7a�����c�l�h�kT@%$4�6d�R�-��&��io+�ŵ�s5�̳������_}��H[�nܫ����Ju�/�k��$��]�B��]�TES�u�p}����^D	4Og�P <rR��r�� ��xj	I��
��I^��������ڢ|U�w��t3�=��cK=<p�Z4���yh\q�~���'�r�ʹ��@{OM��_n-:��rF9J�DA/ı�]�*z�|\= E$mKw�A�Z0�0X�q�3�
,���4���~�����������4�Ǔ_+�_i5�5��¶�"�׻>���ntC��0�)ʉ���v�c���*Y��Wʗ�� K�.��������[J�I�D�Wn���|��j��6��ʵH�w�&�krȏ�o���׾��4�U`��r�g�u�Ǽ��af�!��U�/��m�_hޫ��Z�
ݝ�#�y:Gџe.Vf�P4����
0"J�_�r#�+��|���0'q�ꮭi�M�r������U�	34~@L/�-���Ś�|`Fr&r<ZM�ۨ��з @1�%l�����P�������k���#3�>�(��R�� Y�phx��Ҙ�{e?b���蔤���"�Ta�D��O����n�Uel���i�C0������qs����=�^�D������Ҁ�e.1@xI� ��Kc�ح�:����?D��hS�;�#�6��urfU��km��=�Ҳ�D�PLΐ����Wl�!�%~K{�7���v�ah��TAPe�e��8�E��ԫ����S�H��P���-�ܐ1��1I5i�^k�~ڄ+[+�6��L���$:%U����=�MlE���x(
����Hj4ho���O�%��]C�	д�U�N�bIp�ǔ�v�-F����s��ﴚ��qk|;��t�?�+|,bJ?m�Gww9��>��Ϫ����4�8��y}��2u�9�}m>�r$�6�}�T�\!h=��G��xzm踺.L�h��:�n� ^�$ ՏPTL�@>^��9վv.hT^;����f�fx>^PZz����u]nk���u�)Kq��*k�f�lJ���!:��\�<\Kv5k���v����Sf�����r=;��FS
e�E_�
�G_@��}�T}  �ƕRT����˵>�#�����xkܥX��>cS_J*����b����ߧ��-���U����f�
�X��o�����[�.Κ$Z��9��-�ac�M�9Y��1Ȧ���,�zn����_`!��))9�s�P?�_�97��"�QD�i��w�/"<���$����¬����}>u�Yڅ"�~2��8o�­�Ð�v@/r�R���f���MR`�=up��k \��B��T$ qԬ��$�F(W���"	=qy��p,�
|��j*u��\��S��-W���zk���ϤT4=�sK��E���`��]D���iX���0�Q�� �S"���`�*)3#2rn-��`ok�g�܊��x��Y�a}NA���2 w�ʿ����fʁ<�T�Q�`Ӣ��h9�d�`�}xN;v��۶�s���T9���B�6#LF���q��Ϩ]c���e:�?���w�;��K�+�G�����#���x�������í�E��0�s�%{���@�!_|Ȓ�G�Ksx��O�/��m@-�8��$DU��c�G|���b��p��>Ia�������jܝj��|���F�^&Y�;Ӫw��蜄FX|�E�#;�ܡ�ƫ�@41�W�ɔl*�MI����� [z1���^{aZ���֗Tw��ؿ�Of���:㻗�G����/`�X=-hB�h��[�m�(skz���f ��E�'�����dxH���,J��
v:�r��tGh94BA����^Y��C�&p���)��a���-�Zr�sDgm����-�ð�Ӆn�7��E�1�l�φ;h�0˶�a�:~?>�I��,M����(�W�]XV|�q;����^�g& MUh7|�F���@����.�&��5���K�� �I�k�Q������������K�8f�U�#�I8�&��Q�r*jð���i�/�&�����|i�SKzv�қDiV��""�i��FGn���~���Ќ1��Dƀ*s�ȶI��2�&�&t�-��󫶭�ԑ�8Պwh&�<.txN1�[�	4�FM��Q*���Fz��3�������Oz�:3Ĵg���Тrt��G��n�^X�p��k�,���J��߼�� nりD���?^x��gQ��.�UԜ��J)�DA��Q�k�|���;a,�;q���æ�1��hgD5�3��J��&W�=��~�P�trTlп�BA�<W);�����.�)iu6����j�����\0�Gd�����@�ɷnx"R�*�1Q����%��oe�H�������[F�?*��/��qm���f���v7��#}�R���>�pd��Ru�
�|����[���Gd����`W�����3w�`C�`�x�YO�k?��3<h$],�JIs�`���Y���5�[Pހ�S��7�?��v

r@�n��*yDZ3�A�v�Yy"��ԃ�Шd=��+�-�%ȅ����pll��uUh4���ҳ'z�|���/�l,�i!��nzCgl�
�=ؖ���UN��_.�w`�V<�o�D��P,����:�RE�?>y��q6u�x��+{	.,i<g�OJY�����y��O���7SB��(�ܤ�H��E�J
���V�Vr��B�l�F��k��'�j���2�۬|Z�v\�����
L軃/�x��x������eՠ�ډ8���\G�qhи���t�T�5Vh�w�=�G���`!!�q/��V��7O�1�i�����u)�o/&�i�-�`���<� EUT��x���eS3>h��ql'ktɶ�pi�X!lЩ�D��	�՛Z�Yk����EP��N�:4���o=�>NtTj�HL�}c��B��Y�5NLW8�#N�LÀ��v�YJ�P�5X��4H�z-��m>��Lթ��xx/�sG4�kjr�B�f��$J���2?{���2�a<GRQ<=�����޿%*��5�����/[�sh�2�x,-ܖ������.m��̜��+Ɋ���<!GQpt�12�c��F.� ���&#�������|�OE#��a�	Q'�����o�r^�Ӌʾ�!]��{�Gś��������<�V��Lo+Pvu��9X&Z��y�S��C�I���s�+vF�ǯ�&����'� ��sY�Y�*������W���.�_(ؠ)�Ř7�� ��{��ߡ�$��8�����[w#��^��p�����o5�0-
��',?H�3����1�%�81Ȑ��r��q徴��wȞ����1����.�|���W��R1���e���y9{�%tǩ��Z��@�!ay�����o����\�[��"-S$��ι�����Gk�*k�X1@A�*��Q�QF��@5�,�(�I�����~lf&�_�f.��?�j�E��ӟ�����ƙF%eQff���"�r:�K�Mr:j8�07�Ed�v
ct 
���QM��x�n�����S�}]������H�K��~�������[Ƭ���\$>A���o�Mvi��n�NV�Ԯ�sy�]��p�����э����br�0�Y��2:p0?D�%�OMg�nt�n�gP!�`�"�;�4Q%�$^ܖVm��a�;5�Ers12�Ȃ�0*���ZvN�һT��<�̀��qq��6�r��7�:a��Vt HH�6Q��o<~���Y[��i��N��[�MH��	N�T���=�\��E��K��^���n��R��eb�l�+Blb)s��ZN`�@���`X�X�V���ڎ�7�X�Τ�B�/�K���r�8
&�6~�9ptq�B*"�l5�p6[��z�x��7�~��E��J�=0HV��KI���>Aj��A&�錙�UMMv������9[S!�e�~���qP��z�כ���"6J��p�\�~�_��ck/n��`����*�����c��`#�+��C}��3�uдUd�hn	��2 ~�~��Re�5�+��B䡣c&㔴����Ћ̪�.w/Ր&�0:���:jFCbu4ك�s=���f�����COS�㛥g.6�*0f��&�c�3�7�K>�P%#� ��#��OE�%?��w'R|\�m��F�:��F����8<;�O5+^=�}7_v���y1�a�!4z�J����+L�.����2��cRð�D�0�{�F{�O�
 X�����V_L�ǯ���kkZ����a�i�DG0�ax&���?�D��dk�]޲�b�Ư
[_��{�x�8U=��.��0 �d/I@�� ?�]��Fu�6q���&9����i=��/8(=(:�0��DZG��-���I��+ۈ�x��`;O�\���s��"XF��%��-���~������v*GD��n�t<�r�j/��Z�6Ni	Qc��{T4]�o��U�Ok��$��m��*��[>n��2�܊�.�.6� �u��rm����r�59͡��i�p�!����+���R/2��o姏Be�URB~ջ5��ǝ0+Lv����2#J=����#E;Q��g������P� Q���_t@��c�����K� ��3ϛuL<+͍�1�Mƶ�n ���EZ�C��'��LI¾�A����w�-� �AF�*|z6��Km���Ϟ�������!�(��O#v�$�U�*�B��rK|��]�i��L�^&��]��i��Tf݃�O�gu[���?ht3�T��M��k�fnm��w&UBˎ�����R�ʸ.B��Hll-h����_E��P��s'z�>U����I�E����pb�,h�w��� �H��`��s �����r�4ܑ�a�E�~�سI���d����� }�FǄ�i#�+�_�E���j9E6ٖ٨��AIa�]Kg+i�ޯ�l�z? j%�2}J��)if��́.�C.�^����3�z��J@���.hm������@..�A�Y����`�(����Ä�z甖W���/ n�k\� ��8,�u��ڤ��"T"y5533a��:j��͑�y�\��.�|���i��l��M�I�� �#Q��#�Y1�S}/�]X�D.I�A'��&�c}V3y�]�S��F�x����H5��2Peb.��(m՛YL�Ma{=s���(�Тk(�8
�?@�����&-���S��a��T�}?u�.�X����Ɋ�C
�/[�ۊVz �Q%��<�f���J���zk�*�f �f؎{W���c"so�+���m�9��R��PI�m��}����Z���6�U�k���.����ko��:<���ZESR��ukd!����ͷ`�F�#���n�0K�C] ��6���6���]�}���;�*�&��D/�Ә�5
��l$X�@xH}�8�G�DlYF��O-�y�"�;�F��]�����jU�����
��_U5�ov�֚�Nl���V�JϏ����(�*��Kt�i�/�p������Uϓ��X�b�p�X����b���P�@ő�G�ݎ*@����{-	��~��PIh����L��0�ů�0:���K�}A����|@�F9q�|}�1� :��y�ǝgڗ`lr��|��җ����[�ܔ\yx���)<�D���I��Q��� �}*�y��E�̞��(����%����3/FH� �jpB��}s��N���؟ީ���W/K����gcS$���J�)����4=��! F��p�v��o�h����p��x/�<9w��-_ �?��z��b;#{���>�"�2�_��1dɢA��X��k��0Ѐ��w���ߺl8�$���}?w��� 
��O/�0f�ַ�v�7�-�XA%����D*(���Mغ0��Ѣ��&A���%N�g!I'�`�6NF��|m��m�q���n��6�Nc\-��w��ڔ9?�g���s<2�
!ԋ�Mxpb�����u�I�b#�S������ąHbR����`�1p�R�c���r`~>�L�{��`9�쿳����;$	���`r�*�3�s�2xৢ-��ȉx)G�W�W������qt(�G�=,K.b�b��Lg7I$��g�5s7����t�(j+..:����RW��G�z0hʶ�����{�9^��y��o��V�	-Ԫ��X�5�ׇ�\�̪D�:-�Q�&|��D,D����Z�s�>ؖ �m������"	���+�^:�D��	B��+�:���l�{\	3L�2���՘PI��99�:�P�p�NN.RF�fM֜P|�IB����[�ډ��<H́�T�։�?����ַ3(�L��4��^�E��bK�U���,�$�P��lc^� �<EHխ�V�z�g�X��j��u}TU��߶��h�*i�!�q%J�#8kdQ'?���2}~'W�S��z|�kkB�2�O`��mG�+��>�1�؃�8��+��c�s羢�k����s�@��y�e��� 7C�d̾&˶��*�R�i�AE>cS0�����EGn������_k�p�8�w�Sӝ��!������*�LCf[�)n0�����<&ך�@w⚪!�pBA �?!6���j�7	-G�1�������U������y)@*�K�--�&A|��~��������t��K6�]է�c�OKU��j {�yv���
�t:�vC�4|�����~s�C�G��6�#.�z���[6�q�!�c� p�J�/�3��Q��L��Z+N�,�C���Ċ��U�է��`ZP��3^�QB��P�MW�<W<U	��N�|\� �DF�С܀`�\qf D�G�mRs�"��wY�MX�9�K�T�K�"0�Aԗ.�kTl!u��Y������P�:�^8A8���edl)j��hΦ ����H�Ħ��
p�bWо��&X�1*TLb�V��V��0:zF�2T��P��Rɾ}H^H#.�i�q@[�a�f��g�&Ʌ.9��;�Fy����>b�C���A���2�Ml�X�ךXW�\Y�`�cR�:���>Ẕ��=m���AP�H��Yp�U���|mG��>P����uՔۛ��ra�pLr�Te��ʺ�-�J�gҕ�;��e-�|�9�q�LX&��=}b���F��m���<�w(��M$�c�>Q���8�M&H�;q�@y�Wi�|U��A�_�}-��\�q[ALP�r4@��c�p�7�觿C}��#����G(� >�6$E���׷��J������u�AuPa�;�9��a�E����x͸P�~�P�
��E�J��ͨ�0p�f�OD�4�5�A�����8B_zԡK�_�s�︄��O8i�%��/�NO�fE�?rc�'�f�7�Z�!wI�`��$�^\��--��w	�{�p��j�(s�������L�� �V�3W	M4����zӘ74-n/�bu�	V:'1nǑ1�p�n��G�$����`����lY��!�|��-;#FRV�4qmk.ƙS�}J�f5��޼��{8)lKv�aiO��I�!��8]�^��;�gj��+7n5-�-I�"
[�ҷ#G�����%B��7f*���Q @LMT�/�Ba|������/hХ�pdR���"T�t���hb��h)@?as�Ҥ��R�����SV]��BC��%��;u��������ֿ�QA@P@@Z�C���n����VZ�;�D���:����=�������{��{�k]߽��{'��z����^���tO�y���4	�к���`]���$���uI����;��:l%<�KKdK�B+�u���;�¹�u7hN�{ߡIc���U���Y�ل��&�j@>`<�hy�W��{�\4V~w��T�^0�����ߨI� ɥk��=�܋�"I��[#'��J��!/?B��`t����S�����)��D�dU	m#Fz�;}Y#F�FM�ޭ�U�dqa:��7�=;� �ӈԴ:�Ŏ?܃Q�^@��Y����ϋǢp-�]q�#���_h����M����<�;7_���޸R����⋒�2�� ��q���E0����#'k�soz��أ���ѷ��\���Z�f�b�b�K��*>�k�a��`���:��	v���C{� ����G�ʗ��	�-�|$$�=�}�F(/�.��;��&�M��Ww�F�)���^�ۥMء�iG? y�����N�;g�0���>k��9g��\����'f3��~d���vLN�g�e�T_
k,Ԏ���u݈��g�ָ��P��W���?��Kr����(p�}��1�~M������!D?^�<�%���9�7LΓ.��U�6���½^;�r��E�W+U����f��k�M5�8W��_�'~I�/
�����C�1�!�jOg�g�o�������CXdJe�}Kj���:�S�������r�G;P�H� $����)��g����˘������u%���$���O��<��X��i�����Tdg�wl��8��z��p�p�cl��#��c2BY�2�����9�?3M���� �:�^��x����e�#(3{��o��6($����6�mG�K.����,�R{>�-0��׮��6��)'�$#s���`p� -o�NhM���3�[w�&x�^c/1eA�,��2��p�v����R�sN���G��,�ww1'� �()�����x�nX�@�,o��-� NpT�C��u�W��n�.l��5Q�W7��*jD����j����6�l��$� ֲᇲu����h�[���e�ADdU��`��:0��Y����#�"b�&��=�xB`�@��S�U�d�+����ie5�0�kQ9�����nږ��R}@��z;CJ�v����r!\{X;Ɩ�-�3���gM��x�7?�;���fVR�j��-�e^�=�lU�Ӵ�P�ռ1�8Ӊ|V�[�����S!�St_=7%�쫖_(�Ã�;'P��dD6�h���I��4��������lq�r��_�j��k��N�ϛ޴�moezdX#�z����xw<�m�|�T�.ާVݝy��nc!� �jw�0G�f����~�B�5��ڌ�����U��`�V�?p�8$d���P{֓�1�xr�R�뫠3��)�m���B}�C�nr�S��<S(�i�3j�d�@B���h�h�f�k����`/�_���*����A�~�������勚�����ogH��m1sX�/�h�2	D+�,����=J�UCZa����<�Rg�"�#�eѸ�x�m5���Z���p2�\J��1�}O�r��
��&~	�_�ܸ	U���"<�&#L���х�T�a��
5쏍�ꅯ�]�-F^^Ϩ�C��0��f��`��k/ȡ�� #����`�E1S����S�O���k�&ZE������wO'l�ŭ��Ņ�a߈��t�U�17�$�A����e/QQ%kd����kD��,��ev^
kq)tRv(�bUe����#Wr������ F�K�r�t�ؾ���_-N��5�͹=������՜�q})�¹�x�${@\���XB,�qb��)-��BDo1�Su�b��Ϗ�ʚ�c��D���b��*�eF��w�xJXUP�jǇ^L���iRt�<�	��c��֫5*�q�7��H�dN�w�`2�^���-���4��������_���{�<������84�B:Qr6�y��'4Iw����,�QNϸ���~e��#�����uv�Y���M�����F��!~���j��NOS�I�3�S�|�A�e�k|=� 켫�����F��n͔y�x�]��L��|���`{��>I׸�`���Od/��&�H�>3�����ұ������5<�&�Ax����ka^��"�[�A����ꊦV'�u��~!y�L���s���65<~��Ꞇ���˥�aI����^�]0_�uQ{.�*=����i<��=���P�zX��u�u)Nc���d�$*TW0���B���@�J�D.AѸ���/G�Џ��ςYD�1�_��m���_� �|�C��i~��`8�e��̢=���
�Zβ�9{��;?Jv��kR�j�}W�ζή@t���t�����J����ל�h��3m3-�g8>��m{�_ӥ����^2��z���dȟ��ԕⷎLG���d|c���j���*��S��-�!d��2��p�j�.)¬j���D�*�NH��/L(Jb�9�_�}aʪ�lkKX{P�J���]�2P������s�����H�H�\��"���/�
�[ƪ�6�M~6�G��h���,�D[4S*Go,n��|�Zwr�^����vj��E��'�״�rz�=�?�m<�{�F�_J9J��M������y�W�Rҷ�R�S��ϱ1�LHL�ty��Mt�y�d��1ݕ�\�>٤dsW��WTn���o���Q�䢹G""�nfc���{�Q�rTa%f���m��@��37�� �5�Vi��AZ�X��,)�(������E`��+�U���e��#�&pe�IטK��7Ս���r ���Ξ�̛�<]��X��7�L��&-��O��K���32{���TgNF���y(d��)@�P\
M����9q����6w��В[]�
��0��ǌW�k��P�o�.d�Z=J~�l/f�?e��K�����(� ����(�
9�k@%��s��G�:gc�����*��O��}!1*[1<�'AM,0�9(����UWd�c�{��+���%�M�z(p��"Ρ?|�3�g�T�Lg\/LV���ѥU~�S4��u�1�#%Z���]i'�h1R#��UeژC���H'��{�JB*T��g��]Ǭ��7֫U�����e��L՗r"���Փ��8��;�W�ē$?�C�ؘ1�����LgJ��S]���'���q{m6�PW*�ۭ��,7���{4���^�f��!��?;�ϫ�PSQ榱h�x궖؇O�@��s����=ϋ�!�au��r���x��m�a�� 1����{31�O�,�_d���nxNW%�0FD�*�ut���dzؗ딧	8�d�%���1`_[(���t����z#R܇��T]���)���-_g5 �a͓��F�[���E�WY53���x�E�Iw!�4�*;cͯ��m+m�`3�j#��շ��ݝD��@ l$�����K�W����(��4���|��z�����s���K*xϑ��M�W�����t"��8k��M���eܓYn�x������k�M��je��?2��O��_� G�q�/�E���zw]��`W�PA7������p��a�,�i���y��
!gd��rբ~((X��щ8^�ɼ�e�J]G9�w��ʚ��:|��TǬ^>�|����꿿a-�d��!���U�{b�-|Ҳw�X��_A�͵[��Ⱥ�#�̰�K�ʜ�˫�I�*��h���s�c���o,���ݙ�@�Z��^�p���uF��K�;cjC5�B�֡w���$�b�u����B�������O7�R�8/U�]���4��x�J�����������io��?�[i4��ŵM�)@��N�)j)r��*l����fީ��%�0����cوD7d�j��=,�A`��e�z�]+N�O7���κ���2�Ԑ0�����Q,�����tߣ�b+�
���V9�x�_���	:q[����٪]Q�:꟮w5B�/��Q鹪���W�G�-Қʹ��蜢↧��-�a(~�D:wg������짧%�ѯ��3{�v�s��S�����]���'�
q�~{�{�g��.ɱH��RGm�y��К��f��F���|�]��K��|`������(|1?%ŏ�㇡Q��X%
c���!f3�Ő�a�?�8��5���X�/��R�6���?���H�羡�Kt|�Xp�������|Y��%/Eʌ= �+����c2j��L�6�n-_��W��.&�1�c���VSS�j�~� ^�jݽF&y��j���w�;{8ʞ��4�ͥ��>��+5x����ml+��O��4C��	��W�m�e���wL��.�.��O�N�8T9Ұ�j�iV%0Vq�F���o�$��5jL�����ȫԣ9}3��Y��ÉC<�^��#X�O�<�i����Ci�Cq}�x��E�K�y�1��l�l<2a.��:�O1�ۙj�dghkU�?G#�=�ܦ+Q�_�3�^~�>��.r+:�o�Y�V��'�g��ضcU�s떾���GPAh�ӆ���Q�2�e��'(?����|���|�2��I=q� ?����#>����M�d7��z�xϔ3�n��\��V�s<ް�{u��8��~��G@��zg���+0�/�_j�Ջ)XǬ�$5dp¾�{x�0����!!�&���Y���na>�<8`���nRΩa�_�aU�t��
��c�}��3vS��
�;c���Η�'VT��I9��-y@?(u��<b�a{ u q�u���r�����$|�O���ߟyT9[�=�kBr�J{�_ԃ�5�t��*{�$�}��h��.<uu��</"<��d��V=��:w#ϖ�I;�f�� ��q�
`���\�H_¨A�ўc�6�2�tq1J�8�:�T,ՈU�[sD�(���(-k(B�m�퓩�u��Rn��}�}T�v�tٍ�3�"|.Z��`�a��0/�K��W�.%˪ت�)�'��O2�|eg�_����8�3y]�Pڈ�[id��g����~#������.�`�iG&��A"���������ǘp�eP7����@6�����.w���z\N��o:����B���O9�s{u�n��:��)�v.�݊�;�lC��-���j����ȏ]��Us���G)�%��plks�??����t�������(�������0'���Il��Ǆ����Ƌ���6��$C��ݵ�KA���
���/���I�?�Z<ײ{�U�@����_�i����ՓwK��De{ʓ�zQ9�am�p�U����O~"��c$��2�١�$�|���kӞSG��#$�%ɷ�,_|���%��j;�bdk��R5$"���ǽH$T�Oy�|��O�_��ӻ��-=�'�3ެ�%��3�nL":� tn��8e�qӲ��Ԫ�m��S�s�p	0@j�{���W�Z��!ְ��Kh������\�$���R����l� �
!&kbL���t+2�{������7��x;�-���@�]��ؐ�h�m��A��#�&�}e��'c	mD�G�?�.�9���Vb&%#J� �J���ky��	P	h�4��(�?o�Q$���Z�S֚I��:d^,M%���=���N��Qu��V��".4��xGy��03�)��f*�JτƩ7�zc��zU��o1�G�K`��>�p���u$36���[4����q�nF�BY�vj2��2o�Y/�"/?<�U���Z��˟�|�W��+�>ɽ� =�[��L�D��|��
6﨨�����S��I)*O�y-���7 ��"��%�Y�؜h�ؖ���+_�Lr_x���rTL��	Za�S���D��.�MR�4��/�^с�}c)��rN����k.�Z���jae�UE����1�h)�
ϠQ
,>yw�9�R$�`�Yބ9���й��BV�TѤՌ��J�[�if��2�)#ό�)S���.Þ��K��	��;�U���hǜ�8�y��i?�����6�2iO�]�ΰYK���ʚ�i��XC�C���M�.�sj����HL?��I�y}��Y&�'�eI*(e�~6�N�j�%Lhy���2�QYŊ���$-" ���p��C*���'�Rk�g?�&r��<	�����t���K��^���V�����	��2��{S�]_ A'������@�NB�;�+���7?n���}���կ��Qӂq)���썓�ч�����l+C�I�{(��H�t�����F�	_���ʹu`D0����kH7f�T�Iz���rVMY[[m�%�3$��X%Z$�kO|(´�_SW�p^"u������󅶲��ļ��*��Wб`:�5-M:�R�Hg��,�u&�pU�PO DaB���Sq��9��6�;�^��p��ǀk5\�He39�_pN^�����0�礶�K����sU/#V�f�:��i޽0{�ΦbO�oe���L!���@@C���Z�M:�IVG�(}͖E���f��9@��؆�G�^��J�E8a�<`����o�o��Z��E�9Q�}����/�҅�S+�5-���WL'�2�R֋Z ml�5�TH��?4�����Ƌ�;�k�w4���t�������z,�����x���֠{ z�"�"��|8�H��m4G���\��B��t4�| ������)���F�W���O�IVa��w��>r��q9l�RL���sM����Mu���i���%��x�T$�`�ؽY���n�jU�A�_y�37�x�>���+>%��^a	�Ĉ��z���\\G0��7xLw���(���9Ţ�n�C^��[������/潅�A5	��_�.�.e(�}����E��pV,�q2R*Z�)��E��2����9����-y-E��& D`�u�;_t��CsC�ӷ�c;���Y�=^�K��1L1�O�=Q���m�E�p"�O����qh���fF}Mpv��]�^�Lg+��hP��=b�w��/���Փ_r9v������i�J أn44��� �u�u4,Ji���_�Z�,o��>�^!ib�X�+�:�Z��l�'}.tT	�m@g�nm��Z?�V2��m4�0�R�f��驾�L��# T��� ��������=��eu/'�d�"���R��i��#�jS�ؚ[�?���>�O������=RU=�L��
}�+����hH���)U�7p��F����ŒNI���4Z YwM�Y���KI����*(Dj��Z�������������s]��נT�h��1�|��zj�ּ�̧6���
%�Ù~,�i�����I"rk�,�V\ud�h�g�Z5nWN��ꍱ��؎�3�O��>J80:�ߛ�0��Oka,(�)�ԧ���r�i�3��J9�wuw U�<��J�GGI�۹��pt��
�i܉x=�wUwO�b��z,�� �ܧn6N{����}��ʏ!> /�/��Jg��H���.��_��1�����a��2��Gt��R��]k�A(Vş��s�)8D�ظ�.�:���~�24���h֋��?۱ɐp�)|��;�{�C�?
����ŏ�J*E���" HH ������7����%�g�O6?����E�������Z��X�Q*iՇ��+3;�# i =��[|�2;�;�z[�̣+��Q���'������1m�V��Y@�����c]]N��zF�,(~�YvE�װgj�j�pZ�GD7�9��M�����z�����c��!CG,���4%ҳ��'|�Z�h�f��}X���n�5�Q��)�A��P�hW���]�	r�wi�y�#��u��u�cqS�Bu�
��w�kr�<�'���2���>��$mvغ��]j��V�:od����=����-�9��'%���7�}�

 �+�����:��0�7��=U� *f�P(+�(���=ؒ����_�;�>�s�2k�7�	i���CQ�*����*jD���
��ϗF�pP
�O�Y���ď0��M��3�
@���&>Z-���i�ՆTJ��xn?I�	����J��lIK��t~!cAd⊔��v��3$ֿI���z�����T�C� %=�g�����h��@�ۺ�GE=��b�j�����ݙQ���Je��SM=5ݪE������i,e�D�u������>��p�޴4��Z1�"�˷����Si�+�>$$�ϿB���`Ö���o�󦟍g�oz�C^�����9+&-{se\e�p� J r`z��|��-���%�H��2���ά�zY
���3��}��z��)-�1Z�R�Z��%sQ�t֦k�x-���A`�`4k5Q�ЉTKrl�jy�4 bL�^ \~�z��IҝN��M��`d��F,Rf��EH@~��E�d��9y�c�eצ�̓�l��M��s���y����-���ځF�$vD�"�su�J���z�-V��!~&�^ �����T⛣�'����H��3��rR8S0��MkNt�W�"Y3 PڛM;�R���l�3㹸TX�h��8������I�z�:������R@�G>5�����ݏ��������@��b��,;�(��T�R��3�,�o�X�2��3��ӻx�о�^�b�;�E��;k�?�ܭ��kc��	��i�	֯��C�p~r�,m��p���/e���ơ^M��n���S,V���C�W'�Q(�+�aN��,���e#��d�������72���-�x���s�<׽�}\�V4�m�:5ZV�%�������o},�K�|�_�-\2���*FTET�u ���P:�nf6sD�8��ͥ�fG0�Y�������G�?�fn)l��:�ʽ��>ؿ��ơ���I{�	�:�����A�E��\��W�7��7d7E��=g=��y��W���#䶼.>��7ŦևKo3�<�����{�&ЊDMYؘ�؛[y)}�f*���w���z�(E�����Wk��rv	�p���?���y&3�wn�mж��Ӧ��+��ȏ]����d���Qc�j�0%p�]���b	%���8����ڔ�b��H��# ��X��HJBd ����fl��x��y��!j�	<:�c���)� V��{��y^! �"o�C)@�Fλ>nqk](���?/:��G�iz8#A�s�٣�z�p��o���_�����D��m�!B�j�	��"�QH�	�-�k��i���̕45:����4�@3�b�(�\m��`��v��F�v�����a�`W׀�|���+�!X�%���K�v�S_Z�y{�f"�$ɫ~�/����'an���x��oyu�U���xrjBDQ�������~�d�O��傌ur]É�����������V�0��|H�)���[)0�5��R?����e�K�2Ɗ;�[d1��6x�;�S"r�|��&t�������Z���? � �ֺUqSaydqȕ-�s���Xi�)2����~���H`:��ꐡ�.�L\�o��mM�O������=l�d�6�:u����`4z^a�f�W:"6۾	)��l��T=>9��|ap��ҫ�E{X�����R��+�@�V���v�a"�q���L��&�eU�Ĩؿ�K�'�ZG��2��l������v#���M_f�yf:ս�E �<��J)/~�˯%Q�Z�g\�d�T$L�E�#a��&٣�ϧ?
u� Ґ�E`,)ݺ�M��]�� �F�I��ņ�c�ܖe<�����J�������
0
	�c��O_Σn0�� �髩��k_9i4R�ڽRWM(�>������;H���c��(z����b�Ϛ,���~��I{)|��3�F�����g�^1�)��}��*��b�R��/2�D�ݛK]��=}#��H3��o@0-We���(L?s�D�t�N��x���L]T�z�{w����uu��WΨ����\��&.�г���x Sk�o�&���4||���_g�/��㍫hX/���C"F���1r�M3ë�wS����i-?yr6�'k�,l$�)�m������^����4Ӱ���ZgΆ�~ ����Ӿ�:��28	�IA�u�tg�
WKU�W��΃,=���8ڌ�(L���mo�׳:�W�f*�'T��Jl�]���}�bW�����e���P>���zW:��B����l
�r���;Ҋl��dM�`�N��[��8=�w��:��_�Y�R�-�#觵vf�I��`F���w:p��.�^4B��Фc�v��\XU��B��I��1�S (Z"ױj����d�b&q��� � {�&��[�Q7j:����[�~�g<g�%j�j��6�V�L��0Y6h������P����P^��Y������?���Iho>��E����f��%�Ij�9��a�N��%���4�ң�SG��Y���S5�g��e����· #H����8T6���"�k�������+;��%��O���9{%��?#�$A��o?$0p��|�uNgVb@�R��'SP~�*p�ܒ����Я����,���C�>-菼r��i�8�዆�FM�
�J
����B����F�m𞦖R���.��trёE?�.��t�?�dϯ��Bn=�ā\*�"e͞�Eƀq��b����6�18�bo�����;�*���'O��>b�[�~%�Ԩ�8��|J]@: ~���A�2�-5(u���G	 ����{�q%ǐ��Qv�c;�FS$O����*" g�f��]���a�/Cxŉ�\a�o���W��Pa��<��K����%wK��ǘ��c�Ç?_
>~+��f:&��-1�1�G7`t0R��}�$jB��h��!=�^��jy���f�9��#1�[>D����=�b"1��y��"l��\���1Js��HU��/�����Ʒ�\8���D�nyW3������D�X}��@��@�(lU�S���d\�1�3�Ȓ�;"�$�M=��Ռ�򫧀"`;yZq�c!ρ�����#g`k��~OE�ڂ������Q�_��9�I7ɣ�bo8����O>��ݕ˿�(&.��}��я�P� {��Bv��ف�۬�t��m��p�Y&��W�*���?��%�e�
��ܨ8�*���j�7Ȝ� Cn�&�,�~��.oB�+�%B/�{���/X���ߺ��2�R���H��4�-����tai�c�BR��@ݛ��H�nӷ�&�Tx� �H(��O���Rq�_[�?�Q�@n�+�������g���j��>��VX7�0�dkX���r��$ 4Q؞�ƻ���3s��k��,a��QW��t���������c�l�S|j%���ɶݼ���V��������skMt����=j��4�����Pn�k6Ϸ�I�4�Gv�V.���z�mk~\O���	�=�A:���i�x�[���ZP1z5
���0�l�a[��u�����^�z�FhKq��	=�x���G��)@z����Z}��Q�<>��?"�)Q���hҢ5�w償Q�"]t䱮��D蒟@R"$����'$$�΁���EYSSL٘�^mݬS�}��l�ΐiwm����x8>D_9V }���k�{/����dB�l7e���:��<h��X��n%�b=N�.�߆`�ະI�B�L$@]����
��G�7��LHL�#Qo�;)��ڿ~�z�(3jTw��d���o���Uj#&��]'���(��Vi҄�p���_iKe�N�� 0(ُsm�����Q�oz�/Fz81P�q�~�c�K;(6,IF����f�pJy���n�d2��d���CE�@��v E���r6�€����|RM�G;�U�~N�2m>����r�����+�&�>�d�Mh��%�J��ۿ�`a�����,�>����ھӖ�0g+���fj��T�R˫~��0�ӈ�mK�����yƴ�U$�I{�{U^G���y*����MY"�e�E�>�σ�����ޜ):i�)��zN�� j��C���?���n���V�=N�|���u��S�7do4#[GN\�<����p4i)5���;�߭7��|��k��h�3AG�E���E��:؅Ϣ!V��0�]��w̻�N.
�,a1UuJ�]p�[��\���5����$^�ɡ�hcbM�X��yL���	��R�x�5|Po	��d����F8�����WE�U����b}�v����IP�����-ǔW��}������ZaWi��]Π�w�3���9������F)y?���0̜[��~�W�C�>��wa�緂Z :`;�P�^�������*�(������i�1�ʫ[ϱ��m;��3�vtw8�4��b�D�~+�h�0e�&��4h�0��S}�����`�>���Ӣ����
��WȂ�;g���(R~c�'�����C�a��S	����Ʈ�׾L1���<j+����5�Z[�_�_GD�T,�Q����G��	}H�6h�<<:�rز�qg��u�AŪ�V�� �2���/�s���rp2���89�I���X%�I�=U�ޱX�$�藛Ȉx��eG�~�BE��;}�"�G�u8'}(^D�G��0��W u}���|��ûɕ�6}sm�k��s��#cQ�Q����'�gw��:�����pi0=i�%zr>���-�X�'X���M���h��\���#t�b
U9�#���h���jE�1P�������9��I�5� �w̖��F�j5C1�s�o�/$\A�S So*�Y����-�91�ѥ�T����4�g�g��.�z��Q["�!IK�H���� � [��������g�oȪU l�H��K����['UU�F^TJb1��f_�UEļ�����p@��^`Uz�;���Q�=l��es�w垲�ߗ� ,^X��c�b��G4d4d#>��A��"� `>�$���lAanpi�Y�y?�@���(�ʋ����Zi��6�dM@/0��Y��)#��暵��p����S��מ��:���u�9���Ӕ�GB��rs���LLL(�e�A�G�=�F�XRe�����2@V�������O�b_�=F��k�T_���1��<B��^���-�)�f������Ҷ��3і���;#�����C]���!"V�� q���L�{A��,�Y�ͥ�s����X��3�~�8�4�L���O��쓬g�E4Ny����G<UWj�@TmY$
ָ���
�oő�lk�?��Z/(��Ӕ�X5�&}�z}�'�����hZ�l�P�-�Kv���|R]��B��9r�$َ/����i�n�ŝ�q?/)�,d�(�à�o<4�\���u���i�eG����M	�2���Џ'�?VQ/ ]�I�-�����BiHܽ��7^�{(�F�����Fږ����""��]�h�#'��c_ee+�Gh�����\x��ȴ��na�u�u�)@|�N�>�>8`b�p��F)���?)Ja8!��⃀���ds��ى�M���D�Q��=0^a�|1C�R�%|�Y���&\j������KѦ�OA�+�(�&Z�U&���vȀ����R>ɯ�_c�I�c�� �s��F�?�����טX�հ���ך7�a���o�+y��_yA�������af�Wa�F�X#�}���}�/ 'a���X���bpC{���,���G�KEϲ7�*¬M�r���@gq�����aW���
6/�R2��p2�����qS��F�U�g�=��⥼�y(:	z	�u��>�#���ƕ/
~07�Y�XY�GO@��:R�޵{��%g��w�F3R!׌��t!7���o�Ն���+p*���[m��J��@"�ͮIeF�Ԋ���؎�ҝ�PD
K��T{��G	U��<���c�j%�s:ߵ❑�"n��2G@�>��m��٭ ���/�f�����5%f��6��)h#��fx#5u�3����5i���6��U��	��j��3�H�t�Ĕ��i�\��_�>�g+T��`�y�p�ػ��&�6�)����#mޕ��o�yr�@�ǘ�\�nJ�G��xn�f��7�;;13U�SP�>,��>�X��S��Şo��x�rV�K�r�Tw���z^��p�o�yy�)>C�C
`�AQ��:�Z�c��	#��%�������M�ǂ�E7&>MOxivQ�MP�����t����%��Z�p��ݍH�awf�z^�"�	��sL���7x����_�?��d3eC�)?Oa�
��q����{Eх���o��c�A���Ժb�!�3�Y���y��^��}
�i�7�R�g�K��0b���"�#(x X�E�w,&	���#�$.�Wy�����yx���r\@��w�ګ����1��ʻ��A>�̊5�r�(i"�X�eYEZ��j��%������w�>RD\v4?<���v��ؘGfo�?���Ezx�/��PB��>~����ƭ����G p~�O��ڬ���C�Y��,V��S���;�9a+��ً�.���a�̂��́�P���Z�h�+6��m��D������Q�=�yp�ê�A����K��D���R�!��t��������C�vdKs�	��A��X`"���ڏ����ro�Kx\��-oM`Vת����������}�C�.I�N�X�/?D����߿W���Qh�E-M��du1�ǉF�q��OIM��D��saC�G�X�	{�8<�Pn1�.nx ��Odh}ms�o�y����ϗ��F��f��I���Ma`֨�u�={9��v|�Q��#���oO�s��-�9����4�1��_�*�d|x�d�ǖV|�s�0!��Zh�d�(B�����OTY�"+e�_�ޖ皦7迄��;`�����Ҭ��Gj'O�B2:}�M:Gb22��*{�z>���[�J#�`�~��y\�9���¤�klX8�H�pE~���t�=��5���e��z�$6_9��R�/՗rO'�B��Y���k�sJ�O43�����w�%l!4�]������ 3�9�ȧ�����?�az� 3�џ�od���qgԿ��a��t�!��_�
 ���{�3�o�3�с���Ln��*��B�2��AFf��6����a¾���;ADVSC�ģ�&B��0iZ��	-��Q�at�g��2�(�#����?�3^e<����͞j<��҉�e������u�l�D�=����68��Wo�mх=��jCwiC�P!҄����������"JTn�`�{p�k[��<3n d�pBB��}|�4�Z
2��g�{¶����j�t��ϱ����Y˸u��Nu�t�p�s[�[U�רx>�\�b�@��A�$�p�&�mG��1b�rC������A���ZKZ�YG�՝cE�Yfi�-���k# ���HZں���[���%?(0�V�Y�z���EЀ�x. �͸�k]�F^Y�6���ݼ�03�w�f-f�w�YG��e5�)jut.>�"���TPM-�r�:���T9�$ɓWP�o��F����&��ˍhIx}1��q1���P��\�@�n�%QP�M��r�5ϯ{��X�� ��uO����\4p���֭��$V$W�+��"���}��!����}vW�f���\j8[��9m��7���1`���B��J�r[4��ρ�E{#���aP�Tu�5�^�P�?׳�����&e+a�Ы���g�_"�U�d�W���o��ؐ[Pԫ�]�D���'�	kcЪ�u��&(,h�[�+���vDk��5���֔��Θ�H��ikĆ�{Z�R��i}�Ю���fM����� 綮��������9�13�j!в����;1�C���b0��y��n��a��ھ01���7��}�V�5�oYV��N� VQ/�k�7�{N�7�w�������W�B�D�`����͙� ,�rѺ�f��2�3gC�F�C�Ā_���ۥA���/��B�6a'&�Q`BC�\8H7Hm)�dzw��������*�����.�o��C#u��aO�.���w�T5���jsg�[�WS��ˡ�_+��=ͅ,�!��l�'�y���-�c�C��<��W�2��V���w��:�����0��}�T`�8�61����L��О�^~����\�;��.��ϧ���&m�3D�:���q����f�!����)6����7YT\�`x�����6-mѰ'W{�)9�#L�!]�?[����.h9x�YBeh��3Wx�8��ਰC�terp�Mr��d��e
81R�R�,z��s�>$�m��� x*ףǤw���Hh��`��Ju�:F��D!�e�uo�9��;5�v�h�N� ��ZŶ�n{24-��(�5�[	��*�Ax��0�!^��dF��u�^�����!>�T��ko��W����0���S>���k<�6���u_�k���H�1�ߊ¾Ő���fe���n؎�	��j�Ӗ��/��&'� G����M�La��WN�u�|�P��|0]2���|�@J��"d��
ي-l���v�L�L��n�H�V47ǀ�VB��Z�^9�j�a�t���͘0IZ�X
_X�:Ĩ�5�Q���rlf������50k��cL���[G0�͕v��rV���N���v��c�Gk�G���Q(\rU�j����I/�^q��@��ې?#q
Rږ���jQ���&���J�SU(<��
z �^��'v,DRlB���ݏF!Խ$~ۗbp�O���_���Az�mCs��{��l���"�V�U����8x(\C�˄�sݣ��}� �o9�W-����c���no�V���q��\�������y�{٘�z�H]�n
UD�G(�W�(0_d-	�����d���������t��7�ʚ���+��ԓuھ���]{��=�ki�Wf<���y��~f�y(D���lovЎ�L$'��-�F}��^th4Vr�N���4���)�u)��mcY	C������j����������4HKKIJH#*�Hw#H�����0�k���k��}�����9;cu}�W�n����C��^���+��'�=��I�dZ�2+I��F��>1�(O��k+=s��O8��yl9�z	c�]�En�ẃ�QNQ1���|�
�b5�ks�2��m�VP�4��n$��¾�z'^�B�Að���䨏��[���m����]��}�[խ�{�P(�+z��XF�j�&� ��/CԵ��*u�Oo!)�~!������%+gM<��6�]���׷�I��M>�p�=�A�k�xB�fq-$g�p](�#��ɟ�����C+��,�˕�T: s5�'��e��� �ce���ZQ_a1�I��8��N��n������Z���j��o!1�Q�c� 7+�R'�4jZ����� {vFJ�B�i_����ֶ*0Z^��*�	��2�w(��c���('r��ю��<%���]�;���9���Yjdn�MD��-~�.K�A���r�9��468>a
�@�<��� ;��b��VB���ǉ�]��_��S�f��i��09v��o����i&m�x�%��{�Z�
���gS�>��"�s�O	f_����j�4�̤!�	4`��,���So�3 ����5 ������i3��\���G�npv�
��	�vܩ]d��̷\1xI���g1�I�g�_�"�r��"�HP	��YRޠL���ĉ����vwg��|X�2�+&xu$~�`p���>H-�l,�-$�F�测1��7�Qdϥ���6f�r����u�TdА����sJ���\�A}�� �#ň��ֿSݯ�f�+���7�
�K~ x�u�L6��52=��C��k�*�+	�:(���������g�Sm��s�m�!z����:g�4��É�g��2y�4Y.��+ȇ����EE�z�!ڀ�xF�G�j9
'��p��IK��=#/�ݼ�M���n�T�ᯣ�9�0�T�S
ZqETy#/G��SOS�g�3���ڸ�x\��MNW����9�bw�~\�).0�������@�<L�l|�D��")�9�yA
�X0V7ĸ�
��}�EБ���vߦ% ��N�N&L2�I�dlߚT!�ɂ�S~9���F��/D�|�[��@o(����>��wN����#��e>�~��8r�Ϸ�oܰW;5A�����g�sm�7	�a5��z ǲ�5,��$�>��(���d�Ц���6�I���M�G�;��D����C1&����5�N5�gnƎ`����Q-���^@�����,e&?�t�Kʁ.,���m݉6��]1;>I�I�GWi������#�7��ч����՝e��� Sr�*���۰����*�rg0��e�CgO+6z�
�6��C݇��dý�1iI�9G2�#DϻK3����g��<��|�T.���*,�/2	�51��}����xdu� ���Æ8�v�'�%`�?:��;]R�(@�${x�����ae����b��K>s��pU�|M��V���
/���(h����p��m��̱�=����0w�dQ��q�L�n���7�����I Ƴ�x� ��R?���.�,���8�?�'������j�`��B�ޚDo<:� ?s�Ib�ۘ]^�4W�x�������똱�sNBj��C|f@��o�b	9�U��9[���-��[Ig�XB�LU=?8�klV��h�]���ñS%za��Xz�j�K�{��{��t���xq�[����G}F�d6��u����1�7U�py�v)�"�;�w��R�
�m~<���Ydd$����+�"aŵbg������rbn�w����r�Y���O^��vh
Y)�x(i8��/h(@h�<S�Ч��b�G��V�֏%AbØ�vC_;��;��LZ��s�:�~���:u������d�=m�A��.�"���z{`��JX�V�����z�Tv� ��PxM:Pu�	��1�f�]hb�k�dv8eD�~����j3*�v�8j��؈��ǘ�[��;Os��S\?o��������X>�,O$k}?����S��QY�m�ɖ���:�Q�w�-���|�Y�z��$���f��{��Z������\hv�`Z���	FqA�Z�d�S��o���=�]>�w�izpi*\��F�%�n6"�(_��ҧ�:���6�Nk�ysG�ڪ�f�+֔DZ�����ߵ���8*�j�9�]���kT�����뎧.2in֠/^�'�*�5{�Ĉ���WSeA[��D��%�v I3���6<>��x5x��fH\��$�=��Z�D�Ѷ��o	}zr�1��>������b.�~����+�g�Y�ܦ�g�7��(�H	�w����oz���қZ�ŧ�:�z:AR���ԔJ��0#�������Z��q��x�&�O��?ޘ�����_�+�#�������~LΖ���3=u�]e�k��Y��Љoܫ�[L�vO�'��~�$c�f�Qd��|bI���vյ�㍓��b�r�0�=�|9��K|m9���MM���'�LRA��bK�d�jU�Wу������ F~�r&��V�}�����r���Ap��O�r��,s�q�7]0��k:�R�-�)�w���%��u%���G��dZ|YN%M�{%nbl�/��ԐTH��t�)'��Ԕ(!4CiW�$b?����o؁�j�WX���I��{��Uҵֆ���^7�еo� ����䔺j�-�ַ��%��4>�V4EÖ���6���v(��my���|���i����^<\?\QJ�?��*G��Eѩf~ф��lז������D2
��v�`��pҙۑ�١/q-���"[���ˆ��w�e��j_p)i��}�5�X��9iLk0�0DQF�Z�D&.]
����q#u�nv�b���P�orRvLM}*{��I۟���D�$~��[�!&��"���8|#����a�F����������Q0�z��cb~p�9�ꎗ��MkXΧlH�z&W�L����:���*�!�ʮ���3'z�i��`4���g����v�z�v6֦���N�T�-���Җc�`%]�/eb�8pf��-nկ��z~�\Cci/^v���Kq���H6)s@#§dm����m�.��h���>V<��w�M>`�6r��tm9ث�?�{��=�C�%h��|Z5k�^��;yy_�x��~�֡g��{J۱����Jx9��i|Cu
�п��O�&�r�	�:�ȫY|GA\��©��prrK'݄�jxO���(c��q�Sp�o$<dQ�Ӡ�ke�0(6��~v�`\�4�u���u���V_\�N(!�����+�O%�;�� ��5;Bu>H�����J�7v���h�x]f*�N	3�}*Ӌj��uU*�׹�
j�Dm�V	��.s��IPp���z�O!��~ʵ˳bQrt�2w����N�t�D��a?�8UhR���!�}�b�s��U�e�}�f�o�AO���<���m�W7ƣ;>�c�t]���1*.�?������e��F��e�_l$A��s$�0K����<�|��M*���UW���!ۋ�w�t7��x=><]B ��ON����|�%���v&$�j�q>X"eV1�넋6Ĳ`�+ӂx�Jn~N��[���\��&}Vj���\844B�i����(�&��3�)W�QEd�v,�^�m���4��'t(���|A)�'���+�eN�ͬc9�*4�hxj�o�Z�9��j8=hr⁋�0M?�m��rp�Vմ�oI��Rp�~y�|jiu�u�)l���u0Oѳ�R2��*f�]�I�P�`@�we��5���D4o�����7�����+��.��)#�����ž��>"��E������_A(S��Xr-�F���An��.e�Z�B�&�E�kƎ����D���q�����It�-5Q��xzPR�w{�����<5���.%������ {bE���]ks�9g�<�j��ƈ����O\I�Ir;�3�S����)�拼bGA�z�]Ȃ�)uQ�5/2�An[[UK~iQ� ~CN���,�@/k���L�W�>��믞V�q0s�ffxK��5�+	�㗡��t��	ɑ���;�7������V��&�+�S��z�?��T�ϑ�#�m�kg�C"�����yb��t헁����E��Hƣ��UkG�:}g������&^@|��+���U����)� ��V��9��&�b�q����W�x{����47�z�<�q=� ut4�u�1i��j��beJO�9H����+���"���6/�Cz��Av�_���G��W>��3��8��+Lj
PӤ�U�\fW�\o����v-5�].��y�\�挸X�;E�5��ᯕ�Cܽvk���M5X7r��dD�Z��m1����b����Y����;��1�r[�&SC���ņ|nE]r�����N���_�뮮��$7Ib����;�#q��z�
~j��vf\%��d��g�J��=�FtK_-|hIIF���p"�@I�+�d��'|j� �"�W:����,a�yRt2W�-���V���*�{ϯ���]���MnV�_��f��(]jڑh&{�MP��9�k.�"��f`�`.�*ON����u�$��ʡX)�j���|���p)@9��2�T�v�l�;��5��<Q��h���&�~�~c��q��{�i��3c}�/��{@�^{LB=+���$V�VEX�y�&u�!� ��#Y��֐��I;X=Y�&R_��?isW����Y @��s�O�#F��whf���'��H[W�T��?�9n�Yv;�A�A`pD����`Y(ym���b��>_]|��6]�Փ}����˷��?��a����1��BH��cH�Ȍ
���4R�����YM����_ψ!�К���1�W��*OW2�{+�A?k�($��G:�Q�S�����Կ'���/����)iH�l��ݰZ��"(a���|����髻���A��?��R]���]�g��@V�=�"0"��7Ӌ=�%04����f�|���mK�%K��1����CX��i�	@^~�`F�p|8�>�u�z6���,F�m���2GN\��7s]��MC�OnqP=toRV/r����*m�yBD���$~65��U�s�������B}��\AΟ��%�\�8&��	�Q4�x վ�����=��P�����������3`1��&X�\�V oj�����q����*A6��U�r ����2���!N���o�}��2������5kA���6��=�#����4=�֛-�<�RumkӷةUi�2n����M�c�c�L��$IGw�4�K���Wԍ��,�[���ڧ ��E�xj�cA݇��aIJ���*M
��x;�+ꙮ�ޚ�ň��<��<u�i�Sx�:�UWU��@�{�G(��d@�>ב)���v����S��S�����8�vk����+�b�~��=`��l��n�]��e��Ч���qr�r��L�Id����Sۉ0 �����f��K�;��d�E�#(#ц�������hc\�IDz�)[g~u=]����v�lx="&�ew%����O�ҍ]�Kψ#N{�s��:�}�v7�6
�z������>��Q����
m @�����{�r-�^MU�ѿ�0�h;��dk�C�U�ۯv4�:�/�5,A��wӣ�RS��c4wm��m���[�S�)I{=�^�	���c��3`�nN�g6��g{�4x�a6�-uL�����TIGInЮ�p�d��	��AN��צߘ(��]����O %p�ϣ�#b#>P��|5������e�nɮW�_���P[6y�R.�������L·Kզ/�}�}�ىW�W�S?=fT=14�ә�\�[��w��n����`���ٗ����Q�i�It�׽z}��@���+�@�k 5׿�������߼�\a�P~��4K���V��0 wv�;�,fvrfb�`%�D�sr�S<�>�fR��臩���5 ����9�`����!O�m�ΒΎ|��_�C�5�R�A�6	<o_+�ồz�;�qsF"d�zZO�	��U'FD�A�F����fӲ�3�	
:&�(������1ep-���Yn\��ƅ��fi���wi[Er���]���}�1��*�:&I��K��Qlr�M�L�O���7�ޝ=Ζ��_}u�Z�L�!����yC�+�j�P�"`~��S������d#7������9[Zy|e��48��y�?���&Ća531�XA�Bh���(�6H�H�\n���
�8��q�w�f\v����J��#���1�)(W��	�0g��L�1	\i�;�Uj۫83~OGg�a�A��ڀ`��`���M�V7p��%v��P-J������1k�����������1��	��IjĶ��e D���J�|�1����~u��!&�]zN|����+dfx/H�ϗ�i�!v�I���+4�;T�� 4� C��x�F�B����xy���<:s~DǍ��e*�t���� jy{7����q�<p���َ���TL-?������d�xL����A�p��ύ��z���>7���%����~������=Ʀgd����Z���-�z��~�?}.B�r����p�܍����'o��� U0������w����m�|�d�s�aƀ���}������܋$�g2#Q�e�a$����m/ 4�8�8i��>��q�fH=�{�C�;�j��J�n��%�d�O?�Pp��nV�@.��[hs^%&PB@�j�d\�H�`h��4���|J�� ��k�3�|l����#F�Τt���P�$�u���7X[�V��FX��;�,s`|]���0�Y�Ϡ�����R���t!<�H�DY/�U��sڈ�:��&��.30�0[��D�ٜ�Tm؛]@�\Ny������M���,l��[=�
:�Ѷ�T^�Fd�x�Ru
=����o��dn^D��7����Y�- ��2n�3���R����ym�֧`x+L u� $����
V�DdԀ�W��W�
¥eR�0&:��W��bfKd&{x��ș��@���"��De�"0>����~�^o1��0��n����)ej�g��ѷ�ϗm^J2 <�0N���t!8 �ǈ��$�2�*A�⿑��� Y��7���S7?S'���5� ߜ���}���>½�ߔP�U_�.S#5��n�L@��su7���Fە����I�5�[! �$=���r��AFl�s*܅i����P��_�@JH0}:z�{�J��>!:S����:��&������m�5��C�6�5L�0):�;�Y7�qp�I)I�5��� PK   �EXo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   LYEXG��<�~ H~ /   images/31827051-9966-4dbe-80e9-38f1832eb628.pngl�UP��w����;��wܝ@�����ݝa��`���n���vUw�w��TwǨ��a���  �o��    G�������D�_�qא��͒���6� @cڛ���"�� |�߄�����?���C�黋��������Dc���E�����;���ƇF���������������������(ഖ ���MZB��x���G�w�|�����*�#�C�u�%��4,+��
 ��a	��,sY'ٽ�dK�8��^_W�c$L���L@�DA4��A�$"����4�:]3��*���7��j����,�lc�>{�6�;�(�䰧����=/:�X����J��+�":�"���������M�_�Ŷ����!��2�0����w稄@�Ms���+��f=��݄�0ǜW�	�����[[3k�x=�����D��[��A��=��L���9���ڱ������)߳����s����)��0ş�[嘞��)��d��_��+c��n���G:H�f��@��a��ۉ&�	���Il��C�/�	��|ޱ�O����d������=�W	��֠ޭ�$�
���c��u$)$$��aa����V��m��	�J�<�� �����L�����f��Φv�+��꽀2hCP	�
��	������������C�z����9ǝ�c辁6�y{�6�c.�󭬡w�kC=пQ��ٔP,�5���u�uW�ҕ}���4)���Ǔv�C۱Ȗ�;���X��r��8�����'5]�l"O{�E�R_��2���V��G)z*�����,u��5:������u+v
�϶O����_���k3ܰJ �ll��^��B��_���;��w�2:�U��@����m�;cv7��DꙒ�.�zERG,6[�n)���A��� �GoG���	��2�;o>��{ߙԂ�|ȱ���ܭ(S�*��z�դ�ް���aԖ�~�n�b_�Gϻ��^�w7?k�'��4V�!C0Y1���t����neaA���V�Ss�k�Vi���;���3�1�����eȘR�h��	�nJ.27�xqhG����B!���*�x}�}�j�_?≆i�|��{��Cx�V�����to�8�~4�����c�@�
���\���RA�gefN~��{�ش��q��t�Q�x�u[�7o�S�H���B#�?/�F�tæ�B
BSn|��_N.kk���	�����Q��QWz�ۿ/Wu���,8��S���R(l�ڟ�7��ɴ��Q'V���W-W�1�΃Gk\���n���*җ^�/��G{.��.s�����w��K����%��F�|�F7�;Ǡ^E���w� ��f'�D2i;�lAB�����=P�hT�&*���p��?7�ԉ���S ������i��6���]��2*��N����v*CЏ�as&a����D���� �krY=��&gsM�7� ���4v���6��׵r�l�aVA���_�|zR�&-���RqJW_7g�zu�.p����-7�E \b��{�����k$�0���։�çK�ņ�Z��GR�� O�)'��D����t����|�f=����&b>VS��y���@�X�n�nS��>)b��0�Mчlp������C�Z�ɾ��HLq���K���Ǘ�+�@!�̭Y����7!a����~OԲ�/-��mu	��1QdS<Y={�/U�;|�F6�h"J7���9��SpXL[���~���S�|�y�վu���u?��ج�=M�F�K����XǭZ@�#mm����J\�f��:�='����������2��D��d8K=���+�g�˷�`7�C�"����Vdv�$��7�K�~OLl�4�-��C�����Ǜ���itO�Iۿx|�3P
>P�/�֫��CeeUcd�F�N�}p���zT������nf�!�+&��b����;�{3�3�#��*)+��33������/����v9�G��3���=^��=q|�Z�u�^��u*!�A(t}C��)�� �|s�m�)ԥM [\c\2��ı",mu5e$>1q4뫍���3����	0	�84:>��m�K���!�^�i��b钾+0Crt���'�H�<�=��楇Hlg����C����IV0YU�m���^S{��ϕP�)�����-��	u�����"�"��l���xRk�yU��&��� �(�y�@k� �D)�E
0G�E���R�ш�a��W�_��LM���^9:���W�7����g�Kn'u4��Y����`�QwKG<_,��e�<�$݆M��������(v�d-�ɹ����Ս������72��"�ܖ�r�� ��ꦋ���*\��'�Z+��0|�)�\�s��)��=ŭe.���k>>R=DK~����֕A6��WGJ�/����t�=�b�חio�o�T�L����
�wY�U�G����� ����O��A�������1�b�Q!�֙��ԱQ�844D���ӌ���8�!ѭQ�������Y��`�?�վ���[����As2�Q�A�b�[%�f5�Ǖ�)�
rM�"bH+
S��ְ���P5~��4-F��HO5��xG�^K����Ն�X�}M����|!r"U|�b�ڤ��z7�c(,B. ��t�KR��W[�{z�u�s%c�nĬ= ���s�v�b�΁ؓ���NM�_@]��<!��+�����n���k��Т��"d�Dl�4����ٱ��]�$~B���h]��H P��}PF�vE���Zb�c"�(�.(���ʩ]��j�0֐��i�;+�4a���dO�$��K��Fz����UFMZnX��	�U�OA�0#���P�Q�+5��D�垷�_���6�jܮ[���~c^tK�T<קCU�꾠�Mub��M�X���+����<�^@�$ �+)��l���-D�N���x)D����D!�\"R��Gu3���=ϋ(��F��)��&}��f�>�Wm��/��:4���+x���lh�$�	���C4�����n|Zi�R A�u�H8��˴��!�5�m��h&a��:��<�H�okɭ�תf{��+�'�8�_H-�.�5la�z6���u����qjO�%tv[���8Iڮ{j(T)�[�턏p�����}��*J��r�#Y
Z�:E��T���ׁma[�H�pj��8u�����%݄-4R��+nN!}��r�'U�`�Mb-ƴ����͒#���&��}V#��O�� T<������@�E�MR�N�f��M.Q���=#�����%J|��F�����ZO*;�ɀ�%'y�?6���˻j� �Pb�U+��t,2�E�]6Y�f��*��[z����K�yQeG7���x��#�l����=�)�U�.��R�	1�K<l��,W�U��n������}�_�T.X��}��!���B;����1��i�e���#	j���yys���,!�.�����u4�kn�Yz�|&,-�J&F���Wub�l{ø�}�^�I]S�܃F���aZZZ�@|mlbr�|���w/�i������X��=[�^]�wD[��wS�m��mLŊ}e	��#ґ��4�{ۯ� q|�7�����+	8������gn,,l���ͼ�Sn��t�	�ݾ��k���f}X^�\+{�@=�t˶ԑb��I��}������[�E�}��*<V0���R��$:,�%f��u��Z�ϟA�e|�����p#Isl����.�彿T�X�H��B��܅t�A��&��+69g+�͂���h�Kwڐ�������k4�Y*Rh��q�'�Iܾ`�o��W2��2����RF|1ö��k&8��"҈�����2"���w����I{b��������hɗ�l扈��68Y�b����%��r�O.4fO�r��p�N��u!nz'$QB*�:�����Ыemϸ���#Ym���ϵ�@�n4�|s^O��!�t9RqM0�ӵ@����RFv�ʗ��Z���*���V"gl�����wF��HӳN�n�/�^sK�Ml��͗6B$Aj{	|��o�a�V�
�|����K	M�M�����y�'`��ծ�t���;�h��\c�ܖQ�W^��e��%��i~�t�.�iŵ��:Ę�6b�j����!hq��9(����LOm�UwH5�l�;q�[� T,iD~�h7�����{g=qj��`����Þ�bK ؞��0t�e���r㬜e��Y����5���@�A�1�Ci�r�P�lG���r�{ |jAk;}U���X��ױjNx	.�%i��s�6w�DL	K���^r�:���ܩ��c7�y��N���b&q�W��Hh�fW"bR�V��V^���Ʌ��E_�%��j� �4����E�e�3p�u�}ELIfJrq��G㙄������O��
�z��Qf��d�6� Ty;	5�Q˗Zn�#��h+>A6�d����,`g��Qa�!�[�����R�Nu#���H�:�U�O�?=��Ϫ�D[2���7�K�[J��Ʒ^>��3����X!����*�wT�>)tI�qk �r7��m!�̌�IpsLqM����9�I��W�)z�qh�`?��.����h��Yv`�$�]��sdZ�/�&sLl��/@j� %+��G�Z�T�w����{�̣Wޏ���$oH �9?ʺ�o�Y�{�xKn�(�\'�]IUɜ��Ȧ��u�~�����d����CK.<b��k��dv�-�?���%Yj��޷��s�����=���V�����2�mPS�����eU�j,�xy��-9�19ă���Q�.�PCBH5�g+p��˵�Uc�ݠq�I޵q')��߄�$L'r��F��|VqEX��gI�+��l?��B�k�M��v>R��6U�`]���8T��)#��z^��8c���ʕ��b�1����3��D|����PI;����₸�@���G��/�9�w>$�m�/��c��1�u�Q������FZ��/�&��B���a�BDS�?s_���`E��w��j��ޖ�IA�����I�L�An\��n�If.��G|���6hv��p<C�`ۋ��3��v���u���mC�FC�� À�f�n��G�W�B�H�0)��@����Ѣq�!1� *��N�ސǕ?��:/V�ԑrU]�H��G��fc��󊸿T*��8�˳�M*�.�hs{�l4�*=8w�%�;ֵ@)��<��ywG�MFgHXF��o}���n�(�ٞ�����:�'�Ocm��G�u�b�ҋ�� jx�k����E�{sӐ�w�g7U�6�D����=<{�S_�Z��!>Bƾ
�l5���!�1�>���G��'� �w���������좔��\�S�h�[��t���R��!�5�7�m-��%�n�,�C���$�x�a�;뢛�m(��l���/��=�u4���I�A�#�N�h�I)/���j�Ƴ�%	��Vgk���n4�O�D<&U��ם^A����~�����G'�ׄv�vH ���3X�p��v��	�Hs8����J�ՉØ�`v�W���,�6�Pv��uh~���YLE)�d۹�9�1S{��x-T�r��k(�D*�����g��Xy��'m���f]tUZR#l׿=kA �vgp�T�NQȣ�Y9A�͊�k�v����y��0"ѮiyA��y��}.�%;
�4����.8�my��w�?2��.Vmf����G�f|���@���s��}u�4�����I�n��k����K8�Za��<ׁFqǣ~��<[��-m���Ɩ^+�R�s[�A6xvAw��B�l���� F
AO�Y
�O_θ���{���#i��L��t��h�C������8�e������&gD�e�@?1v��gj�7����^;P�IywZ�og���Bmώ���E+á���e���}*H����NKq~噀"�C�yl�@L�>�:��hZ�P'�Θ��D��a$Z'�R�А->��3��F/�����ח��'J���m�ִjx��md�$If}���s ��!-OX�8~��v۸�^;2S�U>ǫ��g�ۧ\N��$AQ��L�E�әTkf�2�v3Rr�6j�|�˯����RK�UW��C.0����P(�����K��g�A�5�I7��$*b������C��|�ڽ�ri��v,Q��Y4�B:�<�fl�&i�*� \�,NL�v�Y�q��ή�eԦS�#�l�>�#�g�b),���ѵ����K� #�Tb#�[�{8[�a2�ߘ݀�2�O�������C��W�K��yB ����;"_�c��b�1܇"��6�{��>�����W��8�N ���1�|��m ;�!"�H�JQSTf�K�d�X��Kq�b���B�7��'�e?L�nx�C�^ph�Q�|(M�Q���=�x��W�ɴ���(.5�(��yF�v��ro��{��F�Mb �[[��b���V*�#}8�]<�a 2j�(.��$�p�H���r�r��w+�Gk�Wd6�"�b�4�*n-��p���4O�*��t|��g��n^^��B�)�UX��q�5|���������A^�����Y����/h(�� (f�) �sng�'�lɰ^E��]��P����Xrn��q�ZH��Rc4�(���?s��
��������H�J�R�h1|�O+�30H�P�����\kˣ��m��e{���҄����E�rh+A���X�x%G�g��Y��>!i��ޠ��x�Gf�c�71���v~�Q��`�왇��uM�VS���V�#.���J�hA|�\���e�y;$�JԈz@r^o�nF�g&
l?�0�o=ͩx���z'h��1Mt�7�/�#�г�o��_�Jɝqv�E�\�/'!գ�Э�h"�~�0b�����z����ʤD�g�V�S�v��`���u�
)dObsq�k�u:!&DZi��b�E��Ǚ��~y�PUюQ����Wh�%���/*��Y��-瀯��<����;Ѥ���'�Tr��ȸ��⸞�l����J�96"w���j�X�;h� G����$Q5Ei{!o�H���b0\.<a}�G�¬�p����M�����Q�7Y
�O4�܎}�_6�.��\�`Sa%hm� '�v�
#���c�$�?���j�,A��>I6;�������!ʍ��¢X`���	��)?�'+�w�LF�lMB����~S��zs+�ͩ :�EaI�{ '�(�Pq��=���+�cyS赕o�HL�
�b\���Żҋl�*!"8g�,@L#�`�ca�70��=�;�$��w1L:�ϑ�Z�-آ��62h�Cf��/��j/�0���˹Ǩ�'�$} ��V�����'W�cD�F<�0P�("�=�e��%��T��[v�1#����B���y�Ɛ�gH�b��?`S%Q��X�T��h�hdt;(ǩj��y�!9s���y�q�H�^.�T6���W,5v�g��l�L��x��=�p]� �k�*3Qܦ%���S��/����}���2��7�1�^\\�9�Nw��2�W��ADDDL9ׯ�\T��6"��t�Ə��<�첺���S�O�&�Z�E8y���~�'5&�U������0jvTU$(�]�l� G�m�o��ҥ�����P6�n�����֮�~|j<��Ü������K��{�-����v��WJ����@�3h�	�^U�@�cN����+����ʘ4��}�r�Qv��I��A'v&~�ƶ~�l���tu-�D�-�wa񰳐q$�X���� l3�9ׂL��zU�������yĢI+��b�E����2@0�{Cˏ�[2�P��&$��{�i���(��*&�.u���
�)� �G]�Ӗ�#�Yށ�'��)	?��b�$!҅(�u�y�#I- �a��w}�,���7��:Zw���5�(�*�(���(�u��i>}:Rᢈ�`�V�J�zӟ�4�T
"�]6����ю�I���W.�(m�j��I���S]��@.�|yl}_d��G|Ƀ�@��E
����d���U�J[����� ���\�ʰ=v%2aw[�������>���Z;�}�}4�=�g�_�fZ��At���w��HgǑ�7@T�ZM"eY��N�*ai���'�(F�x��c����::��m��������.OTV��)WU�ŕ[�s�d�w��TjZِ;>���[�9"L3��ߛ��������[u�n�h�4����ںA��Vq�Sf�'X�1S���i[�؝,���9��:�%,�vx��/>�3�b	��$�:�Y����g?�=������f!�q��I���~�)����K��Yu�<޽�jQ��>Z-��0��-.�����M0Q�����aO�'��$Ol�d#��;r�=&�%aI�<��3�I�*e�0�
��r�)��y8�
01O�^�$P��N�->���&�8h��V���p ��ȋ�zP��S�o�&���!�c���7�7P�U�ȼ��ap�:����� 4��I��,>S�P��v\Z��U��/�	]��R��/``S\�9��XT9��%�=\t��p8�).��CV�*Պ�^*��QlPc��]gӦ-�j�b�J�ļ�A�L�����`M/y+���ծ���J{# Nw��2*.XLG��$%b?�S�$F��Fp>�Q�.�[��6]W�:,��n�7^j�" �^��U$d���z���+1"	�a*Ʋ�}� Oh� A;_�9����3��7���(`8�+ ��ږ����5�"��(mǴ'z��KF��zf$z��h�E��h�ؒ�؁e��lT�^�y�>� R�G܇M%t5a[sJ��S���$Bv�v����>����
̈Ͳ�"$�64�+r�>6�,U�&K�F�]>�f�_�����.u��d���9=��g)���^���!!�X���aKD�k`�`�������ӓ�t��{G��l�e�b�~�e������T`J�g�Ċ��'�P������L���h0;mn7u�lc�_uJ���^-�J��^��n�|DO�^2�4m'9�QC9�	֐^խ�������~_r7.��ex��{sS�{p�,6�"��6]����S9 B6���e�K2ã��".��d8�q�(�Xh�Kr�ōONp>k�����Q�;�(YEq	�8R�����(��d9��*CPPa[�bX��7B}�<����^Q��X�gxJ��L@
�2�����!�ۃu"{Dt�
�^ڃ#~Q��F�Kb�a�uGa �#�i[�P�3�3�8:��V&�����]L7��kF�Z������g��UB�En��F=H�z��x���&����w��N;��*��|]���)��4:#�P?�!�q���&�ct"�&��<���~۲1E�&��"[R���zE�*��gͯ��y��X`�Ro���m:�W*�l 2W��C*᭺�������b�o>��}���y�E,����*Ol6�R��}����7�6������D��-�`	����h�[^�4J%��j��@�(�������A�W�D�f��y�$<K5�����P�+�^�G���#��y~"a��$�	�D%�1wU��\ ��AxoG��N��	�������	�h���R<��=������eς̺8��ɇr�$�`�̜,�
��S����h��Ȓ��1*as:`.~���pJM�J���R����s���eD}-����p��΋na�&U��c���Y� ���0�+��� X�������9L�s�E!�&� \2���/lV`����S������7g�e��p�P�wq�l��}��E)��
�2'����Z�B����}T����]	^�9�+�jj����1X�?�u+}D�ʕU�{f~C�����/���Ff��o�K�9���=�?=�t��ŏ��CtT]��[���v���K��h{v��QH'�tF)�4�(�S��X֡�P�p�P'���_)���O��l/���Ny������/��v�s�X��_����@���eݱtI���k�����l��iØ9�Ow#&
��%�����}Ӹ�A�e�NV�缣�{�rG��r�����(��V]�4�-�uۑ�R�;&&�`wb�UT�i�Y�k"侙RGS��-g�d>��vz±��]/VK��^p�.�G]��`.��~���<F��4��~�����L�
����r&� ������5g�'Jw�[�AR��r1�Y��.[�%�	���<{(\�����2�x,q�p]R�;�%J
ȅ{3F(4�-0U��Q�t s��]<+����xe��R�����~�RE;�۶ɋE�'J��E�T�#������qfk�4j -���d�D���N�V�vu~Y4�GI��n�S¸>�X�x!Zyq+�TC�����M'��a�;�xCy_A�cQ&�ty�c��চ���a�X
���'��tǥ(�Ož��::�b��'���d��)!w-�סB)��%�ˡ������ծ�@�n�9\8|4�`-�/a2��~�KKs���r�̊?������P�|�����O�E��]��?��u0��?��܉ŽZ�}�����V�^!����qS��]+��(�8���JRDɭ�����t�6�%LB���x���5H7�rWM1��D�u�QF�kܡO=�æ�&�(#�6��+wj����ٳ��0���"���_h���7:���#�Xc��>0���}+����-G�c��'�*D�L���/�J���{� ��DB�(/�O�	]�Ye�A���,�$S|9x��YXx�C52rs���D¼@��Hm�7Ǌ#P��(s��Wش�愕`m�=�5�'Ox_��%xAA�j�$�݈_�*�	�Ľ��	11����Ջ�~]K�|-W-e^\HB�ϡ�B6⦷@�p����B�W(��\A��K���AP]O3E	^���7]� ��Cx#9�JsoAI9%��dї���i?���n9���E�
7�?�t�FD�,G��D2��r65�ܜjt"9
`",n��A�03T�˻�ۊ� k���I��u� 砟��0�I<��'W�q�����V�T����VŨ��#�9D�ze�x,�f3VB=��H����="�k[��67
�����X��Ϋ�2��׵�iZ�r
諮r�������J�J{����
�G+�]COڛs��O�:�O�mE��g;�A����b��*�1�f���=��C'�y9[��:�f��6G�8d���^�� 4Dڀ�ۏ��'���U��-��[�93U�8���˙��� �Cϲ#CU+K0�1�.6��t+1����l��	����L&>�� �]<�*��&l��t�5{t���Dլ��(��s>�j��$uI*�����w�4�h컴���h���wdTT�Z�rSb܉d���N��uK��m\�j�q��5��O�V���'�!�Bw�с�T,�̡�h�V�OCC��H����_�����L���]��=S�����2� �E��ŋ��L1X���"4qg�O���|9�,桘7w8����F��g�W^�ώ|e��>,O��$�͔r6�����t��Yq����]/������C-%��z��(�(����b��Q���'<-|7%8x��L�,?�젧��
���*L�����]�_�����ul���� %q��v�`o�q�~�@���(�\���������У���L|��Уթ�#E�S {�W�����џ��Q|��#�
��;�6p��a��H��&mE|2�RȘ�����J�	J9qz�8���8�`l�q#Si��-Y���W�1�#��jO�:�Fד�Q�=��:z�*��U.q�>�����u2I�b�c��Q?K�<:>����E������G]{�w�O�B�E�S�i�F��%�Us����4=ۧb0y��b%'#��>&R�g<��g��S�؉�`�#1p�'č��|Y����-Gȿ|�lF)���oL�q�4f�#�e\u� X-�;�M�jS�e�Y����B��'��q:��bҟa�wPp�4	xSR��c����~���Nߘ=0����}���3��rc�����*G������&O00���E����i��xtN��
�zv1Z�x��JV�g�џ2
�=T�@qSM]Û#@U�O�)��#$U��.!N����R_z�5�k����ЍB�'�/+q@�%oV����'�r����a�����[Dæ���u_S,��)��_���$�����_U/�V,��Yl*��u��1.|���ۥ��3���Y'@���2�vm��h��	J]�=|$ Ĥ`�c��	�Q�&���~N$�sgS�`
����GxYER�}��5������yi��Ļ�Η�<�o-E2T��4��P���m�J�{����ۖ��B�T�(I��ֿ{\���X�PRG�5�NEI��ｋ�N����=��uWP�7��%��ql������m��ԀU<����U ���ѡ6�ɉ��-�
�#�m�58���E(&yja���
=�S�P���m��%L@!B"Ф��<���_������)`EC3��|�1X\����䊼^_7�B$�C����fڔ�s�F�}�>4�����g��Z½�}��y ׵�I��� ���;��@^�@2�R�^so���0�?�O!(P��K�z���DA+m�A^?�b����0/��J"ߋ�e��7��Q/N�|���7��HŠ��Ur�v��
��O���IRW�7D���4H��&{��Ώa��hǃ�h�/w�Iu�U��b�nO�;o�,^:�I����U��_���J�|
vte��@��c���[y���.t7�!B���ЙQ���4�:��;��э&����L�b�����u��xK���94Cu����8k�Egpr���\#v��s TXt�ŶU=Q��>̞�G\o��%t2$V����{�J�W�p�/��|2ǁ嗓O�8u�XO��E0��F�����	W�F��s��\ 0�B*� ��y4�T	�{\��f�=F��t[��+�Ii[��M<����AI&���(gB�Z�`�:sA^��_8]�=Ufx'!�B�e'u�-~��9jդ��6�)��7�|v�*���ֶ���B�x�W�R��e��i�
����5��mZ�-B.^8�`l�ݓa|8��#��{Kť�������C��Lλa1���@D�,�����l�R���T�w+'���s����.+~^z�u��)}��!�;ggj���?"*.�Pŧ^�U�|%�4x�mI%^{*`���rVx�p�M®!�ԕ&5br0V��"G�<���J� b�*�$F�~t�t�Vrvv�����~U_~���'E`���q,��K��p��������/����=�����8Z)�vQX|rz�\};���ߨ�B�#�Y)�X����mxR۫�>ܿqͩ�!
@���9���)�O�u�fd#ܳi|ޣ�m$W��N䔛+���|���j�/�:e�O�_���f�WdG.������Y����c��l�Ŋ�.�Ĥ	L薶,�et��i��J�\��EXt^�n�y�K���)K�0���9c�9㑡B]ɝ= �um��- >�5�zv6Џ���g[^ZZ
40VAp*��sޑ\p������<-g�&[L�˱W�C+�~�r� ��M�̸~ïb�IY=�>^�WĐ��S����dv�z���Q�_)�>z�Ͻ�-/wV#Ҵ����Vz��?�y�i�;�>@��R�i�D6����Kr�59y�it&9�}r@�*��H0A�.*���8G;�3���J��|N���W�tj�uõ�q��Ƅjp�L�Ź��tٸ���uM^c�S� *U�l'�<��e�|���y�J��}�B�hf�/'���#��0v��>����}�����	�n!��nf����q�~M�"�6��*����ұ+��$�j��=9�/;C$�?�^����{� Hp����V�:�̮������	�p���e�};bw�t|�g!k�5�3B���݁y�.�w%�ݽ?%�\/+�G�*H��zP�I>�v�9^L�C_�D��~!���=�c�uV��)wz���leCm��d�*䒏�w��Ñ��уl$&!;c��#�}�L�����y��FF����S�G^��a�4�����<� �� ��k��")�;�!��_K�P/�E�'�@[�;�i�����C|K�eɵ$�q�����|��xe��s�!�L�03WV�;\=a�iD�mH�*���53�$����ԺkJ%�L�G����Vjh�������k���(?v����x1��mqqc�;I����};�����8/��V�̷�S�Ӥ\�L���?"/>��6)z"V��B��Z��/��^�K7��Kb&�ԟ��/���~����*�D\ZG�,�8�[7ms����òjԜB��̺�����)dتNM��E� &*�.����c��&��(4gE����O�CM��0�/�>�g��$�iS��gE�jFb��,,�3ǵ����FM
�QDգИ��{���1����KX��Nƚ��Q�yj��3+�H%�Q���7�yݓ%A��)��^n�Q�[�]Ͱ���i\ ۙ �,�7�̼���|�"���Ӵ�!���!��K����J\e o�0
RUU����R��Z>��T	�2�j�؟E��]e
�?ʠ��0�ٸF��r�L�tZ��s�;*erE�Xh���<^��כ�G�|�΍ы��۰�~gOT�� �%�.�Xe�������*���-:�> ���΍Z=��Ih����@��Ziՠ++���R��˙x���K�GO�����OGG�~Z&q���T�/��>��Y��&&����r6��_�a����л:�2�2��$���{��o���2��8��H��L��g٫����S�y��J�<��F�L��#o���,��g��j-C4�6���HHk�ύ��8[�z༉��۠s'�kS/�l�9�W�^�f�h�I f��d��q���>x޸���6��~���j�tl����*S��" �j���Үң��`���ed�NY���N�+:��OW���e��W�@��Y"c���'�l�ALY��U1�ha�����\�P9q�as����(�A!�6�8�`�����w���dC��D׶򟿴��Mp䵸���?|�?T�1xT��Ӷ��#,`��+����W�p4�Z��GQ$5�����'�5���Q)-�ښ)YC�θ���_�s4����9�о*��)_�t�d��J���v��Qa���6�ޟ�Hr׿���?�1��[��J��n�f��A6炕�}=���3��xm����'pyaB[�F+�/Iu�T!�7?^~�]y��£Ϲ
 �m�BE�	>ޟ�����dѕ��O�S�%\�^]l C���*��g��G�C��.��T����O# 95��X����9���F"��w�t�5�q S�X�n�G�k$z=r��~��B�9?���-��wf���ٗd����u��c;_'�O���5 a�P5!��~%���yu��p	W����.!(X�Bj��fݾ)����l���Z�+�t�F���!-ʋ?�=�u^�y��j��RX�7��)��]6@��=[��$( ob>���v>�B �m��;�GpI���p"���۾��_��$o����<�U�����$��8zGw�咤��\
�Ѧ�׳�������K������qU�t0xn�:L��}��4ͭ ЏD������D����	���ܐv�:a����5E���O�.�:�g��|"����n1|���ֹ,J�Nju:L��^���{�-O��^Ői�ӳv&�2�'���t��+��v��*��Ab<��P�v����&��|6��uXJC��\�ӟ�e���vnm�)/�b!bW����-�vp�?Ⱔ�^6�9Y���eb������3�E
6��$�tyS �V��p5��ɚ�޺�E�2����*�~�҆o#f#�5��
��
��v��>c)�*��in�%�M=�<�]r����6%�J;��vx�:s�.$⯷lҧ� �B��ӭ7���,�D�q08h^������z�ᜏ�[��V�kBqh4�P�? @��O<��/e�gd�D+@�r�Rfy�ý���� ��� n�@��SY��`�2���FMf���[����d(7��,��U䞸t����<�٢��1dʯ�(`P���@�!�+�|�K�vx� ��F�	�&��͓��ͣ1VR�5g#�ݳ���� 嬧��T:9_���Ef�^�Lu��"eT}��&n��T��tK4@&R�Ux_�.8��L*��S�ܒm��E8��p뢔{����b�8<'iAdw5؎��R1�O�&�5�娍�J�58lf^��ݬo��u��*��������6)��(��Շ��~3���<B�uşuL_+����aAo^�wn�B��p���P���s�M���E�l�"Pn@��尘��S��=��Ie�O��c�O�&}i�`�y+���{)�_�7�ߊ�W�s����9��z2��|�r�Z�������$w1���9~�t�tE��{4Μ:(B�Q�&�����ޣ(��V�"���˻�J%~��������I(o�hPRi�T�9Y-�`�k��t�17ĸ�C��k�E7OW�U��k��T�����?;��{_;v"8zd��
b�ha�ٍ!���
fr��e`�3\b�rk7Ϲ'K�n C6�,*������J�1�!�2�7�s��Lhg��|�����)��ߧ�x2�z��x�٧`j	:ʭa[\^JF�F�9b#�5vG�t)s-Y�m�i1Q��2�buA�p?��
0��%�z���y��#�Yˮ|���R�<z�����4���+���
Ep�P|HEF�U2��7��H���h��B�&�hi�ݏ� C��R`��G���3$pqr��r�h�:���O�s�=�<�p>�H���A��`(�8�e�p:��X��'c��
nu�#�'W�~t�dS���(�y��g��i���Ƶkq�
פ��C!�C@���.�ۆ�R�Rf���t�8����x{MJ:��w����Y�F�B)��n݊7��n�[o��1�Ν;��O������AʺG���T�>N�N�Q�B3	+;:3�anF��8�7�+h���0� ��0>x�;��K�?�o�3O>��Bv�1�LE��M���Lef�#;8T�`�X^��v��;s�t<��3�ϧM�::�ls&���Q��ư����_�@]eBSY��/���[G��ў*9�j����VȞ}�{[tut�
W��`(��94C�:
�����.��<��c���ٟƋ�|����G>���������5f]��QLG��~V�\�S� �@�$����\�3i��V����B~hCsa��%�d����E��ب�m}}�� m�g��bsT��9Ǎ�0��1�o��o�D�H��x�S�mmA���ހ���[^�Pp��׼)@�H(�nE�?�,�?�%*J�M#�Z�	yװ�=N�(�Yχ
�pR���y:.>|�:�J�ueK���ZN2*������pZ�k=�x*���Z��aL��<�����T3��s�?���ҋ/Ĵ.(ngh���lx���]iJ�������ĮXujj���l���>��B}pZD��ܾ7o�(d�sqd.
�4��w}uA#WS�����/PdW(V��i;��o��u+����D	a­�}�ߍy�*x(����}�S(�f�4,Ɖ|샖��s��l�����b����# ��qU5J2�1V���h -�IQ�SӸ����}����ajU ���<��t����\��tQ���Pc	92D��W7}�55,����(�$��Z�'���>��vT�1�M���ʢ���Ͽ�L�ps��W=&Ǝ�m����8V�(�#��I�c3��z���B>�k�>G��ƹ3���������,��O�'c�����F�}&��M�h����]����`ᶭK`������h�Q=V�<�{����]`I�}�E�(��n��'yQ�R�Nm3s�9��I����˛��uD�}�@p�Dw��H���4O�g�(���LN�8�R��Bk�)�v�E�yK>�[�u��	F��b����C��i���-H��PcU��Z��0�o��O>��j��R��(`�S�വ3#i��%�9�A;ϱ�77O�s��N,�,e=]�ϙ�����@¡i܋1�o��#�h��梽��ͅ�u���}���2��
���dE�N��XR�qhR������W���\�GA��*��Z.��₾t�8��������o�;�}���9*�q���a���>P���R��cANd��Ly=�;#�iv7o�Jn��9�%� 	�(�n�C�9�Ȳ`��J.{ k0�J�i_��"p����O�+
š��������"�d��@h����&�8D]��ի�ܻ'nߘ�����t������2�o?�{�X�{�ő���'�^ZX�{w�!��)���6�S��s) ��w�c�����l�R/,����E�3A�S��^Wn��a*�K,��vr�b����AD���]�� R�+��lNJ�W3=�
��2�8�\�Z4�:��S��l�)�z7�m]T�[�iA�	^Ш�ׯt.� 2�n�w��#��AQ�|��s4 N�p���@"q�N��$��"0.l��WF@\�B��lH����ky��8�������׾o��f>��ɓ��mw��a7�m��5��B���]������X;���:�B�M"��	��Lz�}ܻ{��+���Vv������И�ȼ��Pv����Q��-��9R�[cL���AH���+k�==�eT`��5�I�!��jo�\��(��N@rqf�]]���7�]Ơ�)t2=]^�e[�K�X�byI�>3Oą�2֥��j��F�ω��o_���y+�mo�n��������˨LZ�m kf��+c὞�5�ޥ'�]g��J�4�r�
�.��ȐC��#�����`�+k)�WP9h��]��rh(�_�����׮݌�7�R�f�)��6}q��`}�Wd��܋w.]�w/_�7�~'˫q6�#'�RsUԭ�3�+2n��gOZ/�a7^i����Vy��sT=T�u�̴Ր�(u_c��	����?梼�H��DA��v�CIcc����N������[!���4���n=�
Y )�6������ �3P�����ZG��Xy�]���
�x�q)%6Ҝ�b��%^E��	�KW���Z��>�B}��
�p%Vw�C����61�Џ�$3�?7��wtt
;
���C�dbfz۩��>�޶e>���M�R	#��q��ĤՔ՘�s5aH�����l����c�MN���3q����X���H�si���tbv�Q܊����+딗v��7\S�+�r�Ҡ�,pmc=���%�K\�^ ��¾h2����Z�LRv���c����>^��~=q��d2G�t]2���'*���v�����#��a������{(���{X!���2K�����p�̟�p�����.�CE#��Z��Q1���I\�q�ٵ�MZ����n+0��7oƕK����k�(m�y��嗿���M\��n�̃�@.�&�ⱇ�hf����-sa0<���-{��rh��Q3Ν>��v�2��g��o�HuGr��+�|Av�!�m���BV���*ӗ��u_�+���dZn��`���Ay���Gr��@(7)^ހ�kv��ni-�&��=e:��5\3a qH/BCI�L*�5��\,'�9�m�Y������ ��" ��x�w��N2��28訏�tt��3��8J�58^�3FL��� fd|4˴���%\C8�$#r˔d�%�q��`E�
`��x_�A�ru��uq�CG9����ԙS��ǋ/���7��
g�Uj��p|Z_��Y�UI��_��B ]�(���b���L�2� %���xs�v�L�R@q��ԹH��h����\?�Tw�,Zsw'Щ��WG�T5˨�����n��m�u/�OR^�'����?�W�x�v��9��//�*bʜ®��Q4--
R�~�>�Z��vc(��������L(s��d����ɴu�3��W�2K3S�Z�9���z�\����X������v�Յ�~�r��ͯ$_�kW�fv�#@N%qݔ�G'�쩣�$BdrZ�� �\ T.�X�(�6m�N�'����R�G`����b� ߧ�20��g��{���֡����,�b�pAD#���u_?� ®��R<8��cܻ�65��N/
P�P~>�����:	(u*���H 	܊�����4v]S�o�0kI�e�������v��F�q��U&�.������2u�$�Њ�+��m ���[ ��+�Z����,�x������At��D �s�O`^�	M<\��@��}}T�Ǥ0:ɑ�=�:��^|�|<�����^��g�&xv#�N3��3^�`B���rZ;S�gg�p1|d���~hq]{$�6u��	X��L�/m������2��A��/�_�4��ҐZ=���$�.�&��C�dSP��kj-�� ����ZƱ2c�K7��m�v5n޸cZ��^��X�����6X&��V�s�{(#>rS%5�W�(�8��l����ph�3H|�uֵqii���Y[����XXZ������e[䳣P9BB���22�<0
�[&���i��32hl�G�f��ң��F,�ݎ��;�S��I�IB	����ųe&��0��v/�9�#�@��E)N1\
�A}��b4K��^�z�H�!�Pi�*�jxJeS|pWwݒ(n�v�h'��8�;���.��੺*`E��
 ).�ZK��[�����)nln�T͖���QP�uj�������;ռ����eQ]{�P��EY._ ��l�Z6�Ct����ZB�n�2��[Y]F���w�g ё�b��lOJ���G�'a)c9B��2	�\L�w譃{� �� Y$�9�l7�V��t)�Dc-�{99Jdz�,H*4v��6��QXY^�Z�I��w7�廓��q,��yc�\s��a�2�K�� 
����6�k!(6�g��G ��<2wى���j��6�l?���D��(���f
��`���!X�0�G���kkE P�sd���tG�hkc3����U& �8��n�C2�M���s���� z����zh�uTJ�+�S�h�S��Oi@tN�>GqÔ�\iyQ|�����٤�� N�y,�{��x��GSƌ{��N��	{;O���k�P�y��K����j���%'R��~��ZN�j��V��C��A�\�
�P�zm PhS�������!d��ڗ�N�	�}�A2�yn���iMPB�����K.�䃬��l��;6�W��!s�;��S�����*2��8�F{���F�������`�"��7!��B/0�ꕴ���b��X� uzy-ʦ���0k�tq�!��=�����0���	��0CJ�ݿ+Xi��E�P���U[�tr^_LL�:��\r�R!,Eɇ�c���Qn�Q'W��G(q�聤�>�����x��w��wގ��n!T�����Vr1��	�
��ڤ.>T�L����͍�`fj��º.���֫�3;H���g��O���ǎ�p}�XV'6�_˅+� �P�r�V�xC7�C��ҳ�sq���Xk�sN���^���!\@cX�}���{��q$��ƭ�4	:Ȓ#I5�|_~�zO�B���A��{�A���'�����|����ݷ�̀���������G����'���F�qX��u5f�g��b���e}�����Uv#菍�ǹ����S��31���L�RIp����L�p!�v	��|�h}�g&k�?Ԥ�V?�;cP�@}��^	@�E��\�Q5r�.�)���D)s�1S��9�65>�=r1�8q��r8�3�M�sB������k�	�>�=qA��Ƿ����2�D�I�}��6�@�ݐ�&8�l���1��"ˍ��+��91@m�~��xg��$�l}d�Ɂ.��D6� �{�:�?g�>�DA��޾y��fܿ�[-}b|<:f�5z]ǡ���hl�i:S�S��=��Ԍ�j+V�b&���s�'�-.��6�r=,�
	+q����S'�.ĝX]�C��?���^g[�``p�ӽ�������Z���F��"�l5�����;��[���o���z;�7�106g.>GQ&gR���4
Z�Z���\Y�Z�~�P��j)�}hh���*��ӎV����w�G�:6�wL��w޻wfWs�^�i�`�p2O�|p�b �� �J�";[�CZ�7SGF�:��y�ܷ�pw2��������Y�M Jf�5����>u ��P�A@olr,&�G��bsdx"��O�Pe*֗����_�,Efj�-]e���M���m�H�R&ū�ʀ.�,&R���nm#�4)1�B&��p����,��5�l�/�Jw�D��H�6���+�Y�	���mJ�luy�}�v\�z?���z��|%����>|6��<=��;~>Z���Ħ!sR�F��q�2��A��&6�@B�S�р��9��<��X�@at+���ҕr9�7:��1����`�1�%]�ckKo��v��]�.v(��RS7(��$
q!�s�F\�x_zd*��i��
��^�����P�Y�l�T-����sD�pf���E�~R_�zE�◾�矍��x-��.��5���2
@�|�J�w���r=旯���K1�x5�6�&�qdb=��u���c!n�;�ȅGr�VW����9l�4����Y��(&��T�v-����XH	�;mhVP}t�m�^s���o���?�W��e jߺ��H���ч±�����S�  �5:(����G�[�(�:�����L�����h��o-�zs)�߽o��z,�o�'w�D�Nӛ� ��^
�@�2 |۝=ʻ�k �>��cWV��pf\Fa���,��L���������;�'���K���L�����˸a��v�ҽK'N��FA�����������JX^]�a[`�]P?V+q���h�"���>of����p�t%|ԧ�1m�@� ż��ȶS�����!١}7i��\��l���}z�C�,���>�e%.���C;������ؤ�=u�FJ���j�fO�O X�\���� ���Ut�����dڄ�x��2�=�����)tw�����Ԝ�!�{N�ZW��z�1tK���:��e!��l��6��l�/Uj�؃3�.ML���l����U�=�ȏ�C��+��yz^;��A�l�a�� '~�Eʮ�����Z�#.]�7oߊ�wn�z3�P:��m�w� ;U��K ����ma ��E� �7J�L�7>Td�2����~8n����"C(��.o��͑�&���+J�o��(�K�����H�`�ٝ
��}�V��ko�׿�J���;44,��[���c���މ��zT��6��;კ|Қ�|�k�|��C 7k����#kX�\���y5����Bn�e�\AW���;d�2 ��Mƹ3����Ӏ��XL{?n^�ׯ��n]%Wd3&Q��Z<���3��Anݾ���-!�&.�"�q������Z,�/���m��:�Gfp�N�H�t�ౣ3 �|� ���!N43P�ZB}AA���-��;��e#]�<$:�pE�@�;  7a-�W���� z괰 K\�(��|�2�}h��i�c�[MMM����25@=+&����p�Ǧ�pguD&�����V+����!�d���YC � ���0ʝ�~a���35�k��P.,Am�R�NE0�:����ig�C�t3e]�ו�n��5�n]�ɥ T4}�����+��,�ߵF=�*���0~/!GA(���
QlE%��]��'�7�Da�-ͧ@>����(�"����"}v���c��>!�s�w޽o�s��ht�����ϒd���q�N��W�e��ؽ�K�[�A܍��8�w!�⼁X_]����XYƢ�wcc��B/�2Vy����
IAnf��U��P?���t&��B�6�����R�#p���1��R�c&�9(��_�!Y�G���IG�6������'�׎:���W㕗_E�c~~en���f� J�6n�M�h�J�r��q��)�2K#�6�#G���:�cಜ��7������t�����\�Z8�c��3]�sU�"�fVs<�x-��:�._�/�/ E����D�v�0l�ڸ�����W�����i���$��8;։�i)�M�2�L+nB��:>���-3�U8G�-c�+�5���^x��ޣ�}a�	PqO�J̭4c���#4� �p} �{��d���kw`�k��ƅ��3� �P����m�L1D��*�?�+?�Z���L0\F�W�2�粒��o���Z�& .\��NN�ə��`3�tA$�}��a��q	K�����[�t8��OW�@�1��@A�
.��eyk�1|�3dn�~��$��$@���R{h<!݀�D$��Wݳ�a�ɋ1=ZI�D�~�*@r5*U����n��Ȳ�5�[�8E�d0"����t��|����H6
��%��aAv�1$��g>�����g�]p�6� ��.��� As\�\��A�]�ue1p�/���Œ����/��Ш�:��mg3i��:�4�`��9����e����wM������L�?qU26gdp���p�N�=�v���wwa;��9%�&5��ֲ�T��]`� �r�{�>@�aY^[N��3��Q��"/���^#c[�����Zo3Jex����8��� >��d6H~�䙸u�^��o�vܽ?����n�X^��,md�ŧ㕐���0��@1��QplQG�U���Bŵu]_V��$#�UUE꫆ �oʛ#oZv��
��H�O+p��ɉ�8�b��S�F��Fb����p����f;��h�َ��923\�X3�����Z��\p�t������ !�+cGPv�7��a/����>�N#�ȧ�;��/�����1����1����ϟ��GhK�	�:����.�T��Q\P��j����Ĳ�Z:
�.�?qR�Tyw�#�$�������+<(��Y��~(�T���{� ��4�A�1�cm���Z|w�X��X���,�"ʴ��28��_ۏ����,aM�pw_��� ΋Y����ǥK7���٨�@���W.Ǎ���r:�gc7����z�����~���z��P�~@w�2R���P�~���m(�fÇ�S������p���Wr�Kkؿ(�A��GX�h@�WRy�^�o�{).]����mT�lF�� Ԉv¢��6��-��eXǍ+����q���K��n� +����|���Bi����Q�����r4��A��U��C}�����\�u齸z�@��]@�����@$0�ͪܤ�#��iw�ާ��$��������9)���*ܺ;�ǟ�W_'6�|��w��g\9@� 3�2x-�A~�I�����Q�~�^���؃96��m\��X�~Z�����G{�Ֆ����0��s�|D�Y�'���S���f$/,b `W{ A���z;���b�z�U+ ��e4d2�> �0��I��wL�{"�9j�1���{�hK����i���d�4��)��	y�̉�֨[�g���x�q�-y�DN2u�\�P'�w�w�d"I�騛ׯgJ�6~oq%٢ Zp'j9�ӕ��X��)"B�𐝰u/�>
nL%}-:��BT��{8�N
%�P89�"�H�74��N��Ǉ?�X��V�/�|�R�{�2�JwK�_X�Fc񌇘��8x����ڶ�ׯ�!.�S�,�e1�m�ie�5��k�"�\��Ba�v�>�>��P&�Ia-:;��X�~�m�̮k孿V��ɺ*�);>��v,b;��"[�`dή�7wq�Fs�)eҜ�p�=G��6n0W�ﭴ��uie-޻t-�U����q!����ѓG�G�Eu��=ꐯml�ڟ.�u�m�ڂ�9
��Zp�����Y���i�&�eF1��K{X�j���6�� Ժ���z���������X�0��ê��X{D���!�Y�P��_�����['�iX�	X����c��@���@AU��f�
��/Ga��e����c�O"39=<4L�j� �2��6 ��?�՗��w�!�#��L�ޠ����������a�� ޹r+��o�~�:i4��1N��V�����x��W]Vf���Ϻ?E���P�,EK70�u�ˋ^��C����b̞~�t��G�^3��,i�����~.�G�~f]./bɱz[{���w���/G'�S߱>Vֹ������4���B���# V2��
����"�`�,E�ԔPXݏ"���@{ߕ�\[���?ǧ� �bg~�7sY?5DaɆ${����
;#U&�AY�ؤ�4��x�A��Q�k��b��2Ww��`��7�������򥵣㤻Yk���$���
W��iC�"�����}Ƶ�d*�pC)q�AHu"�O��l7���O)�C�
;j���/����]%�㽞t{�~��o��F(�BPD֪�J�\��ɣ16�+Q�f�>�m_VPj�Z6���p�"�,c2��,M�7+��8���QZ4��=�/����{-YN��t٠n}䲁밒o��f���7�}�-	\\q��Pv ��xP��������B~� 8��a�-�B���z��rԂ�ȣ�yM��bvu�h��;���9'NP3m�X9�yM�-���T�q���ҫ��۷�E�\���:��A��;��$t�+z��Ή�Q�s�f�.5`*��t�%5��B�
{~X�g?P��/48�c�{��8� e=�] �9j28��(��5S�l�g&=�ș��%�6@�9�v�g�Z�� Dx�
��9�
�}o	wG�viT���֒Q8�ec��Q����UG�(�t���ZA�s9��y�%�����vx�C#9�P��Re�����_|&N͌��I��}�&��S�����zP���S�]��ӣ� �~qf~��H�Eu}o�ɩ�>�aee�pQ"�3E{�q��t�E���E]/{���ͩ�+����^�z+�6:�H�S�*�2v�
	[��k(}�hѩ�l/۰b�c}o�=�b{--�tZK���Q��;P��޺��-�!(�FkkL�P�>��C�ҏ��aexJ9B����Ph@#6�[�z�瘢��c��K�9�z
h���?Q�2
#QHB!�Z`���r������63����p5�h+�/0.���}�[6"@��ߗ����5H�2�>禄nS�-�>�,�u�!z�T�
F(�V�Gn[$�F�s�p]]��}3`���%�m���߿�SFF�މ{��.��T��>���"�oN/0�o(�L�����qdf�:����UÀ��J����L�����;E'Y�� -�~ߍ�����nC�q��|�*S�iΖ��l����k1^+�c���1�	&R0��1%]�� DR �$.}����3�t�>S8]%I�����)4�,�"���A���YT�H%B���(��s��g���D�!�+�K]W����ë�M%�vݺ��s3+l ��W;����_��g�蟯�LrU2?i�Z�;�#*�O��z6���f� ��z����,!.̺�A�!��*��![�v�hA���TF�65��)��qm؜ヒ	�*�
�A<��6��^��U���
�E �&H�2�ƣ�H���du�Ѭ���� _����uʾNq0 ����7%,c�@-G���Ϻ�=�����<Tt�E:m֤C�
u>D�>Hd��w��B��mh`�:;�x�U�+f�Jŵ}�C��1�~\�v��z_z���j�,��B�q!a�v��	��2��K7(�6��v7��C���d���ً\����6�G���_�;�|���V܌Z�i��}ך��H.L�5���r��	 �>oll�� ����`�0�22G��h�]�©����2��v�]�K�='�IP�|�Vܼ��PR�$���� �N��_��g��dȶr��«Afϕi��Á̆�X�c>4@�5�} ������13QEO}��p2�n���; �+�(�6���"J�%����-����0�Eu���x>�D�*_��\��Y�*r����i�8�"�`���E��¥���ۥ�}��V�,Yc!��(�����@|����ȸ�Y�aw��/�k�|%짃��2�U�R�:�z�&�oue_�D3;�'���I�v���z��N�豳l���՘�[
�\�ev���k�4ڧ�;7a7��.�_�;~d2�p&�%�m)��/Y	��.*֎cL�7v�����2�k'�`aUf��u�����>���X��db�o�Ƶ�7�ޝ�9�$@�X:G�t��u��9r�ϡ!YM��Js����2e�7�A�v�u���IQ�92T�٘��hs/Z͍\�@E�Y��
�g�d<- W�<�{wf���q��}���v 3h�{.:��\MߌiGhwe�`���;�6�j�0@�����9sU����݋��V�6V�1U0zԹE���ڥ����ќ�]��Ӈ�4T���`��D���S{�\�q9;ݙ��2}�׽'l�6��n�ə�x���F�ʍ�v{>��AV�٪8�X� d E�@׵ c?��7	��%�A{eyy�K泩k�穧�9,��Q��Ow��F&��Lw��-�O9��DLZDt_Z ꥛���"@��(%*t�N���;(�,b��&R"���Z���*�_�O��f�`o�e��t:�����|�~ӝ����8
����[o^��m[�"�Nt,����o4�h�.����52���,�Nl��:����,�H��3�Ɔk:l�q���E�����8w�X�=y4N��'�Ν��'���*���q�đ,��fn�yi{���԰L�Ǆ$�+눗���ۭFl�^��5�_�O�ݫ��.��
m>��տ��E�ʕ�3n��^�p����c���92�:�߷�sX� �F5k��͜�b&>Qv�ԇe��9Bg|����V���mM��~��Ŗ��xh��J�@^\\�	}w}|߭�,���*�����}m!K�hm
J��� �d�<�K��2R�ڬ���yyu�����|�_�lo��W�o��Ã1A[�ʰ�h�:��B�60@.d��V��WD7o�%)�!qh[Yqm�)����V��Hn7��̻�V�зG���{��3��l~'޹|#.ߜ��2�}P����P�C��o����[7<�M�İ@���k��3��H��k�h��G������8>���x "�<R���0v��_]܈k��A�cy����_���w?R?�7L�_O��|CXYg���԰Opǅ��ނ*�-��B�:�@�mP�`%@�h,-��!HTզP6�����Cޱ|��d�'��ه������?��+���S�.g_�P2�����J�}������n �������X�a�:J�0`��Fa���hx=W�6{�!@CwE`�]�Ƈa/�h���wt��4��{/A�r�-ba�-	F�u�(��ڰ������"X��p='���Y֎q �op�U�8�����+��X �G�0r���<��dd����mc
f���(/J�iurqbW���H��e��m 0&�� -��+�e>�J9:2��[V]
@O�pm�>��@��'>��8VR�,W�n𪋥��w����h�����N��VE�@��,���5]�ѕ�ڴ��5pG''p�`9���F`�m;v��ڃ1R_#�+� �V#F�BA���T@�R|��	�>�D�If�<�����~�Ñ�������f�niJug�a���G?�R�9n"�.e܏���/��|��(է���<��maB���+��������
��� �*9�@;0���5Vh��k�Ɲv��x������G���~+|��|��t� 2)n߸z�D�����g�~)G��W2>��C�&��@m��j�X�!@�=���;�,]�	x2n�m�u;�Fg�w��~|W�tЎ'�������x����	*"�{=���9���Qwgc�����Rh�P�4�&(��g;a���Bn��2\2&���(��B<�f�f�C��_�r��q����P[���b�$��	H��C0��@���p��¢�b���T�����p;cX�p�s9�X�A�QgW�
�h�\�0����Z��"���B��'��C��"�jj�t�6a����ڲ-A�,��l�@��F^[�I9q�ET�����&�:�$5��.��ï(M���k���o��ȑ����J��?��4�Vpq]��5K�Ռ��O�H�r��~��s�k�c=���C<���p&N��6t�e�^ör8�AD�~��aogpS�؀q�kRZ�T� ����Ž��tF��.r�9�A�R�yAPk����; ��z �y�[:~t
�aq�4�����[�r�Gc������:��YW]��,|w�w7��9p�{	�+A�o��p��J��
�ѯ��pw@��'�����♋��* �.��V�%h��m
����C�g�j�'>��7���v���c�ܣ�[4P_
PepW�F�_�s�	�D{v-�L��1��}��V¹$�t�cӓ���h,�B�a=Li�����'.����?O��ZB��R��Bd͇p���{��t�ںP4'{��9��"��(���b�(�	)��M�vR���j]΋�/ae���(��>�;�� ��}Ȉ�� (���Kw�ѭ���B�{�'��%�,a�1-%�骸%s��s��'Vp��2��n�o�� p����d^� ��`���r��B�Z&�{\O��zN��7hG��a����k�sXS���*�Bu?+���N�0k?��)=�3]�.5}�dԇe�����.��^�GUXz�y�v��䦀� ���X�\N��2x߃K��`, G� kOe ]
�mkWp�_�fR]OO1wI���v��˶�5]�HQ��[��B��#�G)gA��Nᇽ��e��pbc��}��_Y`�k��^��џ� =����׿��K��J)�j8e�(���}n�����ʲ#�CQ����� �H�2��"���835��_��x��hDs>Μ9�l�I�^K6m߻%�(� u����/�}����r�`��]�V4�%�C�f4�t�@�`�W�S�PS~���0�x3(g V&��4�����N��րN���`��s}� ����#��j/�8�̺>����>�v ���2���`:�����k�>�W�����Rl����N$�GC��Ŵ~����ޥ\FH��cF2N`B^
8
apM���-����������U�� �Zs��_��*Q���(9��nN�-�q�#PE�s�;ѕ�s��#��Kq_'����?e�5�Ne~	e(��r((��]�Q1l?�3Gh\��66 ���#�8��2�C��-�)�g�y/�%�Rv��CֱC"[����>� 3�Q8j�~>�7��������sSd�>�����ip�2;�f�[Ȯ3��A��DY\�S/��]{��t���>�ȶ�Ĵ�@b�{ ��}��ϔ�M;���KN�=J7H���=�
���V��ٹ����l����h�c[���BQg۽��gK��pnI)uA��D��!��t�Pν=t���G��o����C�c��gq��7�Ӝ耵ɭ ʸ��wo�H)���^�_��/�Au���#Ai���f�Z�&?��;���LՊWA�}���f��3"�NDG)��4�@'l:掠��ȩcS�w�ퟋ��gc���"��r73�'"mǢ �t� �S�k�b�aN��}/�H��ź�Sv�CG<���X�##N���6�7R`�\��̦�Y.��l�q�p7I�E�Sav.��}j��҇��ΌǤ[����H�AP!,���T���j�3@��.%�B��¢�PPۯ���S8 ;wG�Q�������9\���e������ ����d?�'�0 �BQw�á���ferb*�kL8:��e�*�� ��d��F#"X[/] 3@̿݅� ��% ��i/��@I�����Ṕ�V�sp�ɕ�&�:FJ���a���
ݥd������@��p��^�@.���&LZS�I�g,�A�ס��U���r�`wD2'����f̚F�0f���*�Eݷ��F��P�@=d� 7_�
��ĝ0�|��R4:�ƫ-�E�հLJ�_
D�� ^DJqt�'~�~8^z�XL�%AU�8}��R	$�Ƚ;s1{�N {���\�_��/�:����+Uw����)16�;�PwXWEP��W�Pu�Z�޶�9�Y�5RoŤ�.7W�bp9���ʀ�� T��Oŏ}�Cqrz4Q �e���[-\+v�bc����AVu�������:���E�2z��K#�270ZM��c�p%�j5Tl�n��w�7k+��~��=^6��h��%W�Bh�ݻO'F�]�/����T^����Rӱ;\�9?����m��q�L$��Av E�P+,$%�Z(B��f_�<`G��r��m���f�+#�����W�e/Zj��`��óEއ}���p8]W��������9ʫ2�"��FU�A�\�ʠ�]�^]�!]>E�W����&Zr���e���.� h@��*h$&O�s䰶�+��
	z�����DR6e�E��2،�M䜺��hY�+��D�\�Y;���,X��V#�ߺ�k��s�����~zX"R>bC�'����۵p��u��2cX����n�����*)/� ����ρH��O[ ����v�+����ŋ�H&r��Lc�?e��ϒ�&�p�[����콂&��⫯߈����"m־�4�jOlmn$��s�N�JPH/�>P`�K,跣"#(�X[^��s	 
l�6d���C異�c;F/�l�6c_��щ\��� �ض��?�Qxp����E��Q����8ur&��kԹ���8R�-l���Ak'�s�ܶ-�"��7 aS���>6�*����6�3��ǎN�p�L}��z��h���D����@���"�1?7��я��B���Bb
�e�9?ϽƠ{�h��(�'}�ڤ����9��4)�V��Ԣ,C��S<d�Zr�H@�,����A0ʇ��$�!�S�C�J��R0w��pup�xߍ���v�U���֭=��+l9�rSm��Y��	X3��)pN�W&���1d���n�h9���R%cK����� ���o�!���b-�̙o�u����_��Q�r�$�J&�������:���.��^��c/�4��BL.u��l,��F�cA�s�m��E�	�� �%�Ps�"S�ے �9.�-h;�T��4u�����?�D$@DЦ�r�����$��x$��Wcbb4W����)3�l l扰9�� ��T�;s��ƥ�P2:�N�ʘ,S�:�Q���X��K����+\�����
f��66���*���1 ��� i������30#��m��:�s!Ui�yE���͸v�ṋ������5��ifJs]��r��:}(��RS�[˺�2>�
 ��ڍ��F̯l�`�k�[�������&�^��k1��0�&º��+0��>��6��������Y5*�
,�(h�n-�͍{s9�3P<'fѪ�+I����VXs�]<��l3i�'�a��u[���}���ُ&�;O�[���6@d�)��Z�Ƶ;�(Ꭻ���l"k\o��a����U��s�&���y~^���[��mq�E�E�Fx��ǚ1j��F��$�֫	@lR9�)\]�Cs p� Om*�渶 H�8R�)+J���W�ʑ'�ȾVN<p$�X���ǒ�F{Q��H\��%�����N;yo�����|�G�Ǒ<�ݾ���U%u�@-�e]]>��֌Q)�d� ,�r���,n� ~QÓ�HQ��)AU%j˺h'�G���7O�~jdrWةA�p&:C]m�i�+�d�?�{�|��AʪK�Y��&@�P���"�mB���]���{K��W�s�kA�qY?�
G0�<�v���%-��M-��e���#�^���'8���n6��.��te-��,n����� ��X,
w�ƽ���.#�(��n���
���)9|L#:����ԆFcl�4��"��(*v��� ���zs;�a8Kkm����(�²	F �-"�嘘>��2�P���B�K��-X�@�N�8���m�ێ��n,�9#X%5:���y�� %�4x���_?f���h=NA/ϝ:�g|V�8nF,,�`:V
@4/������͙�K�tL����L�JF�2�*��cN�y0�	���;b鈐J��!9ձ�M�6���S@9�r�f��MT��*4"�����P�ڛ)�h���Ù,sa��/�(}r�zj�����.~6Z9s�����6b�	VZiZ�2r%���NO��Mn����f:��p�n������+��j�qA7a"M��\3d��%�� ��x�3s5v7c������yM.qIYiC�3p��Nrx5Y��D8��{���I1����ų������(V��1��L�d�.�<pg�|��;�hž�D|��+�˿�g���6�0� ���^���lp�����ʎqV#r��[>L��J��вM­ȵ�]+����?�u��7h��'���IY��:Ⱦ�u�X�47j��.���0Lc�y!Rz��76:��3#xgO��i�Q�2�\�>��ߌ�������5����?
(�?����J�ʁ�e V�dlx$�
���	o���`l�����&o�W���et�g�NoQ?-�
鰤9	��}��������L?|d�?&��0�M�/�	z*�q6�yﭸ1��b>�J[@��;Xz�uͦ��QRڏ��v��*\%��h8��u]vh�nƢ��@7F���QH��M �Q���KJU��t|j(Ν���6�� u3�}1�E�7��ɏ2���;��3�M޳<��13.���x�ؑ#6(G�L[���&.k���\|����C+�@Qf�����j��q��L�[�s$�L��j}���u'����hs~�hu�^Ǖnw�c�:���x���ɇ���O=%�`ma6�LO���Z|�շ��HN%Z.�L��E�K`�w�R���o�$Tvݙ@>֦;�a����N�HW;���@����3ɳ�N��G������>�IA�3��ո~g!^{��EP	�1U:G\�>e�!6Y�.������D!E?�E@v�Ough�
��ʹ9��{�KJ�ҏE���^,:��X_�����r2K���������18h���<��~����v���{�F\�v%�_�5itx]���XZ]J�h&+����e ��Z��Z1\Ū��M*8�C����d}���0��`u�k����\�5��@1���h�e
�C�6>��{����cq�ر8u�H�9> ǐ�^�&��wvm��|b�љ���Ό�%�d�P���{�,�#�i����3�I����,��v�Yetȶ�"@(��m_*9
 �a�M[�����(��1�׫�ć���<�x������ѯ %��ԑ) f<Ƈ J@l+\sx��~t|,L���$ ��*8d�G١<搘y*�R�d2��&�qD�
������D���f���?�X����s�]��Ξ���`���V��6���}�M���^|&NL�f:��* �'����g������Ǳ������������=�_8�?|1�z⩘�9�ٺ�s� =�*�ĸv(;���m*c�J�D���@��8l���@��E�F��g;SC��ZKVe"b�4*6r 3���.�X�L���W��9@�& �E���'��r�K�\�E|/�صH�,�� �1�1���O��y
�8�%��uKr!$s�'�k���J��>t�y��N+*�.�F(�E��a�sm�ñՀ	��P������C��q�L8B�P}�6[0���R�&��N��o�����{��Ī�r����;&q�#O>���)r>�s��(w���p��ˢ��D�E�b���Ww������3q����>��`�s�~ܺ;Woޏ��t>~dx f�F���qމ�Z�Pu7t �Q4ɝ�с��gT�F�h8p��㕯Ӫ�A���HzJ�}i��U���鸊�Q@Ϲ�㽁���r<���q|��|p�����p
��6%����Č&���(�Q�c&�W1:ڠ�'����=mC���ʉ@������%s�����`�{W�g?�� ȳq���iX�G���cX�Rܿ{�6��.�O�����Ź㓸���I~Ȟ1���J�������'�G��ի �t��'4�16���V+��S>\������7������T
�B�i���﹡�}���=A����Q�J�<�O�;S�Myi�"������14wmu9A$�s����̘��2e	�"���X��^�Ɩ�/�o��z,�DZ� "-�⊜*������J_Ԏ�`Yv� �v�=6N�����#A$c�U���^z��x��`�1;�J��B���IOg���S���s�a�ǳO<�<�hL@��ܺJݷ�Uҝ�3��I�S#�#{�������OĳO]���\��X����	8��C�:Nv`M:3dw�矨̶_���M�����0�|�NL���L�{X�2���o^J���j'�7�9Qld���p���`�������[XQ�-��}N�%�H����B�)�9<�#D.�/��`���g&��5`8|OA�X���M��Ґ�+���	�#����Q6G�J�;16VE�vI͂aVk�1��ǅsI��Qw5~\�2
�7D���� [���6��8��V0B�=XT�W3&  �H 3���z��I@�0����� P���z'�#q��#��۫7��jcK�O���z��eڍw/�����ȣN���̧�♣iT^������>����p��˯��帳،�'��4h��nl G��)#�9�����߾�}��w�{��$�8�1�Iu�k����*.���c^3B7�����PqQ^�=�W2���{�c�a. �D~P~Q�]ړ�[����س����@0
��S��uΌ�QT����K�9t׆�LDJ���p.�T/��������?�M�ĭ�72硧T��=9��������������OǩcǱ�K����1O��d%��_�X�����x��s��܃c񡧞��(�Vs5.]~7JX5��ȵ`#�&���'���S��K+�{=|�l�?wګC?g�64D���h��S���|��h�0���fߪt�[�N4e<.��Dj��jck �AÜ���O�+����7ގ��tP�M�h���P�8Ng�[�^���u��XL/����뛓� F=��U�i[��	 ]7�=�_�/<M�B�e�������l^s$��Z�9f��6���[x��L����qlfy��5\3\s�2�Z5�C�C�q�|t�n� lld������:Sz|h0�������!��i���#�$�q�]�Ř���q�6F�C�@�2�r��D|������WnƟ�k�ǟ�b\�v/k#q��C��^�o�w#����T<�-Q�Adn>nݟ���x�ѳ�ɏ>�,.�:�5T��z.�N��������o�g��͸zw60�qY]��GT\�=�v�Ш;ɘ�z���}��;6`�� r�q-'g�;������s��n�>2�^�����y��Ψ�)�^ӏ�.n����G8|&��?N0����v��*,�̝"r��g�0��VT o���ϯ-�{�G��g��V���#�c��#����͟��E�6X5g޺0�Xm����Z-�@���'�P����\'�g ���
K7o�s-~��������\ܾ�G���7>>���1�u��ɞ6�k|��_���ca��[W��'���׮ߋӧ����-~��>FI]���ۼ��~� ���6J��e[��V*��Z&��|����rn���E�H�㫀����3P�������)t̈��;;�i����R �u��h��-7Z��>�g>��s�L��G��U��g��߽� F�k��y��F��&��? �$�� �e>5=/=�x�@��Y�y��,�9{ f�`s��(U�F}�L��#���>zP9C��b|�L=�H�8�p�={��8g�y��x���c�D|�S?=t1����f��Run׎սѥ���<i�'��?�T
��_'���{��=_�����_�/�~#Z�X���U͌79�,ȕ� ��k0���O"�������ѿ�(`��#۴���z�6q�jcq����Υ*�b�^z�Q�J5]�	P���\���z�5�RY��;��̵pr&1��9�?Aķ�*lá�B���b�����C<^W$g���j�wX��z�)�˵Y���vː����`�̅suq��sٻ�ͭ8u�d��'?��ήB��`f�תQ��ǭ[w�k_���~u?��'��x&��O�x���޸q7��?���g����W���/�英L���Ŀ���]�jO%���?'��pb:�ݹ��?���~�_����E�ΟÍ8v�l��O�D��D듛q�{Xm�b��k ��#Pev�9M�Ý�c��+K��n!U7'�b�l�at':)��E�@6U!tR���Ey���G�ǩg�W�dnS���F��aS{Qca��.���%%��i�t=���P��J� F�ʑɋ�,����|-�� Ŀ�H�z=H�w�4n�s�<���5mG�:g�]�z},�x�J������������Ư���g��V����x��r\����5b��lף�_��� l��{U�Y��fܚۈ��V����LUXk����)<�ј㠅eg�����z��*̣��ɣS��s�~��/� ���x�����������4����L�}9 ���Z�uX��Ï�ax�Nԣ���Y�����ڛ�p-�J��д����yl���q�u�đ8���7͢��F����g��>-4�;w�q�"��U:6�/Fn
��9M��g�,]Rd\p�Y!�,�{AA�r���E3�v&��|Χ(�p���s��P�b�XC�S��sB�ߡX>I�!4(C����isG/��b���ڕ��s�)ȵj����=�a�C���N��!��X���3��NF?wu~9����2
����B�:6�O�w��_}=^�N����T�oݍ�o����P�wL��C�c��cG*���y4�㍘�;��c�:�����/~%޹<7��Sw�l���2���̥)���K=3ӗ��N2����H���R����+�7`Ymn�6�͵ʃ�x�����ތ�R+�xh*~�'(�~�B��<����#|r�Z��*���}ҡoҝ��A]��w�>�q���#
�.���}��t����OT��XX�	r����ۄ���eKٗ;���ЭMZ퍳����#�Q�miwzc��p���j��h4�ca}/޾����X�������?�_���������4~�O_�_��/���7�����o~��������?�_�������[�[�~9>�����ݍX��k���vo3�������Wb v�y����:J>��*]&��І�-���ވ��z��ˍ��M��NЅ�8`1܏�.\�'NN�c����qm���_�	E����(L����io7bߡH��g��v�:������p^S�p8�n) ���K�]6ߋ�&�]@}N=�=n���fƮq3đ>D�1v��H����!��Ʃ�o*�:-~��NY�5GC����o[P 6��cs?|�+�͆�ڢ�Ί��<����yV����2�\���_�2Ie�i��JHA���S�C�p�N��"�����Td]4��|teʹ����_��#7(K_�������?�����鿌�|��j"��tT��7����J>|iʉQ۽��?���}����y-:���d(��c��TJ-��`�D���;A�Q�,��G9tX��-������ >�kz�k���z)����ߍ��~!��_����_�#��>�3���k�?�Q�ƛ#bNJ1R!ۤ����W s���˽��f��p�i\�!S�����$G7�������+��ut��Dx8���o|娙�}�;|���'��fao������4Te�,p5�a�nsk�������Z#޼t=^y��x��k��;��+��*l���z�4��� ,���z4Ј�.s�n�r�vn��)';*S��%ڵP�ӵ����m���G��r�T�c���vVi3��t2 m«S����l`�N��_��?��K���`����d����^�R����;����Ƙ�IjPE{
yL�<�|���T��}�]��w���.��x�xr�@�Խbt����_�����܊��"~�v�u^�6����Mk��yc�|e����l+h�ױ|���������?I���޹o��V�ş�?���Xu������>�:�*5~ �h7��CP��ǎ�����{qcv%�����ʜ�/���Ͻ��Pz� V�2�gN�P]��WnΦ�1��u)\�훸M��/�R�����І9l�9�j����b���P��C�辸��}��0�dҔ��Now`�� �h&�9�t��أ�⩧	��!T=f�6�v�Ŝ}R�y9��(o�����f��#��6h*�.�7�n��l�2L��[X��%�q�*�������Y|�\�c�vG�Eع�(����K�ߋ������?�_������#�aؼ^�Vk����r!in��P|��H厼��*����QN@��U��w���l�ay]Y��W��>Fu�Xkwc9�� �N9�O=2���He-&��qӶs�`����ێ��o���%0�v;{��\�ieq!: ��47���4����q�f7�Kׯ����֘kT.c�$��A6NO}{|U�����&����$�u�7�?</�����	"��"��̓��������l��
��n�1��zb~u(����$d.9��"�>�U�~��<i�1��.����Ij�t�*T�Dy������O�<���g봎��ߗi,�|�`1��Fk�@�=Ǚ���F��3'"6`9������m H�� �IL���8D]4� B�
�(�����e����!��m�*������ -|���W�af^:J��׿���F������_��_�e���݉��h<�쳴�I�R�,D��54� �˳{��w
Q���d<��G�����f�� VI60��82�ȍP��r�f@���[����HL��ђ���u�:��t��+�}�c�S�]�N+������\�/G�nʋ̯!�h�A	��Q%'�	�@#Ȥ[��mН��\%W�׭���(˩����K����M����?�����w����m��=T�vcc=���[0�F���as� �oҤ����\ĺ	��n�sj�T��oّ�x"���Y����a����Ņ��.h�ٟ	&�y7�8��x�����U��xM���n�������c�@AHjtx�oݼ�!;��EA�����Z��PM��G����皗C��mp���X�sU�,�c�?��;�K26�a;�Ð.p��{�aAo���<�C�h���Fl�-q�%|��"����|���QPAD�a'۸1>�̉��;�� �m�|^C�.?����*�p��LTW���T<��a�Z�:�񥯼�|�R|�k��_~'��_�۳�1�6EŒd�#0�Q
$��j���9�r!i���(q���(�{���ξ��'�J�,�A=ܺ���rP������192�V3N�<?�??��?�3�[�V<��c�̓�`t8R<��n����ήL+K>�O`0�F��>����}�������\-و��Y�q�� V� .��H5�٭��Ū_��;O��G�<?���w~���n4:-*/ǰ+~Pk�����n���Л�14F�\��{�gTw��3�țlf�|��y' :O�F����A��Y�ovk����m�ߊ3l��ދ	�7�tg���[A%(.)w�F�e?��/�����y])�����v>����L:*`8�W�����D���3��#���i|�I���\��	t���f���s�X�C���ZEq�g�j)��+�{䨌k&c�124�g'���>dIKe>���tn��g�W�	j*�ʨ"�]p�4s�h�X[ў��m�k� ?�Rg[����hб-ܰ��N�7b���bns+�/܏+�W��ͫ991�P>��&hS�v�Q��~�0���\�A9����\?CK�����]��z��.��$KH�Q���oYE5 �������h��� s;N�9���Ï>EQ\q��z��i���﷐-�n�,A�(,��M�5�I���W�sW	eQ����>]K�5~�p�T�9��굫����	�G ׵�.�������+w`�|��O>��� lG���܏���n|��ע�}5��#RV�:.N���<\q��O9va4�+�X]���#+B�t�̣Bk��w������S�B����:���Y�B4v���wv��>X�o��y���=�)�7|�+�v�_��{7�*(Y0��d���w`� �x���T&��󋱄b(8��&&L\��U��\�w��å��W���7��h���5�u6�.�Q}��!���p�a猌��f S��ۤI�}�S��@�̎,�nE	�0S +�N������n9�=�b��ԑz=�1�el�@2-��eI��VZ�y73c[m��n)�Ǝ`u� ����~�N�9�PL�K�|��Sd"��æ�;}�&]}N�(��P]],�r&���nLʅ����{%RV/){H:�ϝ���IUngLi�6��Q�����ݣإ\�k�ucJ�M�R&g���UH�Ñ	n���;_�����G}^���2�C$6�{�J��g�,n޻���ON�e�^k3�|�k�[����>����p���[q����Md�d@��W֛��ً7޽��<;_J��\\E�����h����D��ZL��p���Jw�����B2~��[t�����໩gn~V?]�Θ�����n�w�>t�;/!u�e�8�(^ٟ�S=���j��?ۡZ}8,_�fA\aJ�ҡy����5�|�%;�
IW�a+��5sĈb�"����cv�X�nbr"~�G$g��l����E��-�L�@17����s9�&T�̽F���*�W��S����r��JU�T�}ם�ڙ~�+�_���G��U����j���Q?�D�zI���b�n��g[��mP��E��٦�����\�Cr���q�O�S5|��6�P��J�ooFu� �۫Q�ߍѱj�������� �-���� �\���]a�4�c*
_׼�P*(6?[Ly�Po���oC�� �0�j�v���Tmz`	�=%�D��,Zsb �mڋ�*U�P���^�_��߉���O�g����uo9�|Y]]�-�ۢ��i�匁�����%���J9�χu�n֥�������|g?X9�gLgd�X�����W_{;�����p��K��*�`��q���	�л�`{�]���cU�p���S��;���Wbi���뒜f��G�RH�޽���l���^|:F+�g����B?Vb~a5��O��k���`5�7�o��2�av����X��lύc=�)�-�㢑�@�֕�.xxcq�S�����^/� ���L/��o�y�^'�k)����
�_����W�,A�>����x��o":}q���x���l��r��������G���ݸ7�pb���u���,*h� �`6���'_z*�{�|�?�_�i���;w&�Ǉc|z��8�s�k��G�|8^z�b��K5�c��D�����P����/�^X��w���i��#@�G'q��61�n���cX�݅���83S��ND?޼$0���E�Q��6���-���V�:Oph���+��N�F��G+�ί8st,>��Yvg���[-n�eY���&�e�
`h�����W���?�������������������?��XX^��c��	\��T��;.�P4�l$'f�u۪ێ߹�uE��*�u�5�Jh"c_u$6���ݍ�7`r��/��������!����?��?cS3q��Rܼ��)�ꡭK.m��q?��5����o�W_}��y��.`�����6.yp�~�'~"�����{�g���$�|�	��~�ѧ?��q�����D�`�����o������d�����%�luS�Ԡ�g�t��6�=�ߜ���D�8?/VX�H���v��gK�pO�x��~��|�oH]V��*�Y����Yq���ٸ{�COk�Ӌ��K�k���J&K�� �A�߻|#��3����fL�Lǅ�G�N�`%:k0����KO�?��+~�~:'Fᗠ<��G)����³O�~�	�tbk-~�g�?���~�����h-zJ�K�Ѻ��
�>��C���v��\l�z���]|h���$@2����U��S?��x�ɣ��R��G/����O�c�OGgc/�����{�n�[s?;�Ͷ�]س�m�L\b�� �`�C;���a@I�=���l������3����(^x�{<�+z&����-���Z3���ߎ?�ʫq��b�6t`m#���7������O�'�GÕ�\����R�8#?���[�.`|�=�أ?� �}O�Ĩ�R�^_-��F�ko܊����q��B�L������矉��uw5~�������`#���qi=޼4��+�ڛû�ݵ�������X��E{��ݥX�7:�	���ᱩx�C�ą� ���[���?��_��14������p+��>����+�<���ō��`��W�L�3O�[9������q��/�y�	xn>�im�������x��bzƲ����6iH�XFD޿ ��3�7���x�ze�X����D�(E��o�ߑT�H�Pp3W3T��U��ۛ�q����?�����u���~��x��Kф��}�<�;:���|>����5kX��W/���;�x�T��G_|6�w��ӱ҂�� *��x���8q�(A`�܊��5܆f�p����_�?��v#���k)$�W"d�nw�L�o����5�*?{�ن�x���=�:�r�����8L8E]��ƳSϟ?O<�x|�������)(�~|�������֕;J�ґK�~�JN�G �e�#��"t˔o�u��C��ч/����F�������||O�y/^�
�ɏ���\��?��~�r
of���b��G?��8v|2*��x��͸zo1\NR�2�J�r�r�K�J�=�.�M��������m�3��Ơ67�6���n�8��?n�[����/Ɵ|���e�E�pnל�_^��޻���9��t=bܒ�y@��+���S1n/��s1+ym�k�.E��x�r�����/�R�18��_��N�P攧��Q����}������;�K��=>S�tm��a����\P/�Ĺ�����@�|&�n��#Ͼv��- ��FͰ!n�_��޾�����#)q�R��ٝ��`yD:�Ss�Zs.�M��?��\�ǧ�	 .n\�� "�����/b�����;����ø�UD�4��9p̿�c#à��qdf<���t�r#:;?����G��%��^�~~��_�6��򮮯䤩#3'�̉�Q��ɤ(�X��_��x�ч����W_�?��+�e�6��� �uSH��\4�m�+{Hl*_���1yl!0�e�{[�f>�V�326S�3|�#C�œQ�������E����\�{}.W�rH��H��} �\W �A�te�]aJ���,
���o���WQ���Ÿs�n,��2�M@,녠�܀5�J�?N�w�J񅯼N_5�'�벸�y� l����� �a&K(���΢�.�5��%�pۭ(�w�9���X(`��x��\�^��"9�nvv1._�������x+>��W��wn��*�0��yQ�ty�s>Wy׽Q/G��t�֝x��u��R����Nܝ�� �����~�����׾_B�6��}XvǩUyd�[�܋:[Q����;7��؜sb�i/e�����n�ra�\+W�3��>9wtcy,W��ם�X�;����ez	" }N!5s�ٍ�g�㛀�.����_$��P$�l"|D�洅��2�]��� �0�el���*�W�����>�4_8�CC��O6>���b�)�M~����ň���jԆ�����Fw�̙3q���x�'�矍�@5�]�����(n�_�����Ų���ӏ��g��ٙZ\86�}��8�xv���w���ߊ��-�5q0GQv���@*���g�v�v���E!�E�����  ؅��k�~>�dnq=�ͮ����.l���{�M|�?@��_�;�-����"�����H��҅�B)�
���B�{Z+�d�e���{f�v��ós�0��XX���3�Rs�\���iz�������yo%�@a���.+r���f�r�Y�կ|�ոvo.�C|Px�Q�,��郪�Ke��[�.�ZPV����2&��(\o�k���&�h�Ǭ�_�u;�ߛ�Ytc[š��o�WE�\�V��Q��R�|ֱ	��%+�W6�	�B]D]�T�ي��q{~=V�v��+Ĺ-����n�ȾK:wm�z��vC։7���6���߾	B9�'#�q� A�~���pz�lZ&����x��86Y�Ɲ��>~�ؼ�e��G��9�$�}w��k��~�Ã0c8�$�  ���_������Za��sV�6,gk�A�=���˃�����9Ewtbp��p%�����j��s�\L�a�K������t6�*#�f��j稃��o߾N#�Ǚ�gbt|*F�&�s'�w5�\���k����Q�I��w��r:=X�'�WiS}x$��:���f�W���{w�c`����tn�)��i�+�?��Fr{��d����m�����r`%���a�p�޽|#�|�r���{��7ޤ,��}�oj� S]3���hm�u9J$s�2�����%�)���i���_=����E_�O�|�����w�ݑ��s�g\�?ԥ����Ҭ�
�.>%Hn�7�Z���,�-a������r-� W�p�]��lv��D(����ܻ��/ D )�d�_�֦m|��;����&ѹL:P�s�|��yE�0��	}��k���G:"�6{zf5�qq��*,34�F���d�d��KE ��.�n(sU=����D����ߧ����_������D������8�75Gȣ'Ο���>ӣ��\ ��F�v�?_�$��%:���;KkX���kW����۽�v����>Zw`3�Vd�bZY���Z�,-���\�*�=6>���X��M@��N��(T:>84B�}����H-���0�w���ZY���F�IN?���q���h#��O�&½*�����\�b�։���ȇ�ϧ�T�!�|��߈��z�;a�N Lp3�����Ο�I\!����ې�x�z�f�|��r�avn7�Lkb�|�-;1��;��C ��yq^��9-��>��Go�qM�3Bπ6��3s{��x����g�qZ,������+_�s�?�͎>,��l�����HS.���T|�����}�#RQ���lZ^���y�{X��qE�s��^�oŽ�6*^�3�\d���rh��&�3����������t#}ԫ�z�J���̟ ]\˝�,�)����d�uǊ~ d��.^5�ͺzi���E�{�m��f�A�k��c��<�H3|-�]U��q�����la�p9�h�_����o�ĳqlh;\�h|b4S6|����n� "$D\�t5��^}�����?�3���e�ي��vl$�d�3��F g�®��y�=�T�P�� �* r_}� ��W�F�~��h�%٣*���b8C�1��m--氩A`��V�FW��c��Q��.T��(dX7T�BP��p�wh��M��q|���s�C-+B�u������\;Ո�k���7�L8r� @��͠�.�m���
��έ��y��1<��y�K({��dff
������V�[��^�
��(����O8��l�G2��y���o`d#ny?˓��h���-��8
�Y��o�=�������[ewdJ6�cT�D��|��x��,i����u�o9��������<����:�j��D�sC���"��?�K]0j��aG�'�&p���]�7��;�y:�K�'O�Jc�i���v�kR�"�tE��6��OEa�M6�/�Y��&?|�/����8���*���*���xu�2:�k����.\�td"��9�� ��v�tSdN�(��phu�P �V\5l�kI�J��s0(����?X&�ц��0'P^��	"���n�|�m|�^����G!�����������)T���9*�/^����{|�������ſ�n}�-�ѽ�w�i�nY�"/���^����[v_�/˞�غ�@�O��XhfB_���q���ׇ��o��o��u�ã�[~�֯r�X��ݻ��<�[E�����{�;w����z'e�~�C�vȵ:�\�^ݘH��pK�:)�����n�v-t���m�~���p�_Q�b/��8��G�=y�${~X�֪tU��i1��\��bw	,�,4@��0>���7��$hF#@��A0`i��vq���i-�K��J�*��|��/���z��_z�s���p��nRH�Hp���2�����?T�!.�J�L\���y��wC����8ݱ�9L#��A$�����[G������4D�q"r��e��,4Q�H�'��V>�� ���j$Xt���0�	���
���׺W�(�s)\+Y\�p����#�u���KiF�O��k�!>��A�>�E�>̷��y�����ޕ�'^�/���,/y=�V^O���Wqq�/��8-�(�+��J��#͛���D�W���L�����?)T~�y�����������`�:!��J�l�5ѵ@���T(!�o�F�߉�z��Į �#7rC�u���B�oK�]��VG-�c��L�]�A���Y������!坃�9��2�,<�0gP��#�n%�]Y(N��Xt!\]�����9�74���q��S�΂��ς������+��3���̌K�O���	������S���{ �*`�K^�����
�u����������\ �*`�?w ����?�+W�c�����k[k�*\�~�j�(C/Cސ�9��P��8��
":�uH ���/��T�	�Q֕k.�/ĭ�W%�J�R��<\JCvB;��D/<�!,8�["�����N#�B�=���[Q��O��gK�RhG�-��2�麒|��=���2F �wąA~��t��1��@͇�ĔH�j� =�����s���`��X��4�nєd�+�?���"��wuU�UՊ��&����j��	��� F08&L�cـ܇�ft5�A�	�i�3����]f���y�1xůC���8�YJ�$|,T�ŀ�r�@v['�A���u��p������5�_����T
��}�g,jpq�%c!��V�?'��O��'0�ȠN��S��t�x�?�8ݍ�HL�aL�dSX�����e�M�� #7z?\�
���	j�2�7*��f
���^�2����/[��E_0�&0Q�\6�&:˧Z��*�ʠ@G��������p���]�R�%C<x�0c*���g=�V����f �s�?��w5{��s�r�JN�!^1�5�D,Kd2�G��e���"� �Q�σ�i����^��\i�@ q8CA����Sʧ��i �0��N9���׆�m�����/!�E�&T>��JO�
�Ao-��|��m��(�^�I������)�
E�SV�g�$�ƱGu�֖�Y�je_�{]�D�D�����,�c!n�U����pV2X2�vBU����O�!���;���u ��G�a����']��b\�i^pEq��ګE��j�9��e�ED�8�唝e�B���|g���,?o�9G�Ct�������\��k�O�@ʆA��7�� �>E[݈ �p�QBQ.q��<,�8t��G�	;�����iy�.��}o���� �q�H��ϼ�or*{�Y0��J���,2���GXʖ�����ԅ�
�<�o�&�v��.\F ��K�/-�.�|T�0�N��W�^�[X��38�R��*ҷ~�5'�����Y.�`	x.��q�ǭ�	��z��؀��+N�f�}sG�8��ߛ2�N�p��m�ϯt�@D�B�Hn�3^�w궻��3z�"���Y���$񛛙iss�T���+��ڮ^{1�c�Q���nXs5���[��+�OZ#�'��:X���v���J��� �d����_�2qaк���'�d��2eQ�F��o+��_�3�yw���+��lH��㟫������zj[��PGgA�c*��jڽ��]��湎W��g92�0Fa�(�`�_� V�g\�̟�*k�w�Z�x�A��� ]N?���p&iJC��ǁXg�N�SW�o�9qn��s@\/Q�2(d�3[3˽H����];�~��*N�<ץUSs��I� ��Zx�S�@mnڮv}���}��G��O>�+���Z#jR������vELP��S}O&?E��G���W��u0ݤ6&9���
�oy��Y`8�<*́�A���������F�����4�_�Q�ܟ��Ī�jX�Z\_�_��9�����������\��U\R�q�VM�v%b>��b���3Ne�M�յ�)��I@\��.���].�u!�g���(/�/D�-��JD�2����sz$�]�k^�]w�Fy�L#��B ���5TK���ju�}t�[Fq�&�D���Q���O������"�����rn�;-5�5�T�:<�x��>BT2;��2U���#(&/���`��,�FB؟��?a��,>g�xa��{��{7�ք83^`��4N��� mO���E�K����ûZ�/��<��,�w	g���k�<}��7;��=��%����^#����Ʊ@����zW���<�|z�u?\G�O��8�(N������}�Qn�t��n2r�DH�G���S���Vrwfz�m'N�5��<�GJZ��Z�k�q=�XmH��� ��RY�=�"��E��g��ƳP���_�+��}��meq
A@��� \}�d�|�:��,+�����3	+���_�ge�I�� ���B���0*�:i��#Z~O@��ψ#t<N��M�*_)�L����UX�JsT*��M}֟�@)��C�5��Џtͦ��z��s]�sB&N]O�w�]h����^:��K
:q~�K�s��s�.U=�����G�ƈ��Xg]�X�>N��{N���d�N�Q\�Hp�ӱ�]T��j��IG����r����ޗ����`T�lھ���/�J�
�S�����,�����F\��E�l�� �$�!�d{c+�k|s�-�lڢP�:�_��#�= �c����u�jV���9�}urSw���k]�:<�U��0��P8t9����?�dŸ^�&�JzHbH�{�U�
�U����$��<�{Inp�~�3H�qG׼��.����e�}����H=�g��t��g���547D��C���(`��?DN�e��tӢ���$bʵ���ӝ��&<Bvp<j�I�S-�>��#H�\s��CA+�iWq<�����6Ԑ��B�~�QTJ9ԑx҅�l�|}��`s��_�2�j
{�JfThiU(�%�*��@��O���uE�`�*���p�W��0��p�{oN���\���D��*�)c�ipI.���z�*-�^�	��\E9���)���x�W�C�3���g��+�z�Q����`T9<�k(A��R�w�W����k�_��2�~C�eyu�)U^%�E��W]d�«�w���V?>ׄ�?��bww'�!�ep]�X�K�|
屿��fg4��}�~1%t	�#�AN-S�kV��n�R0��x���'I�e�0=�$"
�4���3<I���a�N���K~t�Cm\�N�6���!>�V~˙��1m�I�B{��v{:y���w�߅u�����c�O���{�A���Y[�9e���~"!��7���e�̛��+֗	^Uq��L� �XMG����2���sh����x@8�E�&��T�~q����|2�L:H3o�x������!yz��F�=�Vz@��M8%�^=��S��`����<�BhX��3��[�I�I�xc#[�Tv@��R�g䪿���}�X?��0M���O��\���s�x����]pׯ�����"�s���v�
���P�0�1
f�:&�)h<M���!���q�ߝ��Qj݊Wb������#[��r)C֩ؓL�3t�<g'�ɽ��tLtƱE��w~`wP���p�:��S�*��˼&o$���@���.�@�dP��w���U�G5eX���7��Yf����5�Z?�A��0�L<"�r�� CVZ�I�T~�g�5ʻ�X��q��(%��A�*���z���Q�
�iW��yr_�6�:���������'���kL��>�{h$� D��e��v�
V$,S��Y�w��Y�T��D���G�W���� �����# g�<���4.�m��o�=EΫ�]�[0il��t|i!t��C��.�� �֙FN!݂��ߍ�	�M⡀7�Z������-��,��:o�z���s�ҧ��7u��f�d�4�2P�2vh�;L�	w��t^v��9���@��Ø����~SW�z�r?��]P����{�+��+�.D'��P�L��f������瑰=gy���|��_�YmyR$+�+����gq�ςQNJ&輪]enaE��@ `��>���Es�G+������	�X�'��uȉZg@	�>�M�,�8_�{x��	�)���Sq�0cqQq�Np�#��v��s��TQ����x*��(��<Fzc~�#-pxƿ��s�RB6�Ǥ��/�?R�"�1��4�	��������I�n0�ʩ�g�~�	ϱ��upu��o@�0��i%"� �c�mQ#��_ϑ�W�n�O�jAS'/��2Нu=��gI^d?�>{#���z*� �\O�y��Tz�� sMkh�2�����"!F�AW��~�R��
��^%BC�٩ #��ut��U�&�!�^�~�l�d>�<�'�	?��� �K�\/�n!9���$�(~}���/\��ǔ��ƳP�=�,@\�Q�pM���U?�=@�M<��#����� �
$�FT�1��U;�`d�y���%&���L*�*<#�8�k4�;�ON����9��H��χ��%��NIU���%���K�"u�)�^@���+�S�]�����-�p:�|��{�LV�7�7���F8��'��I���z�Ġ�I'���d�(�
!�D*�� P� p�L�Hا4"��o*�R�ǟ�P��<�
ʏ�f�A��{U�����7��T��I��{��4��g�73=�f��#��{�<Tt H�	�* �I��Y��$�ݿ�CX�3��j�_h-�<׀&�>�n�ѓ*q��_���Ļ�9�G)��5x? �;�=����<tʺ�/A�~���nNM�آ\*�iE�]��f�����hM����
#?��^�z☗H�z���'��#^)+C��&��iy���ĉ%�_xA��:$��aO=׻j�z~��V*ߏ��*�/y'#�#<�֟א��/�TVd	H��	#wQ��8��~p-	���g��wb*Ϟ�Y,�HT����Y໳ ��YEw& }�~5��:�� ��Lx���t����������gp5��_��)�;�ޫ�r�4�Pv��\���z�9˔�=H.�p�ٚ�>���`,�B4�Q��� ��뿎KՌ�H��,�k2�#�'Y���8�]���N��L�Z2 ����@#�@M��3�BNr��`R��e<&���8�%��uڀ~��O�Wx�S��/�����|6����7-�G����g���J�x?�Y�[�� 5+�kY�{���a��])waY�J%�H*^����t��$?��u�>�<}���(�_���)�����z���{��x�B@g��T6N�LM+�Ј4N��.���U
��P��u_��8�}���a�+��Ky@O�Q&�gàp�:��3�_j5� �s-WU��򰒴D�"R�)����1�uPxu媼���Q":��������"ॕ�+sY����ׯ������g�E���P��cZ��ц�"��������U ��!�SR�L�x�k��+�0������-�yδd
F�_AO&�@��FZ�' ��(^�`���=��Bґ!��b~��kZ�:��� :��S�Lq\~��s��tPL�z���)`����@Zj��V�֏�
�4|ga�T�Lr�Hw�S�O�؁˱��C9�M@�q�UX�?��]�O�7׃�ݶ�t���ñ]��&�3I��H��7����a�4���D�ЕJIE���Sڃr�����;{m{�q�������{Ҵ\�s�2L��� ���=:�M�2#n��Gק�ZF���#��bqPtvNR�ԕ��W��}_�N�g�*u��_�b���K��)�u�4>���1�~S8]/^>�dQ���>���8���K�2�L���9�@��!�$67�z���#�JC�V	��0����M(���K��A�VXT]5��%��yY�
X���&�g�ưBrD?)�0��
,�J��A��Ѿ%�Bd��_�zW���\�79e�V%[yw��V�����9��S�1�ĩ<�U%#T�Z藼�;�cq�+3.,̑�
EE:��a�F�b�z�df�f�o���Cd?��R�ʵZ^�Vѣ�2� ��N�ք������d��b�ԅ@�����@�^�yO�#(\���2p���dl��e@�;��3�����g�w��ᡟ#Q锂�q\�����v�n��lo��Aq�9��:�nY}ozp�r?�.oY��Q���N����G�<);a�[�8����P��G[�`�a;>�h�3t&�~��:���-�1�4��g�-���i���(�����i�˝��VE�[���\�.�^����k,T\r��#�V�H��E��"d�����G���o�}����cze�� �%��ũ�/c�)IߥE'y��Vn� �W��2L�aZ�iŔ�9*^A��!kd�0,���@�.�0֎y���s�}3XN�bފ��<��	Li�P�^����8��p�c����e���ʉ"�*ZK�H\�u��z�� ��s�DƕW�w�x�{�Y����
8\q��40���q�`jb@	
���C�'<���>���>�u���yh�h񜰼?�=D�Q^�g�}?t��{Gmg+���7�4 d��3����v(�q�|��Hܯ��t�-�٠��?��~�u����hs�eaf60�:����.Jj�������6?�����8���v��I�����~��uB=��\OSy�|y�orYdhXy��I嚟�����I麡+�F�CG̈ބA,8�J���
�ᓹ�N;���FڗA˺ɻ ZIWD=��'�۲�: ƀ�\#h��¦ ��%�R�1� X*����_��
�����Vʩ�R�N*CA4M�.�]���T�M�l0^�-vY,�R�_�2�EVɇk)ˆ���M|�*��d<��#� ��3���]�~?A�����
r�V>
�FE�A�pT���*��G�P�hH�(\�@E�h#t��P���L���8�C��j@C��PG�(� V���c�Hp���j]^|��/������v�5�&��s.�"�)�f���u�tg�n���Rf�Ǆ��;dWczc��m�SN?�K9�:K�l���]�������pE�||�l?D 6���Q���oss;�ҥ���k��?��~�/�k�Qj[����v��C	Q6���=�Be]��ZΦ��������iv��*��w��\�a�� �[B5�XY8���}�C6��ڭ/o��?��M����?�����O�q�[�Y�W����6&Z�ʃ�	Q')�i����"C�a~�2Ǳ�nnf���V=�H"����旖��.��@���i�@~F�����z��1;m}]v���/qfWW�	�-��}	a� .6���������x����s���( n��IJ�!N�������t�;�]��_��Jj���&>T�冰"ZNQb*!��~90i'�r�N�H������K��M���4�Y����0�@���k�^��*�J׫cQ~��z0>��̧q�I-O\�|���q����������4@u���q%v7��o�����FҰյ�07g%���3&�x}��ٍ�uD��S
68�"�򬴳�%������j�r�r[=7�V�M�s��(ș������?��_�?��_��w��vp<��4۲��t�I7�d�B���4����+�ժ~�i9��.��-3�G��ʡ`]L6�^GƁ�����y�������_�m�/_�qa�T"�t
�pS�6ܼ~�}y�F;��oQ�����?k���r���������D	;��k�(�rlU�c�j��y
�'�N�O%b�/-/��啶��;�D�R)�Җ��$�C%�P&iQ!�,汙��ڴ_��݆Al{#�3b5oD��9�~eJU���ղ���]%\�ʰN�%\�_���Ȝ�"����/Qq��3�~�����L�7r��Sv�*a�K^�S�(<^e
�4�<&�p6��j��4�;���I^�02�(���f�k|P�߄�M���֕�e�g_7��ٺ1݌�௟�Z�5��@���������T�q�f{�"q�'��;�8׹����/$����.0*�E�>w�|���j����X��K����6�n�ִ��nT�D^0ߜ���Cxiy1��^�E�{qN@��y�~�O�O�Y{�5޾��	/O�	���������)4�΢H��#z}թD轵��Bǧ�ԃ��X;�9��i[�]�����d�;D�`I����������;W&�DꘐjH�OwQ"n����޼վ�y:6�b�����W���؎��o����V{7v��F��g`N��B�z���v㘻��>�1����(�!��"J�o�nc�J,5/S	G(=�C["�T��4��!��\X<P"KK�%����"�>�#F]5���",����^f�}E[[Ӫ��
G�	/���su��M��Ι�x�[��-Od���^z��0\��B��A��t nss#��p������O�BAt�_��\ �/-N��W��<[�qU�N��v��v�Tq2���Y+ 
���0�w��T���gf����r�͟��@���μ�d�u^)BK���u�2��%� �,����t��w���䱷[3�=�)�Z"F?y�-,�@�����ey<�"��*���5�BO˩�ө��p�0ݴU��S�xSmu�r�z2�67&�ͻ{�?��������hry B��/-���Rw��U�~�E��p��&�a��mX�[G�:�h���;�i���w���_������.^�:�,�tO��Í�z���g��w��\�>�n����?i�%�;��O",P	�(�����8�����WA{�r��O��J Rĳu�D��������$�@�4�t����<��x��_�I�;�[��-Z�ﱇ������L=���8V�"�Z2h���x@�X�'��k�B$�q�ì�������� ÛN���&��� l�( �!ģ��+�eJ�C�UxҶ3��T��7�׵sk��/%�Lnz�o��g+f���b�2�g���ؓ-ͻ��DYX��4��0���g�T)TZ
@:Y@5��4c�-c����������s	D�7O��i�KY��i��O���8��e�u^��8��S��:W�W��k^�kYZѨݽCyLW `��^�j|H3�(�I�e�-ҝX��+� ���/���mj�b�~k��_���U�㟽Oø�����Ґ U��9�<H?��]�.}���5��JĹ�|�qLl}�8�Ϟo�Ov�Df&��~�u,��k���s�����T��Ȩ㋦or�(��?�8J��o����_���̶ s��]�y����LPt;�u%2@ �$f�����f�B�fAp��Ŷ�����PO��{߾�~�G/����ky*-���N��ƽ���v�{�^�s�n������<*�E����ʇ�3�	ќ�=�v���l���
��W��Q�{���]�R�;�*,.�1��l-��蝶�L�0�
&�8�S�X��PK(C��@���v�m���Rz���ף��[����w*D5R��$��.UM�(
�^?�'�����a���4��v?��	.�'����=��Q�8�r�!��w��h��������y��[j��ni�h�=��(��_]�%^��t�x��{��w�p	�%P^u�z�2팿
�z���g���_,L�w���3+���v��v��W����������Q{���;,�O:T�4-�H�������s�q�����5���y�ʯ<:K��}��Wۿ�/���o]J��8jDû6B�1�T���?mwo�E�`/��������۟��6��Kd�D�@,u�<Cz"����/��P*�)B%r@w���#������J�R���k����h�W_�����G(�Kmu~�$B�C?tsұc~�d&s�Is�)��j�{C�T�	U �`<�vA�JQ:R+�0���ʴU�b�w��&��]�n��cŚ�a*����q⤒��b�ϴM�MY*�����iuFQ �Ш��I4�7����x/�=�b8h��i<��S�U+���G����*��/�;3]���ҟ~��u�Е��qW�uB؄��kǡw1G�C����"�xW���y��N���8�u��_��t�Q��R"յ�Қ�+�E��G����%�/�?���h�������7���>�<����3=;]ǖ�:>]�#�ݯ����yr�2JdbZ��D��gfv�mn��(�����K��3߾Z��4Ν[H�k���
npf&�,R�֖O�@4x�	g<�M��ȿ����R�/�
kv4cA�4%8���Ю�x��C7��v����j���bvݡRQ(Gӳ�;Fk}�I��6>颢Ͷ���������*%A�çtx�w������;�����{��b}91��@��<Z��?�G��(�G��O\66n���}��&��1������G[�o�oO L�[�������!x��W���=?��;��DM�<�����4Ai���S��Q�3�gQ�i-ո�u��+Ca�~p֭ﵠ�J���݉H���e�[�ƪ��*eh�h��`W�:��1�Lǟ.w��;��B�0���T*v��&����.U��|Y *)�JJ�y��"y�*� �� ���l9������tHq��x-�ܸv�(Gt��kg}
:qj��R��ݦ���I���_��m�W���3-�s,<p1�XR&\Z�x�W���e��Y��{��/�[���Ee�
=
�����bh|O|�8"��������r��������{�Yi!r*����0X	zJ-��E��u[X.����Օ�~_ו�&�Iu�Ri�jG�ғ4j�DA-�������VH�(f0��2hr���>�� 
	�f�"h����y)�-}�OŔp*�uz~~�s �,^5�`�Iâ[ �2V���>c����r��Z�d8���ZK?�<��n�]9��Ͻ�.�'�g]���O��-u[�"�|Oc�X]��b5��0���*����S��!Bg%�C#6��b�]��:�^H�\A�t������g9u�'m�&'�c��A�E��һ�=��xXo��8kM:���믵���z��~�հ�f�<�n
޵+#Ϥ���oH�w���t��6�������?iQt�J�g�_c[4t;msc#�|�@�*��GN�8:���l0bW !�	��G�{����3=�M�3��
�� ,��-.-��;7ۓ�u��}�RD�jOE�;�BB��ú��X����X��=�4���)B��JLL*ի����5q���f뢫yǁR��c��쮼�Ep
��N�vL3�)CX�86�x7N��0E���E�M߸��h�lYU�*)�t�����X�'¸f�p\'�/3�U}���~�?�HڀaN) ����z"a�!�
�,�.4Fޑ!eN��W��w։̫�(Wyap�N��#֫x)���*��U׺7N�T��Qy�����T�\�J7�ע�ຑ ��
�^�2��������C��ַ�������_��ە���>�D�9)��f��˴̽
�4��3�s�#��4\<H�(!��,5O�>��U��A�Ǐ������l���Kp�x�������(pO&fT
&/�$��h�-�a%�3h��`0ީ����kE����ݭv��,��66�2#�l%2��
�
bl���n$��坧W�Z�--�~�,[������;V�V���at���`�tU
��sx6n�tT&*��+a�Q.��1�`*�����;����
eb|�03�W%by��";�� <�P���d�]�y��
eT�5ʄ�-c)�^��D�(��<{Z ���xC:B��QL����`M%nr�_��g���'y����*�
��'����vu�FQP��Hw!��4+�.��;|S|)�]Y���>�П�
K�9�.�����eo�G� �E��JV��h��ϡ��3��6���|��������w����x����`u����$��x�QF6�)�׀?�S��z�?��③��|�Zu��u3�]���U?I3�qjHM[���*c芠��W���t% �	bUH<��Yh�I�R"�G
)@�`|eb�bøNa�>�-6ׄG[�B�Y�a��Q�-��􁦿;.tC�˔rf,;3�V%�=���a�78� �K����}�_��]��k��T�u�Mi��=$�5sW�C ��L��qD�&�,��U8|Z�
�����FA� �/K���
s캙�J�s	RA��Na{��-!:	_W���å0�[��J9Tz6v�6.��g��Q�g�z�0BxƆ��>���W��Hy�3񋟊�۴�=c�ޟeʠ3W����V�vl��Cb�.(%����G��Q����\U �%�WȀᣨq��
�i:i��Ѐzl���B{��m��|���
7��8���O�I�B1��I(d��3�qE�%�=����
�4��eJ�H�ъ�\�G��ǘFH]�b���Z�8"W��#~=�|�����0����U.Ee�0�_X��������Q"9��3j/>DRHh�-@PX1��kw���P��^�R �)t��~Bu^Ki�3���0�Qc.T3�S����ů�p*\K��L��y�0��X������x��^���j�U:
]	���,�'X�a0Rх���$��x*��	�{�_��8I��-ǽ̘p�����_<�z��F|#$����?J�+��~�_��e��۰W�е�fP���s<wE���#z-�a�ݯ>ix����W�o�{.X2��]����L[r�pF�M�UNbe.��i��0Es9qݿ�9t��?AC�߫\��5e�]߄W>O�z<�oj���
�����=�]��
֯���8��	�;5xLO��J\�ϣ<����Ɩ�
��G�Ђ�����;~0?�|��&�%`!���{�3l���8Wm�t�?�%��+�A�w�PZjԅ�U�L���:��P����`��9O�y@�g�f��.��<�T� p��AYWf
�	#�?���s��Nϴ���i2���*Qh�G�&u.����k��!�U��+L��0��E"�ψ��O��ֺt
H�-�@�a��j<}_k>�Vi陟i�-�յ����� �>9��p�5��}�H��k�'�'2X�ҫ��Ğ�J�u�]����z��7����ơx����ʲ;�G.�Ѯ����y$b��g?P��T�у��2���VŅ���V����8�ý�~��ɓ'Y��7N��Z�:������G���}�c��]�WX�.�[�{�{��a�	r~�2T�d��N\��J��������,�
��T
$gp�T�C�?\y߯D(\�$�Wy�Rp�A�)�(��tx����(�7��Q	Sa}�B9i�ì���{C��7�I�X�+��R �l��MKIx���Z�цwe��N��pN�[�
����/7ҩ��x�7�g�U�U��I��y1��
W鈫?geWOE��̕��6����������]h���8��	^6���W�$�����_�-��U��<U��[Gңk�$�k1���x�]�4�7���d��[Cuf�+)8C�b^�!ϱ2 b�������$��ť��r���0�B��߆A�	g+��0�yf�8ς��Ʃ�S+C��x��ّQ:_���>��b��o|�)K���,�`��9��֬��)X��(;�k���i���pO��N&皙���Ѵ�|	�Q��B���Aò6�RD@� ��g�� ���EPϽ;T���Ug�~=�Y�� ��,"�Y{
z��k�B�eu��ck���5�/0=XX*��Q"��[	�
�[)��K���E��
��OrB�;	c!�w*V���tY��xM��8V��i�I~֗�-|�鹐A�3 �Q��%.q���G�/Vٴ�%���rO�*�PP���QRb�It�@���W	�]��Z�OjG��œL�k|�p9����8�1!�8�T7��{xpV���e��Q}�<�=��f'f�)��oC�Y%��ס�<�0�_
d�08it��V�KP䵐[��,**��	�J��P��*z��!��`�C���*H}(�u�� u6ԣ�+]�w�ԉ0�S�Y�����'���w�^O)�A�O�9��4�L��NAf�nCZ���c�8���a�C<l�ҕZd�wkU�����t��q ��`T�N�*w��r`��,�̵wi���w\����T��@,���N�z'�^{}Ԛ���qQ�{'���(�D���%�
at&T�����O��s�d�2�Ϧ�<���|ZQ�𢐐������-�
���鎠�UN���"�M[�����!��Y�	�i毁a���\��.�(D���S��V���"<I,��u��Zӎ'8e��)P�D�$���G��B��w���k���������Pɰ���&k�uT�C�_$�Ơ3�i*�'�� �i��3�C>��k�Q {�<��Q�����P!�:�z�6䩢���Ⱦ��;���t�#�7l�,9v����B����No��~Ҳ�HUWCeRy[/5v"]�<�����R�_uђ��
����w��4O�~��3�<x?��A̓$c.�k!�Fe;{���L"�#� ��# �aֺvC�H���t�:�h&x�AϜ�;�] M��rL!rq�~��/S��%�������n;�E��240�AE ¬w4ؐYlF���'h�p0��1= /,�ġ\$�~ *E߃��R��W�ش�j��w�A!Ȍ2�(x��ꀘ0�����ȼ>%~���K�VGQ�"����Ͳ��L&iY�vH�L��r�+��G'fF�|�t��+�� �K��42��Y���8����r�X��l�?���`�-?�!}r���P @��x��]�}�E���,�<x����(~)�R�}WI3� P>N�NPo^�v� -e/k���W	�S�Sʄ�)�W��-�p�9�gFE'���n�)�Mg�0���A��&G��@F����	�.R�n���3�,����xE��У�P(�u��'��^�,��l�O��I�	�?ɔQ���9�&���4�U|�!`v�Ǟzi]y�D���뉫��\<�A0�  ��IDAT�z��Ax�z��ޮ#���^��(�"�aX�4��8�Y�B4�+��5�!a��?�u�a�=�ng/Ў%d*�0�cM�ه<����jt�y.��6@!L��0rM�n>a��VK��s�A��?������Ŗ��_� (@׿�����laAǌ�,#Oڲ*(��T�n�J��A�Y�*]�%6��j�Ņ+���Q(
�¯>3o���-�ǽ~�B4I|��kyϒ�,����J8z�	G����"�%RB�0@q�� B{����=l�{��29I��e�!�̀�J��R�����`�H�4����<Tҧ�FH����Q9x�=�3cmzE0O��N͑~�܏�|ҥ+�2V�<��� ;#w`Ìr���>��)�]q��pߕ���Y���>J%b=l�\~/8�H�#�>9��G���c�ey<&7m��ds� e��'��I +D3NS-]*M3-��ɉ᙮��u��%�!���G]\1��ؽ{UIfr[��H"l
�Le%Q�ޢ��
�(��z�kcJXmè�3�q�}�ER����p�3E�����O�̣BO��ۅ���\֗�,�iDh�U-�0p�@7��\�|O@܉���3i����g�Yǜ�\�c��Mz���a�Ҹ�<P(i���� ���Z �7�5^oY�e�2�gq��ِ���<s��B��j��yN���<<�Y�E=�+��qU�ɇ8�S?�K�RxZ0�[�S�?��eLu`X�zY�2�b~�<�ޓ�Ȗ'�{yB9�1��'���Hv��*v	P]R�����WWe,�鎑_��
�gP�C�v�N�%RnXl�:�iB��a>8�J�C��@��x�30��x�ѣ���aL_@|$�(Ex�l����F1SZ �}x�J��>�s �݁(�:�>0R��ZB+��n�#�Vr�'-���h�G��<�/�W�`ℱ����+'�� �d�Q
A���C�� �3�-�xy���X�σ����b`��C ���W���g��JKZw�{����Х��n��r$��wY�H�Ǻ�w��
ݖ�3�0]���XάJ����_?���E>�Ye��������*L ^r?�fN<�8U��v�O�@�/a)��t�u�y��=��k�W�RϘ�9���v<D%c�S�ʝȩN�&�DO��)?�4�s=^P�>����;��<}^__��!�N;�S�
k	��d];!�>��֝6e5�#�<�e�MCY*L0�L��4,���וJFӛ����X��n*Hs����I�RH��E�"4��~��%�^���"�X\҅E��9�5���u �� ����ѥJ�B�)[�o�Q<@���מJbf�r!���G�x
S�����썲K�݃�Mu���a><|燦:d�����\ҭ #�-���Uͼ;r�~�����-�=vBs_��~ �)�N��p�v�`�m�n��(���N�'OYь2�����ݽ�(�44Q@�T�vyt��Ⱦ�U:�u�"I�1�X+`�1�+�еc��C��(�M�N0����=��޵��[�\}���;C�&��Щ�4�<+SE�WJL�TQ�%�A��չ����t��H�	+����#PIp5��i;��3�-��T"�W6}�&/[5�DQ<^g�h��FI��(e%C�
���jr5O��]�M���s ��A6��i�&))�pC�Ң�U��2���D��i���q>L'-qO?B^@'��a� �5��q�{�%3lC侄ف�<���l(aV��(�!��B���7B���
�=��$r�{�aT�tU*�u*���%���]@���;�e{q�RD���UE��9�ٺ/Y��'2;��ȍ2w�x�#� fuͳ���9V�FE��ӻ�'��˙�:��L[���D�^R�։9�`�ɍ���<��b%�3.i �۰�"�4C<��+�Pغ�*I��*���J?�	E�UƗe�]*~�p'�#�����x̉�~	�P�G��{��]	�����ѳ�GƊ �VI��<��[��}�����y�g��KA'�*nZN��W>�C	��s���3�7�H� �#�R�|O�ޒ���y��;��"������>t#|�J:�B7�ULyO8���(�܉Sp$���?�Iy�Pg�T��|�9+�����x�������^���ί�-,�'MA�.���k�E9��s\��[-t�a�C˃K=s��c��C��ĞɌ'u�7�i���K�]r����.B����7r���� R�Gf�B����O��B$n}���}��1��t�@5gf��0�_�;#�#pb����<�_a��d��(T���v��وY�~%@%8��ƌP.����;��q�-.ŴY�N�* x'#�W��e�l�d$��ۧES�����⵳��w���H��0� \�;pG0yu|��D�H~'�ٚ���y`�
�(����
y�=4 \��e�G�
���Z��8��&/��2�ܖ���h���2��a��ޅM��qRo����:�k�����ѧ8�؆�И��Qq�l@ʨ��p�@Z�<�]1��n��tZ�~�f��yꬺ��.r`#ϵd�fz��E��-x
����_�
�48�J���=zͬ��2B<\{F"�~�q-�$!rų�8���
[i�*Q/���V�r�A�t]��_ߍ�;��:ጊ*�3Y�Π�$��+�F�#Wq��L�t����W����+=�Ta7�ޢɰ��G���n�7<�UX�{���N^�������Y�X�2��^Ҭr��}��������?yJ�����<0L�I�Cy��a�ϐ�W �I�u�U�*۪�.p�+���V�<������RT(�4$�7�姰��T���{�4�D�p\��8$O���k-��� } ����L�4�Aν���Y?K���¢�jq���"�>Og���@�+R�'�C��c�I����D�s�%�ޙ���6]�H!dA�Hs@1Bm��Љ�P����=y>˹?Õ�!�]1��	�Re��̧��{l���Z
C52�;(�0�(.Bq��-t�)�s��a"����21o�
���7R <���Bsthii���n��σ���
/�V�?Nvٞ��.�\+M�w����e�����ps�E�@Ι5xԫ�:�|��^G@��
gGpy�����w���OSk��?q�,T��ڭ�(�2z$o�U๎~�����}�s���?~�<|Dz��utH�]n	���y)�g�N"�Uc�{��S��:��=�1�I�v���ῷhA�T�\и~�M��V�q]<�y�#��ă��h��T*K5����wa��t@G
��B�*�)eTׯix-����`P���V�w�閄8�2�-�~��Y�;++��/{��!�^�K&�L-��7����9@
�ƀ�W����z�`��
�y �����	#���+�a|��q�nA��,��y�@���$H���|J�z-(%U�]�jh�N
�k ��5�7�v���>���̊���*n�)��|����s�����E$y�x���:�OzV�g�H��ơk͗.�n���9R�U����<���Tx�D\�B�ǵ����f��2�/�
���
�L��Cl��^�@2���`��8Ï�4��C��ީ4��~�ϐ�Y`�*�@���op���B�<�ם�7���-���;18��z�&qb�U�&��aF�û�����h��ӽo�̂ᤡ+���&������L���	W[o�ߥFJ$���~&�KC<w�NO�5���Q~Cir7�y�e(���*O�ċ�������p��g{#~J���5�7�D3s{��T�%�35f�d#NC�^O�>�;�YAN+Y��r�{+S-�i���w��_gާ���Oz
lء���{C���Y ������L~p#!B
*�������)��|J�t�����̛Ç`�e� [�yԙ&��3�J��i�e��}6��k~�!|��R�����yz�F����Z(��:P��9��k�O�ax�Eaj:
�:їWf�r�Y�М���sP�G8����:<nQ8�?b�����h���z�Mū����Ӹ�	�G!b�q����������s���*���o|�.O�ѝ��/㹊2����]��8�P�S���/��}p�#� C���C�݌�;3x�� �6�{X��,"�T1IK5�hE�٫Pa��_�T 鞊�e�\U��Y�W�*�����u��4g]3S�D&�90�7�q��t�������Z̞�ީ��B����A����+�~=�}���:�|��"Qf\���>�Wp��G���{iP����#����V�W��Wo}Zᑲ!���1��̹[��[Ü(��W�PJ$�:H4q���A\���~��Ё�3o,//�G5"=Na6(P���-�m�@�v���%��0uG��#w��WQi��x�BV���S�EޓBҮC�D� ��$On�\ �y⌷]���O�=��!7��\��iQ<n�$�C:����e�vp��1�y?�Hؖo��O�l~[7P��(K�u���>�ȷEj������|��Į�$����l؃�u5%\�W\j+��� $w��;@���p��SLe���'`Z@��	�3��Q���R��{P�O}�P e���Ӄ�ƎaL`p�$��V�[w`�A�I���^��;��m����'���D�L����w2��8�1~4B�߇P���	�ak�7�Ѕ�������S�8=Cwk�3x�G�S�}�_.
\�`)��/�ڐU��W��X������=W��Ѥ�j��V�����Y�._ބ�)P�N�L�S�V�ew��:1^�^\��ggz��f�J� q(�V@	��`KX_����$��(�+�`�ʝ��\ْ�^@	����[)e*��<��֞l췭IǨ`*A�֕J5q�`N��K��������
G1�YM*(�IOM�����)o�%�p��������kGzZ&ǚT�ί�c��Ȼ�ú��g30E"-������$
&��-��w@&"�*�C�K���e���O �HN��5Jøy.<�-wR��
�A?�rL�������R[]Xms���n:����mU�
�"�O�7݊��3�~< �t����q^�S���4�>��<�g�1q��4�s..bt����}�n�Ϙd�k��d==�#�4\�ߥ�$�O:�"Q$ ���~�(^�z$�@x�x@�kv�J}V~嬇ݳ�|�އ���Q�`����ّ{�`$/�%��D87Z�e���,M��1�QF��B�E\.�*b�C9[3��?z��mnn�XE����;]@�O��HZYr�,�-���O�(̈́�Keek�M:ئ�B���\����������R��Ync܏M-��mƏT�ϵi��Y��&��~OQX��4�&�C�\���vJY��H"��` e>�8��X[��\f�=Bj��u�\��Т���ɩt� �3:�/  ��} [+Ck��w1��W��ʹ���-�>�gi�P*~��.�Z�`&�b���8�j�̶�6u�����|۝k��Smo���D0vf��b� ���f�z���.;4?܁d{��S��6�3��P(8芰�����*��!���\5����5\i�J�B�j:Yd����h֎��`S�>sSy~��*�!�Si��ޡ5�[T�9#��n�jdx �x�,@������vhT)�&��M9��Uخ82}
<"��T�V-2rg�:c)��*)qqEd��U��P�i���b����
����u�28D	 �(�C�qo��쎵�ö�'NS��~)o�M��)"0=���<0צ�f�ǯ�� �GkDS�� !��T� �	
ְ
ނDm�f�灆g�w`Dہ�I�0��$᪮t�����'(p?8�<ם��S�J]����ƒ�Bȡ=�T��z���?��Ctxn~l�i�}|��}�޾��^�콛�_\�h����O>��y�p�O~�e��郶}���B?��c@�\'�ɧ�~����Y_�0;3^�����PU���{�#�����bSK�@J���a���<�s��ưj,ǫ2��s����f�w�L[)��3�u�Ë��Ծ���6�gf��C|��DO��O��'�?|�W/���?����_�wmsj�H�--��R���nc�L�~����0Nw�"��כq���`OI��DB�OMі�;�6��a"�1������y����J{��ն�*q�Hd4����3o������
��i�cc���})O+9�"N=KO����ܻ�J���ɬ�fv���a�i��x4�CY�x����0�:�L���`�@�I��?���@�>��*���u��k!����&n��r�Ǆ;u�u�t�ⓞ��'�_s�O����u��xڀs,	�3:�ԕv�&��S
����k���X�+ ���������m�J��N���C����0I��<Қ�m�sk�ڹ�����<|N��C�=��ݣ��we��Cu�&A�֚�����Y��sua���'?&i�/��qiKX�y�U.'f�"���j[��LCr���|������n���Xl{vC����BJ.��+�=���nR6����7��N��/���\�����v�_����u�$��^{i�;q�(��͝��'����� p)������k[�����T��?�~{��5�r[;?�С	��R�����Qt)�y�P���pՄ���A�Di���R1M��S�J$F �����-D)����0��(h�̊-�_�}פ�䰢,-h�d�J�h0�zPڨR&�[ǩei���)���#8G��H�##�0y��gȳ���+�Lyx�z�3��ug�~����<�3d��ʰM�bmPfWf>u��S����w�b����[��݇���{(����:��r���S�ˑzS)�}X�42��ݝ�n빅�v�ܹv�ҥv��y�l^\�ni��M�E�w.z��Ӂkǉ��7ԇN�y�q_yMcD�d|bUnvr�-�V�\^~	��|��_|������>���Yh�[��{>_qQ���x���3�R"�q�mP"Q��|an%��6]�<H���V���������ʼ���o�=��hY,r$�C����v���mn�B���������۞�;��?�Y\�i��7�Ӯ��K���9
�I.#�Z�b��V���RP���5h*�xrnW��p�јj�L�+[�q���~b��v���0��mg{��n�{w���y���+����`��=��:y�;4����϶Z���E`	�Əg���c�Z"(��7]gj((�Jn��Dݤ�3�?�^��H��X����I�PL����}.E˳�5%��E�S�T�*��R�`j����M��`�]﬷/>���ö�"�¬>�y��!�M�r���p������2x���"Py/-/C������^|�v�kmem��,L�C?�Zû5�#ڽ����K� $���(G��K�6Z"������<_l������������'Q"�t���_��,WAN�ՙ���4�#%"_ˏ�|~V%�ж����v�;���o������&c�����wP�� �l���.���Dz�xa�n��s��?k�~|�զ5&����לו' �m5�^-�5�V�f�g[��])m�p����E*wa�j�\�
w��".�����>�2�=�~�5�P�%���sU~��Y�f�r��B�Bq���;�ݻ��}�����_~�����ѯ>j���u���������O6��}~�m��A��c�Ҫz�Y�@?j�o�m�o�mha}�y���	;v�x�8S�4�u����7�(�F�L�-?.�����g�;4�ۯ1��.445��E	+�	�K�<'��N��_�6�}����:�z
�oЕk(α�v���?��>��'�?{�}������	ݙ=��m[@�rbY�B���q�0g����+�@\-ϵ�%�/U���>�N�t��ОlP�Z:�|z�2+#�`1�JPH���'�>�B/�ӆʒ+_��8�']�3�����`jl�M��Q��v��V�����<�[56���}�� ��r�W���4])�Pe�l���<t��Ui���/_��~��/����q��+�����t�D4��ҵU~� ����3����S�}�v��yG��F���Ɍ��3�Q���c�7��b�Y���K�LMϴZD��8������-D��/R|�v�" ��_O�E�_��O;'��#�.�T<\��Ή�c���CS��{��2�a����n����w�@n|~#�b�	�&a��a\�"Oi�a�d�)�c��C�i�B/_��~��w�/�����,�<E��46���{�ލ����;m���佛��n�V)�:�!�3�Ty�ի����Yg0�t�u���	U�aX�]�(p
D�d@%g:��W�U6�Ahb��2�҆&X<3�u;1���J������?j�o�m�7�J�f�o��<�(�.
���<U�Ö ��H��ٳ_T$^�h3����>�ϲ�Z�:�A�؅����4�7��H��D�h�=�YL7u�c���4����r-����+���a �NLQ�I,ݙ�y��|�{�I����b�<U��q��/�R��:4�Ё|�D q���y�'�6��h���W^i?z�Z;7[J�O�\�z��H���ە��b2�V��c��g�~�~��m).�X"�*��]��g8�о9Q"�%B�"�[󝞙���s�;��.]ZA�̷�9�V� ?�+�*��D�]6gQy6-�aH�U-��^������	���h����}��v������}�>��G�Vٽ�w�.6�P&*�ASy6m彩��7�WwF_{�����V�7�������*��vn�|�t�r�r�j��v��O�G!�P6�?j�o?h���ý���'9��T4˾~f'Sf��O��V�Ik!H���#7���WC�S�=��?��n�o��n�e��k���$¥q�tv����B��Yl;�����{?}����~ܾ�싶M��)-�]@���ٲ2�ք�͠$i�?�e�!�џ|���\!i2�KO��g�4�ݽ]�G��Ȉ	�̶�������%�½-�L��"�mƳ��Y�{�Q�cX"t6�D&P"�n=j?���t/P���a, )}��,x=t�Ǟ�� .�3s	(M�(7x���o|����Z[�>H��<]�p!|+tH7JĄKM�;��O ���g�}Dw拶O�0�8�HP���T"3�0be�D4=�a���v���_E�XJ)�z�1�2Ȇ��"�r%
�<�>fi]���D���>=8����[o�}��4V
Dszg�2���G�����@�L��0,ĥٴ\.�������o������;�iX!n����oK+�,��_y�������+��/]�_<���}��>�h[OG�G�e�"��*�Y�J/X�A_[:�G�}wR�~�~�W�g�u��yx�/d=��.Jڪ����e4��W���98=M�:���Yj;�{���>i���I��?y�(݌�Y�wI�|T .�K���VYO�`AB��A��� ���vd�
<���w�QxUp�x���n����4Fn��t��:�?��G����20��;��X�!���Ћ�U"����?�ID����_�]i���ۃ{�4���[�:��~�����y J�i�}�K(��ç4�(��Kc��7�jo���%M7:����^5ʖ7�<&~↕��T#��ￎ���=���V(�`�T	x�vJq��L5~��}@X:���
CSڙ����A���o��O��/���Oڟ��?K����u,a�#Ta{�v\��NB�)��o�����?mE��/�l��[��^��?�[�7����=�;�e1>��0<P�����������ݿ������[���a�F=�"�Տ�����?����������6q@�h�ƟB��X+s�yS~XZv&zƝ凓�vM��>����O�}Ƭp YE���� 9�m@^v�j`��٩��֗�۟���ڟ��?m7>��v��]\^l���mKt=����tM0��i!x���S~�hn�M�Š�%;�I>7��fgy���4��~����?9���X,P��2=��nДr�K�f����t_�v��~�~������q�w�!t�2�� x�T�V.V�"��xWɞ.i4�ଊ��{}٭�|>\���xg��Pg;��l=*/�u�>!g��������Ǚ׉�
9]j\,���E����&S35&�%r�O�IؔM-���vgjl�>���x�xquԝ�[�  ;?ӱD_u�bF�2A�3cߓ�^-SF�0O:��<~�g?I�ž�K�gh5�I� O�<>���5�InԺ�H�o�KK��~��~�Gva^ �鶉ea�Jbm�ʪ]�{;{�ڵګ���A�O>����T�����v��������N%/.,F1�r�
�L*��->���c�S���-�x�'����G�ü���>坒ξ3
�zw&?�����>l7��m��ɻ<=�=j���i�ߡkw�x�"8��2�C�ǧ��^=��P_	�Mb��uR���3憲p],��]��7�1]$��Nk�{�׻eN����ݝv��}��T[]]�!^Ylg�J�53��� yC��D*��#PNi3]2�:�R:�h����'m� +�����I}�墜B���?�*�p�@Uf����v*�=��{�腵�4b�k/�N�����^]�n<ݟ����;����sb�p	�3A�1�A	pW�-��ˮ=[շ�K=$�*�
���s!iE�RY�]}q�B�y(I:��r@˩���Oڟ�ɟ��>��mo��Z����AL2%�t�̒�,�B��h<�	�����ggP�e��aQ�*�.��^��R��ñv�y�v��C�������l}J��Ő��k�ۋ���k����X[�	�g1�������G_��?���67�D��v|�*Wp�O=�aRiʜ8i^+L �@�b*�����!�ZZv0B�=e�A�Z~�3�Ӡ+u�ɼ����n˻�x�ݸ~�}�������?�wۿ��'�o����������{����՗_��2����z�}��ys���5�������R���s�Y��s9��Ox�;�N8��ߟ�ϵ9S�O~*u޳�=3��f����E���mqq>i���O>���9<��'�C�1�>���;��	��-�/�cP�Q�ȯ	�)k��:(:+�wZV_�L笚<q�!��y`����>q ����y�����/�lO6�N���/�g��Rb�ʦT-�Q {��Ks,�s�3�;��!-Y�ؿ�Sa��u�{�����|�1��8�j�9�e�%nҨk�"��
T��1	�2�x!����i�h�=���������q4�Lf�e�m�i�Z�����`G�M�Yuv�瀌���Zy�0ݬ��E�.��a�c*b���]�]ZV���~�ܰ�� Fֈ ���:�/���Q���Y�+�Y����Ý��~Ўv����K�zB@#�'�+3"�ٚ��5xC��� �'N�s�������)����l�m�UG�U<��?��Le��B�|0�|��}���m��ö2���z����?���|;<�ms��˯���z���;��V{�oa����sm�.�2�YB��秎P(��i��?�1F��S�ζ��.u���n|?M�ϡ���QP��Ų�s�3�n���Tz�� ��x�sЂz�Ӓ�n�@���FƬ��NNS/�/�Ti*?k�f�߱'�;���p�L���m�)y�Ws($Ä��]����:�i>��S�ʟVI�Mcb\�s\]����e����t���ow�ާ��"���hs����A�xR�:M�E �A4�S�]�(�u�t2�\�"@�	,{Wc*ҳ%T���/�)H�*�2�*��TBy (G��nONCɨDҪ���:3C�d�q�ޓ��?�y{�g��[�Q��>��$h��q�`��St� �@�)����h�e�[��*ە5Z@tyq�-�x�Vnmq�-��$��������v���f��;�;m��e܇&Ӷ���.B�#��&;�R�g�iq��������;F+����=��02f��2V�H�xZ��mk�>�
 �Aj��J�t�`GHoe[_в�f�[�G��a�i���r:F����x�m=�k_�w�m�y�.έ�w^z��r�6�Q���>������ЖW�ҥ�N{����_|�]:w��.� �mme�2XE)���gP��KS(��C=,Na~���t�p~���Q<�/T�9�{]��aA�E3CW�� k9��X��]T�vg�&��/��z��Nl ��Y��?�����?���r�>(%�	����yb�߽�H�)���8c�V�={ܧk
�ז	U�=	��΂ԏJ�,;�i��3�F5���e
�?y�vh��K<�иcN��^0O+�4J�ԘzƼ��V��i8M���K���9�D3�I��hơ�>8���K��;�n�xss����?k?��Oۓ��(MVs6#�b~�:���, `����0�c"y��{������W=.-/!+텗^j/a��;��E�iB���K ��L���Ҋ��5q6�.�R� ���^��~�nݺ�>���v��mc}��@�M�xu �M�"�PݥP���`h��DX(���28KX�Q(��
���#���"es��B���)ZT���w�h���z�������|�v~�|	֏M��c���ٕv�µ��+o�o��������O��V.�s��ڥ�/��+����+�깗ڵs/�ο�^�zm�\_��j���"]�W�{�]Z��p/�|i���ە��+W���Zf�V��Q*�44:�jQR�vW���N�q�q���m�>|���'���yfgT �3�Jٺ�<(5�V��[q/n�k�A!��v���DyE�T�L_����UO���{OXyv� �E��
� :�X�^#޻?�Df���~������O[a����o�훘7�$%q�uU~�7_X	ߨ����Ԓ&��J-��sK���B;~����}�������{�Q.L�|,�&�-f�k��biia�n�z��O��}��,*?�o��&eR��]�Q$*� �ݨ%Ca��mRA�׶Ol~�2��Z�����~��߲F]���h�nު��[-�3EZL�ḿ:�I( �ݼ�.���[���@��EB��	-Ž�����;w��AvD}3�rTi��Ho[�,K�ٕ�t*�2�/����\���B[��05A�&���i�h�h���f����n>hwo�G�Ϸ�}�����ª�BAȴ~fg���TB�Q�v3�.BW�bx]Z\m�+�`���4���UV�s a'��"�Ks���Z��z��[��bZ��8\��ʥ�P�k�kr�-�Eu<K��+K\S��f��BmcZ�ޫ�ugoT�66:��`/
Z��{n�B�X�*碩�C�R��ձ��v��#�V��$Ƹ{���S��#-�?�����2�\+�q�Uv6�����Z����..�#o7��ѝ��L/����"�Dt�ס�s���9�g���TB���h�Sf�
�'���/{�o�����u�n����O~�<��1�y&����J?zJKd�Hܨ5I��)��) ��D�8.��y����έ]Ȣ�+��k텫/��^}������9?B$���>\w f��n��vTz�!4� t��s6�Z�Z�MY�D�M����G���/o�_��W���o��������!m���s�	�G@���B_�s�и������+����k��8�K8�U*i�H�~�BaM" ��q�����f[�Yio��������Nf�2c�S����8�0�Ў���Y�Z��^}������oW�6fεs�/�k�款�f�.fk��!�ͶҖ�/��/�Ͻ־���׾��|��ۯ�V{�қ�)�<E��kIo�}�������پ�����/�B�u�-//��PYd�σ�lX�x�~�I����h_���}��'X[�(T5"�G�ɮGw����B�\���ATy���.P9Õp6����_yк�"�*��ޥy1N�SJ��5[*����:�'��А2l�H
���a�x�{]��h��; []^ż�j�����g�g�ѣ���OE��O�)o�ʣ��tU0��F����.�aV_iW.^k��k�d�iI�<�b��_x5-���(�T��Q���p�'-9��`f	>y��
���h��9ZX�Oⅅ������~?W�{ok����f������A�c�����s�^���3G0iW$����9�X?�P��� ��o=T+]��^��u��q��SY��� ve�R�]^{����[��<7�B�U�Ș��q�'�2�wS����voέ\���:V������7�;o�V{����^x��r��*�W����+��U���r��̝o���t��vn�R�8�i�w����b�!
�����F���������������;�|�����Y���յ��\KBe0�eJ/l�A�)���(�ں栵c#�Q$P��u%����O��NW� f�*N��R�|�+��M�u_uk٪>��W�����Ug�>�Ym�9����rŘts0������R�(���s��2�������s�P!����������Ca�ԭ�i�a����(-�����+�*�X�JXAq\X��.���.,_h�st?&���d�[��������k�n�}��ŵ+�_��f�͍�(i�jĸ_��B��(�;�շ��U��E��F~�(E�夰�C����/>��}��_����R"�}B��2��d�R"���U�@�0��#j�h2�a��d��_%$�����k��ޓ��G_�{w����9����|�\�S�
ˑ��m��D��`� �� oʱD�di%�Gb�8]��xu�|[�.ҍ�$劉�� r=�9&<邃a�ӝ�|�*u����w~��/`1���K��Z�z��v�����B�K�e._8su4����`��ϗB��\o��~�[i�8�)#�Zͮ��݈�=e.-m]^����ųa�~�:.J���B���Y�����I�3��vd,����і�ܫ� E��z�}K̺�AQ͸��t�����[�"4H��ü���Z�� ������Q�8F����6�l�_���v���J��:�P��t%R��|�����=�jnz��o�-����t�~�Ŷ�I�0��)M+u��9��&�h�^j���o�~�w�+/�Sz����=�[[t�-���%�V!]�,^�����ew�����\���H�w��+*3u�B��:�U|p�Vf~�w����ħ��҅�4R1�T�i���:
ァT�u m�����/�e|��q҃{���~������և��C�klqi�-�tp���#�v�G�ur�ܣ Uh�"4t���"~F�ޝ�睶���!�])��x�h�n�.�&�_�{����WVϵ|������=�T����k���q��O�o�oo��f�~V3�27��bZD��uu=
�k��Iχ���)ipN���|�;�;6/i�]~�NE��A)x?\%���f�V���<��?0\�E�>��aH{x��tU��l7�<J��|��Wfg� ���S�Q{���/�@�}�^��L�3U�2���P.$��?��U�:߅ ������qp�f{����B�:I.�)9�8�+��)�� !�1K%�2~��'���D�f��n&��Ck�qgZ�쥅"�p*s�zif����X��[hӘ�cK��ܥvm���֋�w^�n{���7_y��r� t��+�.���f� m�B���)T�����N��=豹�#y�6��*J
E2-�ͺ�߱�}�� fi��w��;w�_����43"��ʮ�G�e�8���e&Tk��V���|U�}���=�
��ݪ��]�n��O��'�s��k�n޼ݾ��e;�E,, �йr9@�n�=�	}�>4�sYT(�
JH��{w���(Е�]`����{�ݸ}�p��㍢����ŋ���mks<���ůڃ�����{���w��zb%���RW �6�%*r���rދ�]����>�Hk�����38x
�����u�v�eP�ŵ5�Xj�s���/r#��s�����5n?���)ǥ4:���C5 Vb5�楟=ǈ~~�unJ�]�,��g�g|��@)qD4�=���.ߩhR$ 5��/��F)��`����l��"���O&�0^�d�CK�knWS޻s�V��ّiv\��!��!P(YdќeX��Wq, @�L.�e����vq�r;�p�]]��^��r��v�+��v�dm�B[���A���G��?j_~y��?�j� H}�)���-�Z$hz�0x L�eKY�vv�֖��������K�m�������
L���F�������\�|�ƽ����PA&�t�J�:J����B7=�s灁��~x���~��.RW\I7�\?�������ݽ}�|iv���7ۯ>�U��聭V��e�_^"GS��1ek.�m�s��([Ƒ��~���ڹ�|t�����mcg�TN��p+�r��c=�������r�[�G��k��?o��K���[�n=��B�a���~׮f]���8����wm�\YFX�n�����Gw��{����e_�-8ȣ]BK|h^t�*@ګ�u*ץ%��cM
s��ͮ��I��Wr��k�qd"B%��iu,���j��K$��>�����j+��޽{Itrj�}������>�oB '���m���L9�'���z�|�T�� "���uo�칠"d�=�O���s��y�g���̠�g���ȗ���g"��R S��V3u{s'-���ť���-H�,�` сG�@��ѧ=�|�������K/����9Z�������tU\��ϝ�.Nr/��K�0�ۯ0�?�⋜I�ɧ��;�ց�=�~Ϋ�${���ǜ4�,���e����� 4�i��&ߣu(z�z���A��A-�y���١�W.a�L�B<��ꆪ��д��_Q:L]�-R9���nߣ�X ?m��jd����*H+vu�B�pAF!ƺ�خ��Y)�m��bZ�-��.�v��<���q����A)d��>�T�{��*i��<�C���d�ݺs;�nݼ�B\� >(�|��Vћ�K�=�N�6=���>٥��C>RvB_☖�[��]�!X@����K����+�#��ڰ:�=ݦP\��+���D{���ۧ��n�
qd��WB..�F7��~�7�K����#�Ư��f˧Q"����.��.ҝ�VI*�IC����P�p���R�d�-��[��O~�9�u���M�D�v����"e�,���'���a�v���q��b��#��2O�]ޫq�Ƽv�i�U�k�[l�)J3�p�M��4�۹���O>o?���b�nelĴ��
��vg԰�yq��z��9���vq�b{��o��^y�]�^��`������������Ћ��.]lK�+��/��>��=��o°�?IMI	��DP���T�[?MpOժ)_��]ho}�-x��lo��;���(��R�<v�ݥ�(�*���t��x~��m�&ҲK�b#�����x��:mB>�,��3yN��m�~�a������y�gr�[�]o�����%,����?uO]��@[\qr݌eS�h����v�����^J��\����B��:z�<�;��|~������~�I2���v���֬�TXA
�3c*;�,.��`���^u�kY<c-i)ՆUӳGVPv�
Η�LO��l��xk'������������v�b�'R}W�ϸ^����g:�3`�s[
Dzۋ�Q ���hQ^�~������ǅ\+�L��� �2b�h��h#3�1���� �8Cr=���� �5Ų�%A`^��i���*���ٳR�w2l�O���ce��i��G�X�۷ngQ�L���:`�n��L$�&�}m�@��(�k��my�M=E�I�Y���E0=KU��`E����c�8��hc�}r��v�	-$Vۍ;��#�1���G�:����r�\[�pAk�/A@|���	�h�����ڋ��i?�����]�N+m�V�v�Y�Pʗ�N5��\)�3R=7�F���O�������+):I.�Je�r�Y�@Pl��,�q�m��~��!�ڲ�S
�����{7ۭ�����St)�(�����,���7E���^U��>�2��U$׿��}���歛Z�ْ����xL��z׊�FQ,��7��φp��*#��
�����ᇝ���Iw�j���m�����\f�\���V��Iv�]�q�����a�>A��݁��9�|JAC����B��M��݉l�%]S���g`�/k�ɔ�(Pe�t����#
;;4�IG� �����#|2���ԭ@�R��*n�0^�����'lq#|5�P���t���l��P u9n��u��/%T0�C��]�g��a�V��B�\�+�"�%����8v���X$N1� ��jf��}�'V��$�`�]�r��l��nw��6?�y��O9�h55�UZ�K�E܆Nu������n���v�{br%0��w����a�7���w�[o|�]D-a�{p���Eic(�1ϸ�u���|����n�H��?�����F�iG���z�+^��g��#�P�<���i�5��ܠ���S�y��Eۧk�����>�˓֞0�J�Н����=.����'X*�y,I���C�ku���5����0Oܕ�ULp��~����(&h�^��A�s����[�"5F6M�H�#�Ώ��HWvzEr�̻<�^�B��vk�5�Z���j��a,Ǣu)o��CB���[�/�����Ա����`k����ɳ�X�ᔌ�ú��{���TZv�ѩh�P�g���MU �����ǐf�@�@zq��9Cȝ̲1Aw�m��1�q%�at��UJ�\浢a��MH�	��VQ���S1�d?���ǜcJ��ۂ����8�Y�p�^�s)�C�R���6�8�&�U���-�m�.��	fa���Z����ŗڋW^k疯���estle��-�ʣN�: �c�2G7h�V����ߢ�O���o~�H-���)]���������]���E�`�C{��N�����T{�ڷ�������Ko����6>s�pn���6���@�1I7���������;t7\��<* cGv'C��C]-
uCQk��	P��mD�"�Pda���`{�=���=~����?�(�g?���]\�CAh��i�^�{�V�e٧ޟ~0��/��oS��f�>�W�Q�t��i�w�����E���EY����v廋 Wp�9��R*�*�qx�-����n�����i~������/�Zr �A`����-X�H���G��)e匍{���?�џ4�l�h�\�����M����jzn�3>�1x'����?�&=�5U.�ǍG͢��B�]�2	�*CvIw�"qq�[YC��PwX(�.,0�!S��H��(5�ӇP���\30��u;z>n�"�0o�'��P��\�B!]�Bjx[��[bo�K�����_ZS��>�	�0�����pQ"(}RS��2�?�2hsmv|��n촻�ob��6�o{�������M�Q���m~�{qr>�0���v{��[m~� ���K�c�+(i���MZ�=�srv���~�����ū/��G1���
!<GJe�������WVϷ�+�������y����c��?����d��/���}�]��vn�R[ �U��6;E� ��$��0���D�/�f��<��U�aj�A���S��.Gw���b�j�x���F�P��lP, �t�M��
�yLD��Ŧ���B]^�����̿�����Xi[mvu��ا�F, ��.�o4(w�D���Hoo�	,��9���͂+yi�O��C��P�
l��͓�"ix5�|��������kI� �|�s�W;ԩ�c��SN?>�@�A=�f�y@ZN��H���̢�'rF*e&���cZ�G���/�ǭX@Yz �KT���#��o�",5����m������kH�+�$ʲ�˷䈲��:���=�Yq9~V��$U��4	�Z��Xrn$�
s�']k�pְ��\�%�8��9j�͌̉�i[��/�=5�Q ��e��_Υ,��U��9��c%WW���jկ�D�
HM+a�i����!覓Vӿ�`6ǩ9� �S(�y�#k���qy�%��}�/�i�=����o+E|�����3n���Z�]s����-���!:B�a�B�!� 8�����������OM��_y����^�zr���E��q	�L�8�i�:N$�nݺ�nߺS�(C�JV�i�F�.q�k[������`_�g[+K�Q�4@cO s���c���MAۇ^��>����w"�8���uCZ�7ӵ�&��ӌ��]g<W�x�R{����+��֮�x�]�z�]�v���[m�Km���v����*�l���tFH:ؕO9���8���%O�w�>�iC��5�~��߬�����Z^;I�7<��蚾3r6��ri�.?֙����4Ά�ג�vbK���{r�m~�� D�O�s�������U��#��������ӄ���@p^�Rq�l����/<9�*�����Ӫ�繌ψ�\�d�V��^8��ǽR�f�mSx�@r�qU.V����sc��¹v��텫�fY�S���^�կ�k��yIݽ{��퓘��q;N�1�=���5��E������1����¼���B���9h}6w���wo���@X* �s�Hf�*�����_���\��U��Q���<bұ��>t�v�Kt�Q@w��IJ���o�o��WF��)g���U��V�+��w�I:��P�9ր��H�l�#��z����矁��m��[�y7���(r�<ງ�ulC���n/��r��o��}����^x��v���\�Wq���7��,�G�:�=#
�憸l@��(�[m�<c�zViذv�X���;���.w���J�+4=W嘉�[-^3.]}��`:��S`2σ������/�CI�m��ٹ>���d�y�w���3���(�0
��!HͷO��3��ֈq��
���}�_�@���:��9�+T��^�,m��U�G�r񳋴\�(|�0;�uE+�4-�]�[j�V���_ik+Wۥ�/��X�q��v���Ν��f��Ï�~�>��o�L�L*� >
�U��EqAs|ɳ@����rΕr���a(8Qv*s��F�|�������9�3'�-���m�t���˗��o}��v��e�j�wh�8`�3@YZ�1U&
F6%R�ҭׯ$T9u�y���)aABe,��#�����]��
q��<M�x�w���4�*�Z���ƻ{woc)]o�~�Q������} � p*es�zC�\�iC�5���Ǧ��Q��/.�E�Cu�M�8��*aa�T�_\]c���KI��U��!���Zp�t_Q+~%%�$?�o-�,+�{�8IyYG�t������u�ދ��t��*15�}>��4� ˋO,�D���ijw���փq,ĥO�D�Q����oyܼ*��$3�2�d<3Iy��M��pj�or=�	��or*��eP+@�����bB��%2\y�*�)@�\��-�-����
��N�y͹Uq����k����P��`�s�Ϸ.e����m�CY��E�6]���h��'��h���a�J�f�v`P)?٤UE1��Lb�ə�(��>�[0��+-���.��֚�j��>�E�����E����*=�̼?a�g�~�����3�z\ӑo�Z�u8�~TNM��-k�)>��,t����{z-��te�Ԩ�;�s&j������Z#�������*�g��́@�М�rC�bݺ���W,�K׸d���K�Օ�v��U�e!іI����kj��q��!�WY*#�Q��O���q/����g�Od����]V�ڍV�PWfi�6�5H��[�X$�UHi��9�4MvK��ԀK�2J�;+�V��VP]�B�3�U��U�I:��u�+�x
���K�_�����1������I����iz����J���#��A:�H��@%��i�]��v>�p�|�e蝘֏�Znӂ~ؾ�~�e�
q�,��{G�`�0�0���<�ck�;�����~���@@#X�HT(Y�-��t���+0�9���g΍a09Đf֑氂�O��l�Ϲ��C݁�EjC��_�N]@���8&�-�<3)
D�����)����R^C0s�3�x�����q���@�jժro��-v:[z)���h�����}���٧���w�D���e���F<U*w	��{��XK��6`n>S᫨��������W_k��+Y���� q��U�TWR�Į������dq�]�)a;QO���-�㴶����K���8b�l��5�F�m�4����vmJ�d���\,�2���;��"X�H���B&��r%���WU�Q0��D�6.��?	�����sr�S�]l�uT��2�8�S�1\�ْص����|���Ͷ�1�#x��c�9�������w�~�7��*1��ť�b��=�Z�bcc�.ԣ0��/o�௼�j{�7۴S��Ř����9��-z��Z;�rZYt��|�{�nw
.~����t�ݣ,����<ۓ��y��o���,'�dia)P�B'�T������j��n;ѥM�z*7��K�����W�m�.V�$xH<�`�B\�R�4��v�t���5P>* �6�
Xe�f�I�,�3_
�̀���m�5�>����eKPPz�ӲP�x��g�Nӕw[��׮��_~x)���t����s���������"ﴠ�~T���r۵�>Kߔ���S�CE�X��6���i
w�򳻶AY<|���j�XU����������z8/��,z���#<�
j��t"�4r.���?�~O�)���3#�P��uUKY)5�S��J�lf���D��z���&�I��V�0=��G�m�$+%�r�O��
�F��vB�c�O1�an�:�{�-ؒ9���c��u��<�w�Z�u�!V���aև�ô���Ӯo���@˃��^��W$���e�l��k�s�ګW_o?���w��v{���+o��(7v�,�ҥ:�.�]n���Mwhþ�y.�4η5��S����v��XS���f������́�S��ݕ��:�ꂿ��Tz������:�~:Ǭ6h�u�
�W�z�8�E4�F�u0�gWө����ڕ˗��������Q�a}x~�K�s�,�qZAqΠ�x��vP N��B��*s�x��L��u���K�f����t�B�v^�a�/]�1x��C�H3q����n�+�WA��cˮ���Y,c� �[~A�םq����Q~7\z�G~��{�V8�t=�!ҿx��7���
�>i ���[�5��:��򯲚���S� Ҵ�ܥ�}��
�	���H��I��P1kp]yt��'a�q���t|*����pLD�,��qS�+��4*�a�D,S�M0MY��F &�00J��[S1 T�>Eq�t-�Ɉ���� �W���֎����Ri����T.�w����2]:w�}���j��?�Ϸ������{�ݮ��L�����CM�W^~�]�x9eu���?��l�qr���榃ܻ��e��ꊙ��h��^��>��Ge��X���{�(�^���I��q��[-���`�&����qpR\��@�;Vm��#���2���^�r%XK��Sn�i:�� ���J��b�EyS���gj�]>W�b�ٵ�lvg���V�P ($�]_�qo��1�R�|�R{��U���"�e!�Q*R]V���+�~��w���?t9�F��.
��I�x���A5�:��bR1��a�
,��%J��=�h�TI�>���svְ�Xi):t�ww����z)�̴��� ÃB+�*�Ҷf�;���ş��[y�MO۰V���l��+���*+�!&JP������5�ꀰ�w�BF�%��{b4���w�_[����ø0��A�Tp��PQ����ۉ�]������b=��0����.��^��JN=s��G���Z��Z��؍��4}]��Ar��ϯ�_�����{�7n�u�hw�v}�������5pYc �*��MZ���;e,-So��|q�%�g�}/X~��k����!3f��iz[Wn�W��L��	y:`)�HJm�M��X(QX�U�ۙ��t�\��ip�>���,�4�ԅ��/�W_~�����<����Կ�� ������+�EA9�&] �W�9P��Iw�h���liq)�6Z�K(-Wo;�T���k6�*�F!x40"($@�jg\!�-r�P���{�-���i�7
����yy[(E"�L��4ĮP����XH5"�ת�J�wN�-�������AX+uz�E�dʉ�mI%���wF?14������R�4pi�!~�W�R2��nM���?e�ђfl������%� �ٵ����!�EE

�S�R���;�2�A�ݶ�
�,i�!*�t�4�H����(��r�Z�xRBs�|E]��%c+,�R�m����]��V����>�裶��Qև�y��N�D��������1-)���T$Bgk�ޯ~���������I��?�������ݸ~3k[��hٸ�����S�I�_X?�LEc��ޞi)qR;lN�S�L������y=�20��ր�&�WH$k4��G`R@삸&�k�}ʚ:r�ɶ̮�"և�`_X���y���;�br74�&�kUP�~��۵_l��]mWW���Y����Fy(0n���[��j��[���ˁ~���/t�^������ջ��)g�_3k�膪MO����@g�}~���x��GyO��
_M��S�}£D��q(7���ΒS���՚5�Ζ�豆T�'"�Ì�n�1��-���)��
�Z'%������׻�i�@wy�8�r�Vnp�4�T��λ(B���!L��<���M��Fe��T�2�ȸ"�sR�V�ܥɷG|[g¹,ٴH��@��u��]���4�0����@��*����w��#�9Hz���v�����~�<�H���%pX9G�j���
�Dj�mY5oU��[;�����]��p5��"�&�sӖ#������v*;�Ӯ����pQ����7��ttQ"�/��R@Ș-�U��я{G�z�_<���$v�=~�6���l1��ni��{�D��W4�=�e�n*\��=x@w�z�ӎ[ćĴ?��E�}�n���~vN{����F��$l�:wI�8:�zE#�U N�[by
��~ة�V��써u�H���A	�\	p��:eCE$���c�Zi]������ur�l����$D�C��饭t֢r���+�ŗ."�<-�������WnT�!@!�,<�N>9YQDP����)W����������*��N1-f0�������_��06L!c7!�g%y�����2�S���0�x�O��Y�z*�	�HMW����v��9����b.`z饗ڛo�ٮ\�R�)Ĵ�.�rL�V҃u���Ids���h~�q^Տ2�G�.,�Z�0;D����Sޥ�/��R��w��~�w~�������'�^�2���Y1~��.����K��ta.p=� �I�&�E�2ҵ��R�d
�F�͋�] +H�tP 2���\iz�ޝ�����r��a�ʉEf
��(vu��r��/ۗ�oХ{����~=�֞FLu?w	���w�_��?��}z�����[��G1`AK����B� �<�n�e,�*��@�?����_�r�kP.�,�3J);?�b��]g����菟5#}#�VW}Od��ϦU��SPqk��rU��+�C��j��;���1�K�:3�WI�T��D���
�D䡊��R�w�Tr�:�L5ꛉ�	�����W2�i�����\���h�¡|Ԋ���!g�����`h���F�� �k�����kÈ*��(���|�&>Bi�Ѫ��@w��	�M�(�* +��g`v׌�/,Y�r�=Ek��9��l�y�v�����i͸�ai����Տ(-G�5�H�թh+7�]�rY0�����Ɯ����Cʵ���^����߮]~���8�	�G�{;��7��g�sڛ3G�c(�����eqW��:�>v)�Te�yµ.�'���3~�\J�)>��~�:A��n砦GXs�<I�e{	����O}��&כ�㬘��BB�q( ���z�91.��~����&9�29<�j<r��z���n{@7r>Ytz�����C�n߹�F�����(�:��vi�p�+t�O����O"�f�l��m��c��f�<I�:\���vn��IHyW�G��C���{�RN�	��Kޫ*u%j\��xs�n�*���JR�mBkW햵Օ�Ii�1���-��i#}��n��3/�n���$��+��V�>0$�W����\��V2J�<�|�N���e�iG��M���˴�0�x�+��&��jY��;!�8t|�fa(���X�0/��Eh�	LT
p�^�u*qu�b�\h��(�����x�����m�o��ݱ�X��]�)��hd�}���%�2Y>�1��?h�~�~����ڇ7�l�]n�kmii�]>�"Ap���܄�A/! �M���'�ޓ�6�|��zAc?2��-�Ƌ��H׊�9B	��}�6�=��r�f�hE�MiI���8���Ǐ60��^a@����Es�Ԕ����*4�J��^d|z9ƒ��h:�E�c��hb:ӗ~�r9���b�jI���m�;��ݗ]��1�3�c\�*٥^�loE�9P{������(E��R)��x[]�kWί���Kmmn�-�"�G���n�{Pn���$��x����S�SX1��c��HP�ש�O?��ݹ��ݺ��ݽ���?Zo7��m۔��'�������M�:�K?j�y�&��=�������Vh8�|�S*H�ֲK%[z�z~z*��.�[�LiQ�̞�F��)�R�z��3*�����q�yz�v2�` wj�	?�|@�#�ˆ+��q����^l+�Z�5��?���AP��^�H�E�BW3��lyu��{��ɨ-L����T"SН��X�^�ƌj�K���c���e�Q$��6M���[�w�ojd%�B���@����
}��\(��{�����?�}����az@�B�E+�ՌvaT�Z��ڑ���j��n�hG�[(����/��b�x����f���.�r7�G�M������,�3M{�.TڧN(��0ô�fe��f���a���a[^�D_^� �]0gE��p�LmH�U��<O7��][�L[��\�~���"AH|o/��Ow!/�.��66e�;n@+��S�Eq�G3E����.�`Z2�V��۷s���3��Jk�֯a�k�����]Ěp}��~O����(fW�g��.�Pe����14sq�)�1?jf��~~��>�ï����t�n��=��������B��M@�!��w>˯vŵ&"xi�|�şt��׎��K]u�/�5�qt�n��Je����]��}d�d�.��a�(�Kje�<���	oy��ҷ\�W��;��H�i�o�%�?�:�� ��#1{�R��9��c�u�6?�-���jΊ(�T�5q3�)����1e�gq3d��t��hvo���b�~�z�}�v���Փ�c�9��λ��V;����A'].O�R����'�l>�����6F̹��:�z�5ZK[W���|�t�*�m3�G�{R�����ή-0�����a�-ϡ�b�Q6��JRXL�����e����
�{����_�9;Uݿ|�8"4=@�0<BCuǂu0��� �����:��F�u8��z�:�����gJvR�<t�l��+�Z}� O�{,d��"�9E��n����X�]�r-3<���mաV�Vx��uEq���:�yx͙9�`ֿ���6�1�}�Y�}�]��to���h���2J_%³�)�Tv�˴������}�ީ���)�p��ӠC��}=�;�5�U��)��c�k�B�B�K�X�������j��+�	e������J�U͓=����u�^2�~��q*�F���*�7��Ϳ!}�Y��7+��$N�����������<㝄�ZBW�:p�̈'�?�]o��l�w����L{�o�����k��N�=���.�w>ﴟK��s".�j/�lxv������d�Q����gv��"��m*�1v�!ݑ�v�҅6�VS��/�m��w���)�V�o��PAT!������y�I�c���y������c�I{��<�7��ow�L���~�Mk)-:�n�%[�
�
��h�Z��~Q̽
�oԺΣ&]�RV�1����N#:(��Zͻ�tg6a��i�ޥܵ��i��M7z�w��Q���$t��WZHR���r��������J�v���[kw�� �8� m��f�X�q�=���:��^n�����ݛ�X���Kѵ:4�-_)�X:��T,�����i��q�P�����y�{���Ga�䩠��~�j5@_ട�m�P����=yLgw� ^R���0����w"+��l��.<y�%"S"�g��p�4��E*�	8_X�:�&I�/����_�ǴNB�UV���Ld��G���Z�wi$�J0}h%�`X�2�����'�?�ϼO7��ǝ��͕�_�Ҿ��7�|+�&<k��a"�t�Z�z���	���
c;�����2�����Ӷ��*v��n߽ٶ<�
��rL�)_�#��j-9��%C�S/�?̯i}D���|{S|�a�8���4Р��؏Y[sw�"]��6�N��Rw��x�}�v]�����w
�V����;�m����>P ~�N�dw�V;�"�(q�E�������n�Ję#��2�v��h��*Q�qu��3T.�����_�_����'�f��7n�8+[/���V�}<��.�{��Q;@P�Ҿ����}a!ݠ˞؏�m�a�L+��j�A����H���Ҋ��P��4�cu	]>�I��(=�ݡ7����Uz������~,�:��Q���A�7n�׳A���0^�lT�PE-H�0���/�`�bv��@.��S�*�LZ8�W.�@��T�i�%f�Z��X�� ��̵����M.�,d��P���
W��Yԣ�7�1Y
��kEW9�/^S ;�K�����=��>��q�����ߦ�E��eS���R[�]h+.r��b{���a�s0�����8Ck{��VZ8:LM�v#>���l"�~�y��ۧ_|�nܼ��=��p����|y�F�K�\S|��'];��X\ms�m~֣��k�g���F�\OZ��'��P�+��8wa�tl��*z[�ԥ�5�h�<X���U�;�DiS�'�/ve.\���gMl�4��_�F����A�y��c>�X%��=pl��9,Y0���k3�^��(m�I����'�A�n�Śy���'�}�~�F�<�!�sLV��҈�I�,���GCHɝ-\vvm�AD�`���*�:�h�}�3���
�A�Tq��BW|��9^��i�N"OE��W�����.����e1�p����I��S�kø�cA�.OIrh�1)���ρk�B��^�֋1�o=�(��XT��m�5?_�0�6r�g!"�@i<�6�+%��C&�~��U���+�p5�D�BL'�H�+��ke�$.�ć��`�/u�V�p�idX�A,��(�`�=�~�>��W�W��>��y�+z�� �չ��./��p�����
B��6�Ç�X	;��o���v_�R��~{�r�q����w1��g�Ϣغ:� �xF�Q�*�C��q0�*�!������]Y� q��9��K!�u�&2�g�����ER��ִ70Nƕ��\P�j%f=���ɠ=\h�ρ�U�"DIIc�H� o��- *O���(-��iKO�w��V��Hi�7۟��� �//���8֡�-*J����� ���G��Ϯ��5 �ck9��n�sZ>��Pkd	ˡ+1-bǛ,������%�匳�!�m�T�(��(<
k�o�(G	C:qa����z��;�F���`��7�Ʃk�?��;�
߳UT
�zSg֟)�p��}Y �i9�>��j@Yt����j���G���T�
��ԮV��-��ن^+��.��kp�L�LE����b<�0B�ʂ	���A��	�yv�L��f��#�x�nW��S���������w5(-!�H�/P&�{����M��}�^�q�&�_h�>�~��}����ڋ/^k�����aj?n�~�Y���m�1���l�_mSc�-Wiz�~�����q3J:�3V��F��`i5آ�
�r���zQs5p���v����޾�8X���J[Y�DWʙ��|0��Sq�kd=8��.����ҭ�:��d�G�g]�)��z}{����V�h.(�U!Y�+W/�w�^.�r\���
Q��]]#�U�U���fHg�D��b�֮E����$>�g����p$���Q��T k�w�T$���\+��Py8�q>��U��AL�4g��]����~b�u5���x�eQI;(�Q����������n�� �ʪ\KH�ɬ<�gC焂W�o�}Y8�Nd�蟔B-���({��ҷ��a���-R5_[K�m�f֡xʟ��h[��_��2�OWJdp��i� �#���ݨ��	G��Ѕ�΂$s\g���S�Zq�h�"}r��%���2��&���L�A1L��#ϋ�jO6��o��w�����:�YFm�(�x�4��inwi�f�]]���q[~�E=qLK�V�.���ն<����վ��zZQ�����ϭ�=3t�Vn������pɱ�u�G���o���XIۆ+	)�և�r����a���I[_wt��R����pveV�K%��k��?E����\����z�O�2�������ˣ��cY�b9��a���ZW��7�|�}�?����i�@�/��-^�P�5����hn7��o��V{띷�/��"XK�J���6��b����1N��µ&��vl�3U7�ki�n�GO���}h�ڎ�m�ͽ���Mn�p���.-|���G���]h~���
�O;�9� �S�+�N*d��r+�Ι�8w���Mg�/����<m@��w<QU��-�(۬1
�#�O��n� ����<�~C�	��i�$��Am6R$���
�Ofq$��F�pK.�N\��V�F�5S���4^�#���G�!�`���N�s{�	��Cɝ��� �&hݞB4�96�n�{W4�\g��������MЕ��^k���ڥ�W�^lk��*�я*-Ғ����b�ln `�<���Q�/���^��^y�J{������%��kP�{�wn�O>��}A�֝�t�w��<�R�0C7��_8�^x�
-�,~5�*�N�Mwy��hQu��NZz:խ����Ϸk/\F`<Nr;erq�P7�����۷��v{�W3��r�J���a���l����/����1F�LA�����J�uk<��:S TJξh�i���p�j*@�:`1h=8�t~�B�F�n���ϾQ"(��.d���`�W?u�����ex�1(�m�=CȒ�R$��WU�Ҡ���s\�+!��n
�^E$XP��uL�"DZ��I�FɐcP�j�gC	Y�ҭ���%3����`
K|+�7u�b�f}KA��a�a�;a��EL\�$��ga��c���/��b
ξx�,T��(�F4U���CZ�/`�Ð��O�������v���v�1�d���V�SZ��.�K���mZ8���/�[/\��^v�(]���[E��H��	��Y� ܿ��ݹE+���Na�,/´K�_mW�^io��F��w~���������������]����h1���?�I�����?�G�M�����}��GX ��O	]�ۃ�4I�W�]iWQ"�3vq\ ez�~U��Su��>���
[@R�e�}h��^y�E��%��6�����tP��ܿ��>��:tx�)Y[���Ե4R9e�d���#gp�Xl��OI�»�������Ny6��Ĺ��ߕ��-;���S񭞫���q�b������Gʹ&��C]�GN-g�Ɓ��'g1�c��#���k(,M�g���d��^g �Y�����Hc�wW��g��� O��\}��\��J�� h��7��$�V	
ܔ�-��O��߳+%�g
"�k�XA�7�$]ekA*��Lm��00����a�B��Yx�F ��+(�/&�]c��A�6���u{�o�Вn ����7ڗ����X(��tSP"�)��;��؄������_�r�]�����cg���  @濳y��r( K��0`[��)��B{��嶶�6�%��b[��hc�H��i�Pr�(��[w����������������O�E�<�{�jz\3��1����U�AziQT��A(��ZK��z�/� \,h/&?g2�z^|�
�p{��ը�]�#��}���������c����Q��]�F����2�URv+S�܆��N?�&��8օ�,�0�	�v�u��jc�l��w�?��/]����
	�ey�(�~��P�x���K/����q�<�l�
CE"_y����u7��^{�[tW�b�@��w(���k�E�6?�ZZ�#JR�Ȳ��5NE�Of��IC��~���#��#J�ժ�,����J\+�2S�H�JB�A��C�D�8U�z�M]�㩂�m�6]~�k�犿~���*��X$�7͞�'��^��,w��"V��+W��2�~+����o����Q�����{�n���F�5��Fv��]y3�7o�n~���q n����m���BC�w�G���4U���D�=.jZ]^j/^�J��\���to���w⺊���v��;�O�?���������΃/ۣ��(��������g(�[���r+ Hu
Ա��^~	�~!].�n�����6��D�~ i��E���>u(�E�k�����5���/C��D�λvkN�ϟ�>��F��O~�~���~x����J�2�NX�H��k��4���΢Ք1�Iz��3KU��Y߶��������
qfI!R��R$𠵊������5�ȕ�ʋ�Q�Hc�w�x��������K�����F2�hk��9m��/"�� �T�����p��
�u�\W�z��.k�
1�՘�U��I��_^�z)+F�� ��cw�Qc-#�J�$�bʂG+���50�<�d�����p�߆Y@&�_�t�0	����/����� iW,��ɑ��2���F�?#���ի�[o~+� ��㘛c�1��V�}n�K�y��A�Ccerp�����f�V�C�<|���C'W��Zd&]��'IK��5ݝ�e�����oĬ,����h98��B���2��΃�a�/?�������x�}z���I>���ʬP�=��G�:� a�Ofvn�]�t�����9�K�D8`��B�^�+ڗ�t|�^S��	��� I�l
����/��%߱ ~W�:ȩ��>w�~��'�����M���nW��W����5?���b-d��e+A���mqnvrQ�$��n�R���U@�M��n���_~�����*����h3X֋֒���o��#��V���^i/_{��.b�L�~��iw���7���zp��E-Ae����.]��ʃk5�ܓ�ֿ�2����E��OA�3@Y�Z�Q
��f�\���U��3��n�a���0QhSv�c�Ɓ�J­���N�hn����/`x�����_��W��c�V��d�(�ڵ������QQ���Z�,RAS�{�����p o���Y���r3����w^kW��!�[�A�&���=5��AJ�7���{��vMN��l�dܛ_|ٖ�g�����W�$�c��37����;�t'T��)�_[Zg+wS�RLa���`��lR^�V]�n�ݥ�a�H|�\*�AZ���_����	�J(q�HE�p�a����v����V�>���Xqv
����6�7���������ۯ�����._���>�+�Mm���^��ק@�֒��V8�(}�O�T�L8��׌���]��~T}Kk-8~�ɧmavk	a��9��p�z<�iۛOڃ�b�\�����)OM�i3�l\��
˵Օ���/�k���Y�u]�����W�^�����N�*QZ;�v�]�}Z��^�n��:8.~����]��ƴ�D�C���a���x�����`|���������P&I��6N)w�O�4�����fsQ����8����n�z���<h����*�	M�R>�j���SI��d��&/��u2%���pz�����}��j{��+t�fP���e+�'��u�����Ց�=Nk�7Oon���A��%1`,`�3$\���5\Mb���<F��V�r9r �d��U �Wv%B^��~��cZ����e�0�Y7T��S���! @���&��1��mP����a�Y�'	O�k�w�VE$��*'��fP�Z�m8\�p�]��_���m�ʴ������Ab�;�q����h�x,�&����
r�o|��46ۃG��'�?n��|�6v��q �zhe���Pg
��B(q.~ZZZi?���j�z�v��ӝ.��q]�����1��7�����[��j����ZL*3�'�ۑ� c���Z\�aN�e�a�~� �R,�L��w�"���Ց�d9��c���W��X/��݉�X�.ֳY� ��=yd��2����+�ܹ�����btG��_��Bq��[
,�8��?��~@�kڏ��Fv�f��ٵ���F��zL��b��k��{����5U�U��.���f3( �#�EH-����0�Җ.�����vUQl~șp�NȌ8��L7�D�� �8��z-Kd��QV^�B9bҊ�c�����_j?x�E���6C]�%�7q�1���i�wjr�����ݏ��Q+;
�)-�ZZƷ�Ց��Z��;/���!"��#"&L�u�Q�A�;��y�%Z��+�~�a�H�-'*U�NP����i:ߏ�a�����eiP[�bj��V�I��A@+���ϘIK���k���I��#������\WPX0�:�y��y��y�
�E�����M�����wf�/o~�nށ���pP�%%��a]ݾ�����.��tl&'�����o}����h9 ��:s ��t�����(,ZR�6/���np �j5L��P����T�3�ڝ�k�T��Gu�+:=c5�!�f�gl��cSN�;f�x�-�'�;��Rz�.\���o��Ţ�q�О	ݏ��.]%�-���<O�>�I݃���VV!��Pae��Ӄ�%��m!�Z�Dej�zS�=\�nܼ��zn�}���i�z���n��Z���6��
���1�	JdJ�N.����v��f��?h�6���Z���O|���E)i��o �3SU��5\*����3�)�6�~U��ߺھ��e��ͧ.�3���_��`�x�r�ut��f��}����ۗ6 *�RЮD,�Sd�HZ'��vV�%��C�Q8a��1�YO�r�GY"|qi�������.0��
|	�]�ޟ�%Ϥ���yUs�XF%�'�Ѱ�<���K~^��E��y%�������z���s�liQ��W�b���B��3`�j�h�(����/�����ل���v���v���F`{�I�=B���X��NC;���`?\���fR���)`��G�����W�2a���*[V[Rg-��B��+��d�T�y����3p��ϐ'�VhB��]>�ofQ&.�v�І3e�3ߺ�"t0�b.5�A!�we�%N6��f+~>9��!��(���l�Xkz�����o<�GO�/o_�V�:Q��8����յs��������F�b8�����'�(���cylPG�ۍ[_r�զ�&Q �wP�Y{B����'m���a�<O�xv�������,�3�������T9Wu���ݍL$H$A��Dej���F�,{�e���kfl��ƞ�g4�,J)���$HD"5�ht�Ft�\�r���}�}�Uu)��o�{�瞳�>{��IW��܂_���Mŷ��R�."g�3*�AI%���/���J���Y�W/��b^�W"򂝯��oC�V��Z[���ێ���H�dx���}"f��!5i�K����[���귞�S�Х���ia�"���M<��W�G)��(�V"\K�L��X��b0�?Dރ%��?����dAL�σS}��)�%��{]h�����A;s��]13*�zѭQ[Eie���h҆$�w��h5���Lin����橖��!es�z�9[RK�NT˩9��B����9����t,���m�U!��E�����E�vO�HDV<U��x~���8v�x26�W�5i�k5ڢ�ҥ⥠�*��3�9�H�T�Z���f���q��dփ�>s'w�\�;8��V��p����_�B�MCk���
�-��+��\���U��f��d�Dk#-4Z�Zq>�a�;V�Ҫ�T S�qs�+�Jd��������Н&}�^tMc~a����=�;e��w�T�.�Ǣj���8���%���Q<�
�+SѶ�<R�@�(����lkF_�p\���>���_&-$�ӍOܤH#]y���"�̬����?N��ّ���z#Ѝ�!�S�ԡ��DT"��r�R�vgJV Hm�R�i�-�<>�W��d\��:@�c-����LLS�B���I4�+lZ�Q ���kbH�Zv,��D|���!�����c:X"H5�K��"�A"�EZ$\ہd˯ g뿴JE���m&�ȫ��l��0��)���y�_*<�VC{i%h������n_��7o[_Q3��uZP[�N��|*'D9Sr7F%2���XC8�b&��7�¥��O�s?�cЍrq������ ��թ�N� ����HYO���҂+��P�0�Ƕ"���R�:��<�
��>����dvo��x`�� �������mg2&��:����Z3s���XFi��]��qKB�
�cc�0�T!����lE��s{��J���C�4�k���2�����VI�h;�U*.^@�L (u�'����^x+.`-F�J�@�~�-1<>L��7u���B�Ǒ�?��I������ɉ�x���Dַ�~��d*IK��P��<�P?���)_2�N��u߆)G�#c=q��P���^���|�eV;���H��ɶ�]\^�ǿ�|L,�3b�#�x��'.Ss��>-�2C���� ������'�����{Gbt��Ym�}*>e���-k����R���؂�D�H�Vs��5�Ъ\8{!'��]'89S�4J�\�i;���^]+[�ĭ�T$.-wRS
$i�W�Wc-��k�`��"c�`���O��Kgi�.e+���nG��N����j�
�뱑���W.�a��C��q�(�S�irG�=z�"�1d>�Z+�t(���C\���@�khA���N|���<.ז:w����ݕB��}ex��c�֠���3j�|W�V�pߨ4�P�(�
���U��R�����L��8r���%�2�����J�f
KwIr�
.��ܫ�D*�K�/e��Z��$f�%ru�J��;�ފ��8~�h�<u<��Q�W��&]��D�T�H��|��	.7T"���h�@�tĥ�s��3��D�3��i��N�NT��yVr^��� Z�~����D�����������;O�����3�0�#��rmg�J$g����r5�6`�I�P��<��+�D:hE�xtz��Ĳ3
FL�$�Q� f���Z u�2m[�Rt�7��D( oa>���o,c�`R�r8-ݙ�n���1�I�/S���	ސHm�؉�;t��y:�ٞ�i,�+/��բv�M�I[H�% N��=����'u�}Q��p�~N^?��聊R�Y�axt(����ws˽��O�س�����2ndN9&o�W���3x����cb�*u�g�=��~2:���+�0��c�b�2��9�4\ۓ_�j�+�޵_��d���돌S.����L��2�52D��|uS��q9�K�m��%��y��oߍn���3����/g�ڒ#oy��i�.��am���*�b8`��.�i�TTL4�N���/�])]��Ts��7*t�!��]؜|�;،#���܊��>W�֡�}Ok1��|ɏ���&�W�mf�-��D�v �13�/��vL�.����4Mi]������u�]֝VN��2��y�`��Z������d��+���������A���HB;G�L��T"2����Ddr��w�������>�g����A ��t(	.A�p� i��W
l?A��cǪ��S;Y3KY���1�S�K����fﾑ8~� ���x$̆�꼍4�E��˴�A@��+����������5��.3w��u,�agq.~�l�N�Z[�A+�;A>ͽ'����u�+7T���e(����*��������k/�k����2[��5Mf�oƊ,*!@(��z(���P�bq�;0'N��=ô�`im�'��[�#?��ޫ(�Cf/͸.��B��s�y�z���W.�lq�?��_6�S���)�N
���e�*Y�I���K�g�^7(�n�g]E���Ǚ��\��h�b��}�����M��><�,���3�w���;Ή�<�ThM-�W
������[��c'g'�.LYķJU��m�R��I��G�H+���W��]෡;qg�7q��L<������X�y+/��ϴH��YeBf��C�Td�������+����ew���oo?2�C�c�}Ѥ���^7x�,j%RZq3q^�G+8�ɹ������r�'B����Q��l�dZe�Y$�d� m}�)�d� ���?�Ej\·����?�ޯ*-�@�DҴ��]�Dʥ��'C��o^+W�ڟ��7y�e�.�*Tɖɷsg4�wtIȡ܁����i�R w���+DҜν+I��$���T �3^z���4q���� �Q�d|����6�8\��G��A��щ?4:��Cq�Ⱦ8q��سo,��e�$�9�
���֥��P�?	��ڡ��hX����r�^�����U��Ry1[�L����V����<�2<2C�9�Va�����q��w�_��d=�f��\����ɲ�������?��͏�w��cb�T2i����PO�
uT�~��Ŵ�4�����$B�k}`4N�v,n;}k����O���B%������*$=�(2�43��Ah;�9:��֊�W��_�y"[N��U9�T��ڙ��m&��X���)��p���L�<�c�ј��nx��K���}q둱���ƅ�$m'sj5Y�fQ�3����p���./�귞�Ӌ�J���sz�&~2��H�8��� _
 �7V"v������>��ԡ̊���1��?zl��w�")�*�
C�D��u^咣£�ϻB�r�-ˬ��ʰ���:���*�\S��3�yMER,?�048��<�ˠ4ڰ��(;Kg&�'�sS�^yf~"�_>o��Z�Q����sU)���ˍU�w�@JS�V���Y�����ԭ'���9#�N�ZQd��Jܒ}�[kD7��0�rH0��&���ke����T����(���L���΄8�|�]<-:C���#"�u���8J�f���I�l��KޔCe'��V����5Q)	P�($/i	ml8��M�Q(k(+���j�^�����I�����q�������B�X_9� �v��츭���_�M$Q��p�7R".�s�f��7z�qyg��'������(�2�����뢼3�r��F��!���h�y���|���	n��m;�ֈ;��IwfKg��㈹�lɦ(���bq�ҥ������񧞏��v��!�T"�F��W�$,o�\�K���{�9�l����P�b��V}�o�ǝqt��me�MP�-���Uy�t娯$�����;M��B�/���:�X�U����\w\
'R������0�
X]����0W�qq���UW&�����w�y���@Z �S��H_�k B��	s�-�����=#q���ciQ� �
�r�z���%�D,�4�V*�Iw�^h���F�X����ذ��S�N�^]�5���p���U#�K������닜�:443W߾!~��c
������I����br`��_e�@#���I�W��\���4V�@ʮr���ג���q���8z�`��C�����"<j�
�(����T�n&e��
dg*a���wSK��AC݋���W����߀��pqsj�z��1�F
 G�e� �����J*�(�x�(���3�W��W҈{n9�u"F��=@�~���2i���D�� ���w�z'�u`U�d3�`�P٘�.牤�(�D����z���u!���H��C;Ղ����Y������\���v���LX�ǒuѷⵍK�Q���S�ć
OF�,��~��/�	-\�	��e|e�$,��B�?��8������\��+�s�r��9~r�2.��Y�TVy��߿([K$G)(c;��ܐ>�!��u����q��DW����')V�Ӕ�cю�9����Q������_�Vԁfٲ)��\�m`��ߊ4���fy�\����8Ut�K]�T�(��풡Lʭ%���Z\p9�������*	�>,�һ�Ҁf��[��-J�V�2)
%;�0]�K�M�p�<��T4��@W�AI?~8n���8v�pNco�:�Fk>ltcu��K�k�Y i&/[��uU��D��Hy��fJ�mhR�+Zq�rqg�l���J^�.=�~Q&�aVE�(�%\^O���p����C���.����ȃ��ĿF�vx$'������r��<��w�&������y*�S�����K�Ź��b�PPg�%RAf̣�Y}2�깗7V"%���Yd(�Eh���)8���(���(8�E���H
B�s�ɜ�)W����#��r_D����	ɝ�pkTǎ���h��O�ٽ7�T��q�3�n�]���V�#9��x�$&����<37��pc\�礥�)*��DJ)��fF������;o��g��aӥ�KE.����K���ͨJ����5y(t�XE�$�n*Y��r��w�������5�V�r�}�a�y��(\*)���0L7Nk�>����Z�a�i���.-�B�b7�r.�g[͢�-�J�2H��o��P+��#�@%�ػ�s>n��D�>=q�X��L�w}�
O>s�]�-;e�I��<T�j��r���2 ���X%"O����3���H���������`Q���BJ��y��P���i��0j/�b�H�y��v��X#�;G�)6.�(J��gN��'��`�K;�+_��H��vg2S�	����Kn�=�«q~�/�c݈�fW�#
��7[�,HI��d�w+����cڹ&~
�NI�*��7���qj.�2@ ��%?�U��2��g*���W"�@!<�WH.�"���km�t� |�G��cG�>��V���nݘ�4P�nN�g:�I#�R��%M��+q��٘�p͋Ç��Θ�ٿ�.V07/6 M��4~d_�z�6���{�@�GЂr�a9dr�8��s�'��j9Ay~P��R2�䓹y(*h$}��C�5oH�Z%�yG���smb���P�f�VC*�:��9�2N
#�����x�)�~��2��bd���P��Fwo#�U¸z��+k���N�R9�P���F	��G�C��w2`����8z�H�²;y��8���m�j5���˄��*O��T�KA��
eK=P�b�\�'��� U
.~3�&=�8;�)3n��F�\�Dhciyw�5��ʉ��I�"b��Dv�CP����l�	NF���@�en�
brD*/���'�]i�R���
���N���ǉ"��;�[G�< _ydIIH$qg�<oK���O~���/��e���@���H��"xOST�r�[��P[p�:��B�Ԅ)4��T(ۡ"�=��ݚ�/���.�&Z�4�m��'��{�"���@+=k�[���i���HN��[R3�d���le���� ��p�����+�'3��x�HI/�Ӎ��¼C��j�MŪ��/[)A����N9�4�������6~��ŌTP�H�� ���+���p��')(7����xM�U�Ω)E��2-����w���Ƶ�
#U�$�ʫE�-a��-��C�r��Y*�7<������ɼ9;�f�Z)2�u��8tud�tsn�JN$\ZX���e����l��Й��������A�ӑ�Fot���g�F�W��{^Zl�x��ԧbN@��!��̇^�$,_k�M�׍��5Eg�Xu��U��Fol-��H��x����_�B���"�l>��2?y�<lI';ei�Ra�{6Nv@�&����m�H�C��L��(rv)8�}y9�p������?�Ïġ}R�26-W�:Zdq1HR�X`�(�?�B\��&Ϟ����o��^x;���� ����wS�a��-E2�R�hNIwG-ܣc sU��_DK#�j����]�K؏q1�i�zL�NPЅ4+Bu�%��Mk$	�)e�i�	Y`C��yk%�Ṅ���:��^ɘ�0s�-;օ��.,����a��(x.׵Q��{�1�
��U-����.y'�4�_���n� ��#cn����ݽ�XW�Y̲ ٓOX���b����Ujْ��}H�j�N0#���B�a�/����<�pti�(�,�����I\8�e�aQ��r,�ʹV0΀��*]9�N�8v���pF����-?�����A�I�e1J����v�o��7?� �TqZ�\���L�|H^.bk��Bu�y)���ѥA��H:7iT�cq��j�گ)^|u�x�2�/-�t�H@͂壱�rx�P��TA���(����������;�k�������#�����T"m���m^��Eҫ��)�Ha���;�֌'�{9޾<�ʹ���j��������T�"��׻3j|Q)p��!^]U
(e-F��� "��c��!q��0�?�-%��M�5���óY�U��?+��f�l���' {�9kznw�W���.�j�7�ӳ�svS.��z�������F�G� ��!7�9�/;ǎ�#���cl�X��tu���rf!ץ�Fs&��б(�K�-�4Hꖢ�/�Z��Q��UZ>���|ҧN� ��4�}}Ժ���N��RS>.��Y⡰U8	�!�5M|�kG��@��e�<�]7c�:'���K��9��ʧ���Nt���v�= }uT=릸�Ү(�^"y=+��QOy�|E��"�k`i����}'._�;B4��}�M�	����['�"W�+WuJ�cٴZ��)QJ,~�l֪�;:�'�̟�7w�<�� +Ks�u�n:�A�̒��(y"��DX"�a���Ԯ�'q9��!�#K�����*1�a�^7B�5�p�a�{�A��P��D��0�6�T:I@��k#yM����`euS�(�-��;��la:w�G��3z���7҈}G�������~|��GF�Љ=q��#qۙ[����'�y�L�y���;��ɣ���!|�n,��n��o��U��j�죰uͺ@yB��J��,��PT��|;N����ٽ=I)
)�2aa�"p�vMt'�����yxemX�Y#<Sȳ��θ�Y�ԍ.[�f����F�),Z�ZD�]��.iHM�]�|�{�Q��:�|E�h��3}1�q�΢]hυ�	YMIw�ɛ������PS~��+�!�!���l��� ��� o�n&n.��I�4���r���8'��"�tL׳��&줭�w	���T�r�@f�d��f�0�D�-�'��r�F�����a�0U�er��JC_��ߣ���)/�!�;)�G�[yӟyl3CI[B��n�����2��t�1�ۀ��^��W½,�J�+��ՙ�X� ������7��ǳ��g�]-�J,����lb��@�l-���ҁL���Y�M�wv�L�^���ڮ���z�_Eo�����׾�
�и���U��O��2�_�ï0^���sI���amU��_ �{�Z8#8ib\��s��ı�5�@C�m��W��-t�P������ ���߁B�kˠ��{�!~������4~F忸��[`� �;������v�S��lq�����se�u2�,�'��>�\T�Ȝũ@��3��u��q+�b��G~����$X�)�U�^k9�;3#�>�Bm_���O?JAT9O#�W��0@呋�8���˖8ߴ"�#B����%�0E��c������k��M�N[�ˤ+[*[�n(���J^�1���G�z�t?�'}	�����48Nu_�٩�	�W�<�-;�:�������՟��<�Zƶ��)۩��w-ĆY���!�T�|���9ė}@�O<M�6��7���u��:�)$�ʻ�'��Y��. ܺQy�6[��-�8Z�Zk��"�*;꭛���t�
n</
�R�eZ�8P��l�ZQ��ɾ�k�%\>݉é��R��(�X������iT����7MgJ��ӹ1(
Yu���٤��Sߕ����dA������9i�G�X{(��F�rL��M�Y��C���!��;�rX$
R�YA3ػgO
���f�q�B<���������5x�gmj��d���zJYy�x[W?:�J_׼��'#�C�%��Ix�t�P�yx�䟤J�=�$\�d�d����*N��fk�cq���bZ��ȽEL�y*��f8+i�����m�j���Ȩ��b����]�DY.靋 �L<K�'�佐e����EZ�[�I)��p�;���q�a�����I#�����T6Y�XH5�⛸��R)�$K��|�tM�tvA�D�qy����!~
��$>�;�}G��
���|��dL�xW�Y���Ǒ������J�
HW����QȊr�x*�)��R�{	Ϸ2Mxk��N�ny^���@KQ��o�C�4N�'V�Z������f'�B��h	VI����S>�.�ᗧ@���2h<�q[v��3�eѳ+�sc�.�/�;����ky���&�*x~��c�r��D�C�,���<�%�:�A��!�(2�����-;~-�"^�V��1���U��!��:���
�=����� %K������?g�¸V@~�&+E%P���/�U�Y�QJ[�|��E�?�� d�l
F��5�p�I)�B�9�a��05���g♦�w��k#��:���VXe��ʶ���k�)���Ԕ2��m�mu����c�~���]��N�B��t��w�{m�Gy^ũ�����$T�wǭ�LGi�n���g�dci߅�?8�jvGO�-Z=6�sX'�х���Y��W�Fݑ���e��H^!y3�(X�����c��B9�Ѿ&^}ɹ�L%�&�&�ƷG۳Ó����ʩ�S�a�?�a2���SY���~N=���E�q�ڼ�y2\f+�%OyY�E�
+�@U�+B��W�D��S0�T��K�s(��B��ӺH�hA\��R �/���I0�̷�%��w��G*���kA��
Ҧ�1vʐ��(JoGQg�Cƭ�ITU�+�xҹ0j�W���ۭ<��lMy�`ҹ��6�Uu���}N�����I��B���L�r����x�ED���x^��
M�z��-!z�����A|�n�u�=o�n~w�O7���m��}~��͵.��<V�i-��*4�@��Yj�5���ٴL�<��>����ְ�o3���"���]ɇ^ׇ���S҂1���q��՜�k�N  �����Y���g9L���eJ�Z`���	��3�|�����Ez$��k�g* ^*�V`���r+�:��h�J��44�U�*S�U�,��Jt�X��tJ���:|��'��}泝_y���H� ������-3�}m��׼0��|U���Ц�lT�s��ӫ�����Ļ)����Y�\�Ae}����F�� �)�uM���Bґ���|)��uI�k�U�����UʣV��{e����a$[��;( a�g����]��ju������q���x�='���'o��~�gxǥ����ߔ�m܋%Y�4����0p����%�eZ\��ҩ����_�ླྀ|�R���>�8���:C�z�R����ւ�4����R�a�C�����$FV*i�`Z���$JI���W��J&��,*d��
�qȫ�}�@���)���2)S�����f�~�0bfEo��k@�Գ��+�+P� ~����2��X�d��:�[m��Y���T+��ؼ�\]���`~׃
��v���ؾ��v����3\�S�����,/�xo��y|-�]��Xc��.<Wೊ��>���)�E�h]�i_��[��B6ή�*K!�bx�w�}4~�c�G>zw������G���݉"эvG=WۈY��U(ul��)��/��ڣ����/� ��2���[�@�a��kh�Z�����(�u��S�)���i� ը�W��bݷ/��ٓD����1�e�/-�,pŘYх�Va���*0+�s����n���ôx�9��
�ԙ����$?`'Yv�A��d3)W��A� �_*�l��<*3�e�ʹ�dr$- }h�e���VC�:����-w�>�.c�l[j�� <'��%�N�]����m$�	�!�r&����<�H�ymC�w3�>n�}�uUAE��\�K.-|%��q�(���c�����\�U��9�(y\��(7�^�V��0QmS��6���}���=~��M��K-zRH��pxhʽ�I���P�}.�ƭe=��3)E�x���u�(#hv�y��{���L���L��X��*�?��V�;��\��A�s��C�N(\�����aKA
Q�k����Id�d�k�JU1��#�Z����uZ���tpm��Ȋfe��X��wh$.Ii��2��y&�_*���亻�L�%��k��\
��IYF��������!���݂�3Ӫ�z��ޞ�d����)}��r�o��2��C�u�R +�ʹ\�_i�^��ư;޶ER=�y��q�YѨ�s�z�&�i�O$M?��ڸ%�կ.��A������8�m���z�wmF�K��K��ӷ3�gcz���n�9�gDy�4���%����y�rK�
����,�/{���s�ukxF��	%�5Jģ��f��K_�'(��HP32��8T���\�W���It=��"*�B�G2�x��x��d(��/]
��"r��Vg�4�c}�1s��js����(�������𻪆��jx++�������L3��d*-	��rS����X��uY|�AE�y�V�]]��A�xA&q��t�p/. ��2�U��B�PWkc.p���Ê��U�(�F;�WG��U��8	�K�	N�/JM�Jgk_�*�.n��M�T衮Zn>�s�U� � �(Q�+'Rv����I�c�jeS��@�3�u��Iڭ�Ժ���g?���-,]W5�t���ϭ������<�|y�.��<��nG�u~��;�Z
G��<{/�:rԉ�I�&���,�e ���?^�C��2�θ�w�wË��6�s��ϵ+�+�������	Z@���Mhٌ��������c>�J}�um�B�r,u�$P�]�<�л[҇��Vc|�/,����	�`}�9%��J��)���D�Q�(��FN�PF�a������BWg#�hy�>L]a�-��)�vANsu3���Wbk�u#
�����'2�^���p&�-�_
��P��J������ȠbFM�-��~L9�7�YNW�zC�mY�ą�Ԗ	0�[:���ҹv?��� ܰ�w�6[(
�\*�l�2����6��ޱr��ݰ��V�Z��?s=D~O��Yܛ��C'�.X9����-ye+L�hB[A���\J�3óL��C�I{��OVXV�lŌ+Ho�@%k��s
V���R�`�)Oߗ6]*]&'+�w��e0L�6|���SQS�.�*�^Aș��+<s� gP"�s�.'O5��-��^_��6�ɓw;*�9סM��d+}���~�>�wH�C�ҁ{�y}͙���:���i���)�u�U�MXل.m+Њ��2�E��6�AЗ�ban���l���,\jȯ�9K��5��]^/畍<�hs���qw;���|�b���.S��3�6�����Ѷ��I��~r�����я���7�Uҋ�Q�Bwŭ���*y1���a�_D@�T�#�!c��&�<S��w@���b���4�i=MH�N߇gܡKAHEQ��,,�HTez���N<D�C�qT�C�U��+�؃��Oy���,0���	ک�K�T�h�������YF�����g�0|����¹n���\�ya�M�����{(�FŤ����~:��wf~@�MK�5�V���ʨ:n�����$��ݜaDqQx㺚��������^�CI�+V��hM���e(�A]����B�Q����t�����T��)~А���QO�ހ_��	R��<������n�>[�̛roͥ��*�>�M�:������Z7��Yϝ��=V��V�h�) @�Ϸ6T;�=	�>�m��(ꪽ�xKk ��J�}`u�����[bVs�l���P���`���8�@��`�Y�7�v�j�uSoPmǩ��X����6���g�AGy�4�5��aܡ�+ۍ>G�Ȝxk������ZE/��8�$7��Z��z�
��د}���_��D�uju�`���g	��Y��������;r,����g��zD�L��V �\^�6�V8Oe���CC�|v�n���5�Oݺ7y�����x� 0~�v���������eh2ie�<��E'}�瞛�by�4�(J(��D����1t�5�V�n��֍��/��,J��2�D��6��g�>�}��o�,'�%�Vh	+8\�t�5��<u�D�7��!(j����d�7����>˥�pƮB[�1�G�P8bS��Ia�LS����I�&�q�5�y�%\��o��֞������s��C��ɡ}q�չ4\��9P׵���F\�*]qw��ue�5�5^�q��(�^���b��\!,>W�^���)c�u�{��NR�h敐.h��m�Qf���h~����Q �N��*V�Ux��o8?l5y�=��/})^{%ӱ?�n�<�[�4P�:�nw�R�ϴQ�X@\��~[{�����-��7w�Cw��_��{�S{P�+1:0�VT��-mD���
��E��w��Aɀ������_��M���c���k��=��P{|���/�z����n�|�����|'Wa���|nR|�P_��=w�s�x�,����眢\i��*�bUHQ&�Ҕ��9{��b�������U�X���m��A���D`=�_�80mI��g|-<�;y�g2����8ޫ�m�l�T2pɧ$c�݂�g~
�B%3*�{�{	�p_���c*���r��dn�Gim�N�b$��ِ��ݷw_���SVOz�Ϝ�S�dIS(��h+}7_�e�˵�od''�QI�֥��/'::���嘘�H�5��e�~⟫Lqt��(��߼-�e����?rG�l�sHj	�gq����q�C�D��rck	V� ~���@�Y�)��*��DR��}���xQ"*��4I���SS��b��5�OZ��DO�PL]�_�_���j�$�������(Jz��ϟx�?a��~dlOQ"�N2-��ό�/��#q���ն������7v�����z��cnn)V�L~�3_���çn�D���.�l����C୸|���7R"�S�!��q�o��nE+ vB�����ď�?�s~�,��٣՞�Z4i�P�5�(��V�S�ꇻ� <��s*�^7b���?+�}a Z���c��L~D;�y��LY��"ВG�0
�S�WP�U���?1?�DZ��yk�H+��{���ɘ�e�Q
5��
q'/�JJ�� Y�H�x����tT�S��2'@wV��^�}xd8FGFsMS*�֒��ȃ<��C�Ѐ���H#��|i��e�4S9�X��.���.*�g���(eVX�t*.∿�G<�7n;U��Q_{.��r�]u�6����:�kI�Wv�*��}I�]�不<����)`��֕_�����U�t�egsI;W�SW��=�1;و_��_�7ކ�6G�]�>��n�BNy�P �r�$��߻����wxt����cGqw|������z�{בT"�"Ɣ�Ũ�ֲCXH�P�V����13�W�;��>����ן��Ap�6=<0ˋ�ҐVE��� x3%b��E�lh�"��=���9�#�xocs5�E�=��mM@���Pt�4k��42���ݴ�T������̴��Ԋ)���s�3��Y�@������P~WWi~n>&&'c����`�֙���O�TI�-���'�(�*���q]�a2$/��i%.�A3�L^�m[E@���e���m��ܬ��K�,��#&-Z�6��ʩ���o�'�HW���ܾ�x�ېQ�*Ӱ�k�l�S�|��'M<��g�(�#N���%���@�B���Gމgu�(q˹��HT�5_a;LՍ��g�5��Ֆe���W���H�z%b����H]�LO�W����Ӂ�Nכ��7���Dw����T"kmc���u�@�7�n,-�q�-L����{�J���Q�HO���
��p[>t�x��O�/X"n鸉���s��K$���tg�~�u
،�g�_����w��".V�B`�����E�P!�aQ�~�Q>v�T?�}�mB���H��ah] �	%�7��`��f�/H���Bo������}o?9�=ZƱ3)�<g��rB	�52?�eE��r�a�l����](C� jES�� 
n�)+��O�t��ָ�,\W� �Z����5��0e�W�V�W�uk�;�>���c�����C(��y��c�Qh��!u���GZ@�CYj�ߍC��˹J�[�<��n}�ޝN��_�Y�S+����q�{פ�ah��%�.w&����uX�}�A�ع��ե�^�JL�!�pR�g\`�����Z"(	}ZR@n.T)���;qɊQ��hHװD��)�Q�S�`����������ߌ�έ�F�8�_�N;�G��������؂QᇄJ�������L��i�f5��������G�11���u��間 �+�a��2<x(��ݛ���5Q�2��S�j�g;1}��%��(Ɉ��t�rL���L�����#������f��@�W`߈�Nز�a-�����"��_���#�x�b0�gg�� ��I��i��Z-.����T�/����"J˥�;�$�s��jjg�Vy�Y�u�#l$@N�O|t�l�
�o�m�d�+ê�%o��g^U�U>U�f���e����z�p�̓4r����3]��4Lw����n, �=�1�k�,��m��v�����A��͝�*�Z�%�
�.�C�����W�2�J�����5|�נ������J�0�O��2�e���� o�C� ���Ů�K�SP�h6�Y�+rf�BQ�*	�>�Q���������U�p��-nd�˟ƁǶ�N���ϗ�ʮ��KŌ�\�.�4vCʲ�V�~��EhQ4��JN��I�D���3��>H<+@�VD~!^Phy��9�	�^{7��Ţ,2cg�ܾG������Ռ^��s2?qT&v�jFk�9Q,��Y�i���p�7�H<�!���#�����v�;<��*_)�n����V�)���
.�8i����<Oa�>ү�Aqn>�Q�B*������B������#�e������o.�ז�U*�T��fGY�"��E�T�Y�o
v
8���Eq(���ŧ�wN%%�In��-\�N��uW�v䴖U�<��k�)G>�}- ;ZK�i9Q6	��M�r��^��m��I895e��=�i�V��F�c�2)��Z$5�b�+>��L�w�HE!AU +ɳ�o߱�ڍ��2*�3�T��C�m@ Z�"�V�-G]��a��-=��y  D�4�/8Eގ/A�I\ t 8��x��QE�RP���x�K޻�/kp��7�:No���V2�Uy�ݽ��ou�Q��YHe�0K'�=S1��T+�]�o�*�k�Xf7߽Qx8��& ��l�n^���R(��+����=�N(��+���T��sy�r��Q��q���|��^\
���8�ǎO�����,ⵓG��ׁչ�#��!���f�Y�0���حDc���9V"ˀ�5�c�2�Bյ�L�p�2��_��!�M׸��L���PM���R~��N9��2}���H�|�Bj�3w���J��Z�׊��k�w�M����y�y[�*�21/�%���{�(���kP<��gpK+�k��W�N�& j�0�,W���ʚ�\_�w��Is��Tr�A8a���?�I��f�����}ixc�)���ޭ$w����� n�o�M���3AyN�y��~\�<X��q�T@�Ez('�ƜF߃��<�[����$�b���XG���zQ$�N@��vn^�A�>p�M/�!�zd� �25�o����ylk��97�D�������HP$C�G�k 9��H^{�a_���})����U
D����c��:ׇ�Dl�Z,J��GeH J����#$��J��O�}b�&����N��jV@sM�����_ȣ�p�Y0R/�Y>{�K9Kz%����Tg��<+�lC�S�6N��f@����7�M�*��[@ƺ�l�C%�]Mt��M�s�w!|�ε��Rh�ˮ��SA���|#��n
ES�
�f@y�&�
��o�s��M�x��5�\���蕊#�M�s�Y�*�r%}Wg�:�+�e\�f̸4�F+V����ū���������Ȏ%�ZNR�����u>(�T���&�R'�RQf��݇��a!d�t�A�w�-�	�M�j$#C0B�S���ɘ��Q��
�F�mL��l���w���
%���W����B�2Dv�Q����k:�
P���T��}B��,�r
i�t���w�9�\��o��W�wZ��<d���i���v�X�;"�y[f�� B�0��f�
�˔e��U9I[Ʋ^�����P�ʍ�Ӎ!��x���Z\�-h�䇛AZ�U?л����y����)�IU�J��ʚ""x$�+E
��VO_��}(�DpY�:h�Wca~#������^�o>�����K�b��Q�(�ݐ��W�v�r]r6nQv�[7$��S(�NRT�k���!G�J;U�D;�)p��3nˁ�bر�ڌ��p�:�X�{��f���I(^���zVhs1�$��=���]X�kD[#@�:�	�bɵja|B5towo4����;~���$�c,۰!\�PnY���ؼge*�2]�VxU��PI�������B�[���*;-�u�/����n�a�����v�����[�C�����|N4�d� �e�.枳VMKW��u`+|�p�)W@S�m9i	�A�E���ɚ�l���Hfk��L�i�7�
x�C ��Z�X���P�F�ҝS8o e4�:�MWWƑ�o*��A�]��er��aݻ�r

�ЍR��ک�v��r8��.�v�+' ��
6���q̍��ɩC����Jx�'��}�g7������'f��_���~�||��oǋ����f�#aIۖ��R�s7{�r��,�v*O��P	dt�uv�[�������esu9Z���}��C���W��RR��̚�d�<&�Vr�E�w�{~�.�YQ �K�M�\�'+
e�]p�h�:����T'�H,d���0O������ke�S�р�˫Y��^�nJ�2]Ϥ�2)x�4`za{����S���(�jE�V���u҂�����i(�S&�����v�G�ʇ��J!'���Vl�9i�I��e����	��B}�J+� ��bʞUK%�,��(�<�n�v�Z�z�M���:���sE�]�mW@�R�庄�=Zn~��f��/������
\^<���-��\�oC�A<d,��2���W�����í�X��x�[o�W��2
������ŷ��b���b�-Ѡw�А�ө8T")u�b��� G�W@�6�ț��TH(up�36�������7�Vcu�缞�Of�|7�@� ���Zj��R��^+� L3�(��W(��&H�$P
T��p�C�(C���Gё[!v�pH�P�	EIԊCa���>�%�Pݮ��٩�vth�Wf��RFy�1tw5iɜ(�Cz����BYY��[��x7��B�g�l�i=n��ŒV*�F��- 8�硧�)V��{�>.�Pʒ��r.�u�`�jy;NW	o� ��5�$�&�Vu�� ɮ���-���V���
{����5ͮ뼗��4j�<W����{��߳{����J ���*�+p����A�C���re)ff��~qy�:�jp�JYy�5I�ZC��G����(2�#oE��s�?
UF-צ�����打�s��O�y�G�jB�S�l��]A�B�̅Y���3A���JKQ��d\Z���ݲT����;����J-�v��A�'�gԊ��)xd6��i �?���O��Y����)m�����vC��6��|��5�B��SҦ��z��7�+�şr�;�n*��iqXV�HE��Qi��ey���Pʢ��E�ן�ќל��q��5ghR�a���s&
�=�)$��qn�r#(�U�n����w��<;��s#�8U
ݞ�1��&�==���L��A��z[�����]���s�.��oF�Q��U]�.��n�̿�H<�nĠ�%��)$�g��{ߗ7������u������@��#���v����855�%��C@Z����,�]g���`'����l�a��eN�M�`ՙ��2q�c���9���,ў�+(���ܤD���Δ��Z\4��[��#��xf�E��>x�Z����jE`\}����אqJxGG���q�ׂ�������R���m�Ҵj7������ ]&�a��D9
m�w�Mt���2Q���7 ��]�� ���0��>�wCgB�j"0^�c�_���@aW�k��?RQPֲ+�/x}}����띳
�!��Z�P��'��̋�J��#'�هh�B��5,����ox���6ܖ�m����\�A	݆^�I¯�LUJ#�~ ����'�4\�A�~��&&r������z%��߶�E3vN�s�*�=�j1��=3տ�Q�B�:��V!X���3����Jx�r�
:�]e28��}�u֪%&Q�j�(4Z�EV,��>��Z��*̺�>�u�(����SN��v�ۚ�zVC���C:	�OyV�aZ�{=d_B�g �%�?к��h��Ȋ��?�b�21�.e,`��q�ܼ�5�u}&�>g�ҝ�\=��+�&n����!t�������3O��يrH��aX=s4�)y���^����/� ��Q��9��9�����a��:/�VN�O�"�K�n1`w���w*�������{�r*�)fRdI9�����"_^"1���/���
�|����3��sE7�l+���/]~F�����������
L;eFi���Q��Dݤ� fB��@�l���,P�}�R����e�1>>���Ҵ���'Ӈ���
N��|tϚ��$��0>�E׶<��m���l>+P��u�������<�)�EA�o~�/�3� ���M��g��n]�A�1�f8��teR���S�^mTe*���B;�ut��y�sN�޾�a��0�tH�J�3qSaTg�������&�rcPHA�={�c���Z��)�H`^�s�6�O�I�,�rgc��FV,�2�E��Q��mP� 3����;��k�<w,[X�E&˒�u�x�&��Ű(IP:���/�Z�<��	�IKBZ ��az ��n�����[7��g�9	��\�mV����0��y��fh"�ٸ�<9���{���L,��n��� �SX�<W��yU�΂JB���NA��4m�Ķ(���v;�ʖ�ݝn+�K��`2�̽ȝH�1 û���{nI�v�坶4�53yӾliXme��$r�^�L4�˥uk'�a%����� a�S���M�״�a���9��S�Y�b�"���o�ȭ�|��XoM(^��i̳�_��m��^z��y�;-�&�ε�������J���7�Qg��p�lm�M��يu�qņ�z۔Iy�v�oQ������«I� 84�Հ~]v�R��Ap�����9+z�7�w��it����-��,w�Va��9D���-�kG�@^w6�I7�!�Ƶ�U7=�]!����Q�^e��F��6�܆p��喆���V�m��&�[4�n��J�0-A"�2�I9�_�9�#'���h(�*N�'���*�O�	�$����=G��˦���N��V��˸�F' L3N*�|;�J+q�c]�r5?`���Jޔq��vR u�* ��$&�Bi1�}���)d!<����/1�{���E�YM_p�WK��=�z��Ē�R�`D����!�v�պeqգ��6�穀�b�*P*���o}�
�RM竸*��&������E��� �I|ȫ�@TXŵ�xed�V=G?T(�b���XO=�O"S�U�r�G9je�"0n����E٥2�Q�
Tt(�Fw����[���Ze�[�g���nZ]Uv=(cq�*�*J���i"�QiP�N7�F��v��uP�N���/�\�T��I�q�����4�i�s�k�&��k����I�-�ۄ���K�ZC`��H~���57U����[�,6p��4�>�&�o
�dæE�Y��k=7����4tz���I9�����Vc��P��PP�����W�V?Ŭ��Jd������`#����"Y�?eVT扠<�a/C#�F�>��N[���C(��G�ϡ�i���bbZe���0Ja �NSu��V�Dw�%[�ڋ��7�Pv�x��Z�3+o��p!p�4LHK���:QpX=h�.��%�n4v�D���/;8;u�4�6	��nt j|�h���4;UVe���c�Q^�N*"�4K�X��*Ui؇P�֎G?�l���ơ:��� p�W7q�4�oK��� �#��n]Ɠ�`� ���F� �e����U �ll�rBQ�o�������ozﻰ�Vy�Ƶ���(6�L�����'2�nW%��m���[=�'�Z$�pS�Q �O��W)��j�snj1  ��K<��s�	>ۚ�e^X�n��&^�׀��g��e� �#�ע�� R�.���"Z��nh[팵xq+:�G�:�Z�o����K'�݄56	]�w��8mK�0ٵ/���y�5O:k����M��W��by"b��F�_Z��(�֦Q���<�_(�9C�$Jc��/��g�cy
b.a!u�P�}(��>���ʓ�fM��S�R�*EaU���~)��@���u*�28�xʝ��0�R�ݰF�����%Le��8*���v6󇸠e�7;A�{�{+�]������>�Tn��F���:�W���T���b�E�Τ��z�i���:�ף山���]&Lʢ�iע�_o�얊�LO�l!��{��~�Ѹ��q�P�&�����X�X�5�4 �N)�l�Z���-q�rcf𐜰8�+�9B�B��F&ߧ��ׄ*�3�U)�rÕ
�T3��(IL�2�U�(��B��f��Jex'�~��}6�#?�J�J��+Y�;��������<��\��/����壚al�^�c�g�W����g�'c��+<������L������lh���lQM��B�n�(e�Ѡv@o��# ��R7kN��[v�N�07o���້�O���0߮�de��٠�7e���ʎp�D��V:���e���]�6Pn��c��@��u�V�=�|-�B�9te��_r��y��=<2����b��@|�w���o'fQ�kX��R�{���>"�)�P[Ң4���R��̊nƷܾf�K,[���Vq�ȉ�ԇo����0}Ey5G�l��$I�G�ȳ���2�V�3�z�\*����w����I|[*��W��c-�N^ŪDp�ų��|~�(S�?-?ȩ$��^�װ,�(�[Z�ϬE�@_*7�u�j���˳1���'?gn��S�7���K�󹃚&�g+C��.�TL��T�����JZ-4K\Q;) ��)a��D	.�r��beY�)�yM��∅a.b���+�~*�����kz%R#�Z1��򞧅����W- ���;�ub�̡�8Y��։��et�U�x��E�Eׯ�Mi�*�Z"*�eַ.�3�ԩ÷
����E_��fO3�f璄
���J,.-f�[__ne!FG�rn���"����v�K�z�L��x`�M��bI����u��+�n��yJ��E�&
�-�n�&]3b\�V>p�ui��l�8D��cG�ġv?<����v����)JllAo�.���s��	=�M��/�^�������|7��f�Ի��";<�yB�&a��P�s*�@+�|+���|�׮
��峂�66�7~����g~���c��QQ��$����� A�K-5��o��N\�Z�O���7���X� ��Z"]�11U���@�Wm�k�AF�i�s=��e+d���l��
B�D�D�GrG��h2�V80�J�޻���$q'ci�i�*Lc�6}���e���`2��&�$4��O����2���|g\��r�W�"�+���VV��e+�V��Qe�L��ΫL[���k{��}~A|��>���,���`'������B�2i�Ւ�ⰏF%b�2��E*3ʐ_5#̏����D�߹X��R�VӲ���m˻0��ԓ��z��Q�De��w����;ʩܑ�����̲`"�/,���T��C��q��;��'N��˗���s���*qƬ
�ʕɤ��~��ոzu2;DW�Hj�������C|�&?�fca���5aAjU:���`[\�F�m���,�u�`O�J{��P�TXg*����u��ux0�Z)���Ӗ��Ď��ٸ<1�X��@���WuQ����^�B�R(��|�.��8�\� k"��]ֿծ��C~��>��3�ÇG���rX��m%���m�)���<�̛15����3�����C�M�Jd�*��%�k[�)T�H�
A�P�3*]���6\��	\��U�	��D`�AM%B�R99t� ����]���� Dl��6����31	؛O��DVb������}����D�Մq���$�+2�B��VZl�+�a-�S��@��U ��;�
��������N���*�X!�qj��&#+�2W
����è2�������m�:�"���&e�|zb��Ym�{�+�/�w4�7]G$����ߍ����D��
++���;
�ߚ�Qi,�����(S#��F�WZ�v���Bˡ��r�A�6��/GQH��o.+�������QX�Y����$
Fˤ=fg�)���A~�º�g�WwOw,o,K���������f�:�~%\��,ŃwlT��ft1��=i�c��{�oD=d<��2g��(���g�L�@Qc�Բ�k���n{4�Z�+�a"�[H��ꄮ[(<;�M?1柔)ְ��%R���s
�J$;��H�t��#�<k��u�\9k�|������cq��x*��gӔ��K�D,0�
�@�͸|�\��lv����ܙoSQ��0�+�ڷVQ03X��%#8�
��8((YqT�ڎ�� ��F�2}�RNp���Mk�5����X�'[B���il�/����qߝG����p�i�_�t1.]�0��"pk��+('�XiV�0L;62���UHv[M��/Q@
C�dH+b��i��b,+��&s��T`XG͞={s����w�FOw3gReI|�/d-FG����ño��x��x��ߋ*q=��y2x������o�y"���OS�GG\�E�*�2cQ*ߪ�Bz@w]1�ɖϣBu�QphA=|�ma}�F���Q���6/�Sp������pq�Ph](�8*g���`BOӮ��GΖFH:�^�Ō�������O8�)X��4�(C��W�����ߣ�yZ!<�-�SM׌KX
</��L��Pmf�&�yk16�
;4rI��[����M�4����x�y��mM�Z���g��\��ԉ.��X4d}�X�'�0A�������������{���M'i���T(jE� ��~7��[o�o��{��}�y,�'�;�P����Q�1CK�g!����<f�&
be��Kf�`
�.1\[����褥��|&�_��*/�u���c&/�|+����½Z������>,���+q���l%ռ�JJ��݄�K0���3��ƚ8�2dmjʸ�����y\k^{8�[��weD+���[-�0װ��!ɞpY��7^�933�i�[���s���q��x����/}���s�D[s(h����@aT v�,�*� 1�R9�y�����⑖J%���x�C��ʲ�i����p����[��Dĩ�.�ê�e
r���c7��Q��?��;�_��g���?���-�K��U��;�����5�P~Խ-~�
��*��:cT�
���C�MXr$�}��Q�<��,۵0o|��F��3-p�3��ɯ��`�J�(�6\+���a�E��6
&���wZD�XU�o���;�o�Tܺk��Kȝ�R4_H�K%zR+	 �Xv��ֈ���G$S��|Wq�,�Y�C�}O�
�Z����{����)>���L��D鵷��%��e_B��7��QS�����Vc���+)�~��8� ��|�~��@3��3�۠Br����f����f[|���G�'n��@��wRi3~.�G�q�1~�@L����ϿFzmZ4�]�N\��}���sY|l�i-
�9��N�S�:*�$��}7�	�g�d�h�v��+D�Sy�N��e>��!֏|�un��®g
;'�̋)3A��a��`[T��i���AA�vP?e��u�uV�1�h���$3�6B	$�9ê8f��D��Ƀ����h��Q�Ŋ!�-88�ΙvE���d���u��z��/�.�� K�Ơ��)��
��(��ӣ��3q<�>�a�Oߵ�u�<�@������^���{�My�s�P��@Q�uf�Bo]2,q��g�fHd��̹%RУ~/;s�4�Y�o'��qJ�N2������z?\P�V��U�NR���G?�|�wY�L��S�[��N��0;���d�wC:Y�w]� �̿�����Vo?��ӳq���8x�`<����>��z(���[n?�y������bfa9���3qab.}CX��r���A<[��r�]�д���J �Jǌ_Չ����4ߕ���*
��Y��W�~�4����&�[��3�tK�R�J[�ciW��UH�&a�~P*��E��y6�gu��%n�d�ӃV\��h
����=@2�,�l���pM}��x����~bq-��U��'��0����Y*���>�?-H{��_�V]�K9M�"�k����
��0����/�ߝ�j��m�߱�"���RĔ�'3�q윔)m%j3�>
�y��I+�*GnAM�.DQ E�gEq�Ff��x��$"���>Zl9b�>���	q<on�|d�N*y9[%�}n����*`\�hVQ +k�<_�g!�T�M [�TTM��~κ���2�\ʽ�Nr�������/�a�s�R���[���������8}��1�[��'���߸�}P[���ȅ����NV`��ʺ�S�T׻�7�[��,X@�*T�����b�����$���8�|F���
�����E9��E�E�z<o+�p(_����W����i���`iQpm��x��/�5u�kme�A\2��P�� ��>�~Wٶ��s��.�v�������e�ۧ:�Bk�[C�X6~�sQ�dk�E֠G6 ���{��#��QҶ���|�PXݢ�D��(/y��	����H��)��R2+ĭ��E�Ng[2Mg����X��/ci���ǁ�G����==~�ݡ7�u�C��Ž�)�Fg��7=�.�R1�~*�d��̳T0�L�x���
��`d�����$.NJ�n�ų�};�����w&cy����j+�{�{�/|=^x��h��fk��L\�p4IS��Z����lUJ�d�HA.��8* ����3q%u3 �R_Iκ��b�{�^�#p:xQ��e�
L�Lڪ �
�;PJE�1��/�Aқ���p��獌����J/�9��䗴3m�%��3��X!�]�_�{˨���;q��(K��x'����ƫ�\GV�[;;��N�r�AB�v�
�\l�u*xyB ��>S����\ޫh����(���I��<��e���(�,�%���-�eM��?ᳺRJI�}�6�y!�n��J%/���*�H��?�rQ��C��.�ko��s�<���SW��6�8��Tɴ�S��+a0�a�͘�Uj����(�wC���i�¨(�_�)q���3�8���:{��3/_��?�j<�¹x��7��b|�O�k�_"����?��0(�-GrH�:QAZ�$i9�"�>�p����͸F���a(@:�̓P�4�����&�形�K����Vi�3���Ee;��}���]WRp��,�,i���,�=���-���PZ��m�Q 9�2�<T	�с������J<�@�"�x�MZ��)��%����յ�#^t��[s�p���.�����I?ix]?�HŊu&����Z�vS8�`����ǣwR*��0]�*%
�f⬠�߷/��;�m�7�qzd� ��%.%Mo�{)�}�4�q|�x�ɃXT��NL�
S�u=.\���LP�
J�e�p��VA�K���j�d����h� �d�
��$\K؛@�|�0�	�s���oO޺T�p���~�H���F���D����8wa������֌�6�����Vb�\��D�ZEy� {N�iI��>�xY�"�E�t�ʵϴ������c�Ul�2�S:Kk�>;��Z�i�y�u�Q^�62�a>"�҈��-C��>'4�Υn<��;��Qx�tdv�>B�M\�����~[k���h�6��|F8��Qn1*�f�l,͇�3O~�h	��2@��"d�w��ڰ5�3�BX�C���N�o �l�a��V��w3�m�:Z��s��J߉t�ޫ�Ώ�svҡ���D<������u�Ue����X�l�:G������;}� ���Uhj��u>�������0�B�6�4�s9�A�%�D���&�J�_����[�W�%��<\G�C�1����S0Ԍw��R�k~c(����U�DB
J��y�%��p��olv��y�G�������
į�'��~���T�G���&�yT�e=l�E>H������YAHӛX���H
=M|����R1��*]9�{pp8'�%_��x�Wp�_|s)�CU�2pn�C��z�ߵr,�����*�,W]N��HΩ��SnF%�x�� W����\F ����̫>Wt����p��
���m�ꁯ��-,��k��sۙ�Od�F߻a�CŃ��௾25q&Mi-a�3B�z	�.q��3�>�}�<˷}]bJ����8{�l�rX���DGhu�9T��6D��	�D���n�V#��/��h��~$s���0�`%�
�D�<KĪ�r������̀?�����x>--�&# �YdF��7Jj&Ľ[�h������6_K��?�(/�A��ݐ���վ��&�
X��id?��`k3m��{l�)�E�_"]a�݂�pn��lx�����Ta���lq�=!-!�&e|𹝬�<��֊z����!�䑢!�U�"ni�܄;gt�S[�"Ĺ�n�~r&e}�}}�YԜ��gn[ݔAp�o7����KWwg���v���'�h�&�n�$/��v�9)���$��S�S���,bܗ��<P�����
���&��뒑z�/Aky͌�S�� ����2k}T���yݎS��bV���Z������(��Q��4=��"7��?g.�-�k��3��9��KEiXڌ��QX�2�:\��;�/e(�uqj�T��'T�3 �|f��r��m��a�Y�E�R�8�L��PҼ����F �6W �*��֞b���r�c�V�!���������s��B_q���s	/�!�D(���o�nE���N�Q�`�����^���\λ�M�!q�,��{�`˧�0�2�(Ö�ͦ��
8�~��7��t�L(7�!^��õg�B�B�jg��ayc%V6Wt�+E��	8�������xE~*��b��Xj���G��C���M���S�E�C5Pp�PQ��r��7���(�^ht��ϏiWrTC��|����y6�N�:�>�Q�� �+���T����P�*��z6�q��(H�v�e�\LA�12�L��2�a*�Zqԅ޹.9 �UR��"����{�}��ך��|��(d��N�j|�  ��IDAT��{_��s��d��nyn)�oI���������nvP"����N��
�r��(ė��fx�8iYK��6��f���2�4حl���a7�Z�r�����M>����+@�=n>��K��5[z?x�lf���׊������E����~�¢R�ܔ_�IbИ$�z����£�!���{��;�h�k;x)$m|w�s?�k����h_&�A�XCV���J;:�$��t}B�vm~h�J����b��D�r @�3j�^�|��v7** �ká]GyT'��cw^�������8��Q-ˢ$R�s6���Q�
8d:k�K����=V�h5S2U��̵͈Z�3�����!f�=����6��tJZ�n��_ċ7�x�4�2+��n�%[D߮c�k��O�F��7�,7�4yH;DNP��\���Lg����j�%�܍"q�n�E�g�n�-u��t�\Cu��^����e�	d�U��&�(x���P�$g?�KÑ��t���^+�Zٺ<�����������[i��+~�u��{K��e�O*�T$�[ʎ%boX��rt�F�2n�قzH��ptc�t��E��Z�>x��jF/�Y��۬� ˺��1�*��>�]�ZK�I���xR�L:��5�o���śBǦ�/���-�����fIܶ�{�f�����a)S x�����Z��V4Qa�L���дQ�ԃ�|�Z�0��3V�Pq#�d."��%0f�(�g;'�,�U��~����Nz�z'm�8mk@�+��n�e�9|W�!�$�j�.�g��[���%���� L<��2Ϻׁ�]�^�����c���מ�ܢq��61c���!����>�$?iW�P+��P�������O�Z!m^[N�Bi�\+�>��M��riF��|U�7	_[�K�2,���������5Y��X��O}�VP��* �r���#@�f�D�{VV�A@ ��?
=ƨ����F/��8��`�{��s7-(�@�Q]ד�zʹ0�����;Mꨏp�Iu�w;�
�m��[�)�t��ѱ���K��X#��ڣ���^���b*,-�C��+��G�S�ڝ�u�r�u��S�c_���, ���d���+����?�F���ZL,�?v�`����Ƃ_݂)\��T��ڂ���ʅ�� �N�d}%��
,�乷�{��,��Ӣ���Nkܗ�j�*��jb6�ĕ�c}n�p�Q��,F������@NLCup��h���&=[�􃫣fnѕX�#i�d|�R	�Bj{E�LJs��
-�3'uI��>���;GY`H�]���"?}�-��-�&�-��e��l�ܘ���H.8v��f�Mm!::��m��jv��:��J���5�(+��T��e�Q���Yn÷8�%���nZu 
���QPH�2��8��]����bph_B��� �T��t���;�A�a���>,�%����+;�w�5�Ni���¡��q���\�v�~�t���乂��N�sV�eSx���B�Riݩ( <q����^W�.��O=��y.�zcy)s���{i]`�U�g<8���KwH�/O��*�5hశ�ol�r�Ąɲƅ���Жw�k��G������ފ���m�pF��ԎX�W�+�R�
t�]q��73P*;i�Q�� ����M��+�F=�W��8����OE/�������Aҥy��e�A��0�03y%�{���T�|���7�~<�y��C#S)]@���:W�N��f[���`����JF�����<�z��D���۽���D����R��Cr��C�;ܥ�+֧/���T�/����Mp�V�`�Ų{�@\�|��f�*-��\�t���������_�]at9�SFe@IԵ	��TX��*4Sٵ�w��PYAz�l�i���MWזiU�<;������Y�&y��D땰vn�G"3�9���\��ݠ�j�=0�������0�NP���g��a0��r��8�C�CI�����A6[�BQ
sAd�5��<�brF�;{����]]E���C�n�ؾ��N�u����k���g���A'�F[w{��*�:�^�����u�_�&��V��D�߻5w����=�Й;�����0�C��I�m�{j�L�qi�~�Bm�|�щ8��l�������W����3�u���?]*ёP,TT��,��P#z�t|����{s�vY��'�vx��'�\^���W����V��YN� /�[\��X�J�;�zs��3�������[_x&f�{b��[S��9t�%�a����J�&m��ʕ:�N�~�'T"�5���?y�}gz�ޘ�å�Ƣ�:s �Ɵ���h_uo�D&���lȣ�JHu8_Asw���x�W �@|��7�?|�;11��xc��}X%}�t��D�#hY5�m�l��b�&�t��Bt`%�6�y��E�('�@k04<J+���2��N	�;M.[4�[rm�R��NA�b��؍�����`.]�lp�����i�8[0�>��~*I_��;>�Jfff*[%;����4���)ݡ�Aنz��*:c~i%.NL�w_��Lt��SY��S�$R��t�+��n.DO���qd�x��� �nD���싉��X\^�=�Ƣ��'&��Uw�o�SXh�����}���;+�:5�s��g/���F#���0L�:\�� �@���Ŝ����b�d\�m�NK'Z��	S!*���)|���l��R/w�G���s�h t�O`�<U���э�*���S�� ��*��&
FkK&�gځ[������ǣ����Rqfg-V���ؤ�t���Zq2���*糨(�\��s6����:�0j�}�w�(������;�&b��]�T�(V��t���k�Q�����O%����@� �'Ό�GC��Ӏ*D^��Fy����_v\������]��*Ô�e�"�M@��џ/~��_��~%./Sw4����T�l*��	i�%ѵ�NX���*Bkح�K��uJ�i�ڈ5q�Z-��L7�j�;O������n������!�x��&Y҅�U"�ĶE��q�����oD�5�x����y"�O��Vg-�`c�,!�K���mk�X)�!)��پ��-MNU g��1>Њ��bL�}=MޕdL
���=V��`o;�#���ˤ���C%\9[0�K��N7��pg�ga��8y�p<�����x��Wcnj2{��:̕����(�j%3������ϡ8fc��ju�0���&,+~F��~#>��_��%��.L��L�O	*[�Υ��G�;�ч����h�0�O+N]��~]126�0,C�E�K�h�g��h����TK�f_��p,,a����ZZo��F�֗�_���B��aF�C���U"��8��%��ew�z��̞�O)����4!=}���]8��lb��x�+����a�0�����G�
�[Q��íܓ֦�Z�EҌ��@�:{:r����������?�C1��o�W�~�RLNO�p�7x�4l�m��p��Eȭ]f;�.�^�U�ׅZ^Z��������8w�r<�GO����N�_F��6��C�� �윍%x���~,x�J0�VOy�h�i���Ce�ž��EC�D#܊����y���e����6O9{��bl�?�����_�7�k\Z�b�:�B�ʬf���K�����QP�A�r��Ꭸ�h�;��w �Q�X�������ʏ�D�s�/"�O+<�o嘄:D�z�D��/�;����������V\���|�e����r�棗��D!h�9k0�g[��-�VE�n�~S&���N,) ���$�p�10<K�d�0���Pe(�:)� ֏}"�&��&/�u�K����࣎�_��O�ݧO�/�1>%��^|�6*i�W�,�N%��ߴCY%�߇�A�(��h��a�9��H\������'��o<=�#�'�Hl�����.�Zم���� ���}"��7cui��]w���a��Ų��S�׀��Ҿ�����-k+�I��:P�-�e��/|5~�_��e���e�M��`����@3_��z�����j�>�":�j��ϥ�S��f���ީ���.3X^$�]M����G67��ڭE_�#���v�eA�`�ٹEp�?�l_�����P��6W�S?���O~$?@�����?�����Ob�ʋ��zs�[+z��Y�e��t��dx�$�E�a�e���M��\��j���*�@Ύ�8�4޴���	6B�?H�ؠQ`v�:��F��3��2U�ظ���L�������j\�Gu�õeޡ���������=z_�3�?�x�����D�ݚQ�R"�r^�$�ۖ4�ɕ*�]�⌂����MZ����A.uQ�k?��'*%B|�1O�`!����������bːj��쥙x�s�/d�?l"~�N��0�J����AFSw�q�L�B�9d��s�z�+�}U��S���LOѳ��/K>9�F�؍�\[��5��B8̡�} �4]���~Z��ハ=}��˴�-�w`6+�T�SmX1����WeՃ�l��'W��Dr�5\)��M�UD�I�Fna��ko�7i���Ҭ`��G�\l�@��~M𘝝 �������QG:���K��Ǣ��'���m?ܝ����uclZW�)�ه��uD�ޡ��F �ںh���|<��s���(*p@!:��9ف��RGB��m���VVu|��Յt=�Q��<[G	o��ɳ�V[|��}g���\���K���.�[������Ĺ�Z��;�}����4>������?�O�<|�8}�x����_~���[Wbey�:��O��kmB��n;�����VP4�����}���}ii���bn�]��������X֋���S����v��zX �*��]Xk���J��.����>B��*g�_�<V���Ū����͠��	p�:[�*]\��)�<��2��̃��
��:ro�=#Cq��bt�o��Z|�b�/g3#����O�l�`�تX� AcW�;��xVN��F�4Hd�ᾎ����8~`8�Aa��U�4eW%�;cB��nT���g��J�y����jWM\�\`\?�d��{��hb���8?nnt���Q>]�d��T�xc݈<�����^\*Ʊ��ل=Th��iv&��
ff_�������e��ܳw_�y��q��'��=���팿������T�����jL̮���,n�����WgV���2q7br~=.M.��+s1K���BLϭ��S�=��3�9J뾔���;ro�8[	���PsXe�q���8q2��W�����pi!^}�|<��+�o|;�y�54|g\�X�'��^|��_{���֓��w�{6�y���淟�g^x=^y�^To���uq��\|��O��n�ꦿ��� ܺC0�F���Cu�ٕ�E[\�<�7PX�+K���AIl��4��C���?z�}�27O?�-��`�Ȭ�請Ѷ6w�v4�"��q��|8F{cl�/�I%��芧����F�lt@�z���).P�3��ƭ'F/<��0���?�+S���N��瞤𒝨9�o8�Q��y�CUs��$��i�),�m�<m�h��Ф[ǻ�i��f�i�����'$or��T>tF���B�Z
-��0�:��>;+�q1�,hAu\.;���������C}���S�o<���8�� �: �A��Y��({V�h�x��Y`"i0�ˎI���tMiD�CN��a��D��[穀H�^m�sȸ��Fu�.�0`A4@��x�t<��;��رj�H�$:1Ea�%����L�EZ���Ac�����K�S�n��ř8�$�zb~�
-�b~ k��4�h��������������� ;2<�}�-�M��������vGM�z���q���{�sO�?G�Ş���Ѹt�j���f����%��"̾�٨ce���*+�Ң��vBj޺�{��uQ�LU70:{��?���-�;xK�)abHB��Nk�OT�a}4`�Aޑ��¤��\���a�o�̈́�V���O�89*��`���������'��^[�����/�?�����s�A�]����>���V�xZ��e$�:��&G�t���w�r����!� �[��V����g��o3������>��0��:>������=��z~i.�'���x����������k�<l�-ڤ^�P�{F���/~!>��{�Ss������y�{���֗vLg<*�5��{��a^G�VP5�稛G���Gh�Q�CA����4rB���-�V��!�t���}<Sie�v���@6�сi/�BU,u�[t��u��EW�PZ��k�~df=>��������x�g�����87�u��(O�(H�4��j۝��m���U
_����J��s���s�i,a��-�z�?�X|�}�c����JtK,��%"A-�K�EH柚�F������x����HD�b	���Q����F��1���(3��Ko_�����x�����a����x�������ӷ�]�ʲ�5;ۨ�Z�сV�v�@��v���f9�+�|���	Z������8r�0V̉9���C7b��=q�ء����]��s/����~9^y�||���xx���8w�r\�8�p�{��q��T���E�\�����,qΣ��x������I���C�0�f��'?e�Nk���=��0JW�۱`�凉�����5���vPc�L\����U\WR.�N�O6�2n��(~�A�E���{�8e�������bL��fwS~�$�����A6�����:o����r��=�� <6�=�i��%���#0�\����;7O�zp/(/���4?����s?��LQ������o������c��9/�Ol|��_��+��O�nn
`n� �-��G�;n�W�籄B���?/^��C�*��gJS���gX��`�7��X��;����K��=����n�C\��!�-b�t�(S'¹���s��Ѵ�W�O�n�/g���u��$r�Tw�����QUl��gA�Q�H���í�U��Z�[�k,ʯ�u��H�{שi���_���A��s�Fť���,��K�ܳu@��T�Q-iY�ʝg�x����� ]����J�k�{N��#��n.A�����Ρ���m�Q���Qm�&��2��Z�yyA�A]���H�^,C���),����'>���b<|��q���q���{��'~$��_���˿��qs���0�CV�}��������ſ��k�r'nNw�yg�o��ߍ������=�o�ވ�_x:�����>k���=����E�Z�Y���S�}��^*��k�m�k��@ss):��gk�gK�-?�__��K�}���V��+
�;�hC�۹Z��=�10h�4��G��N�m��,R�~f1e��%^O�	g�*���׌ɩ��E��
ŵ�8kˋ��VO2S����/�1V�S<W�֯q贾�B�X�u�}X�v0R�T 
�.�֛��]U��;s{�����ܫ�������ܗ�_}����o>��� �H[EG�\ćr��]�LnX%X(�Y�FZ�-�9-#�(�7���Ź����؊�>�� �ͭtZ�����Z����Ҋ�uYE�}��C�tX>��������@���^,N�����Sq��a�I�����ᖷ�Fu�߂���VW���+�W������k1з����:?����O}�#�w�'�`ų��L]�VJ�����Ŋ{���y�uŀ��YeQ�.(N��7�&(3���E}p/��LK�j^��"�Ԍ�x1�~ww��B�13�O��d.�IP��M8���*D�=��?������T�<�?�H���������i4cϞ���������!��H�2i��{�����{�䃰ݴ��鏾�|v����J%29y	8_�Xb-Ǵ)ݎ����Q�E�h1���:�aZF�E+ڽ���A��l=*��ѾH�`8�+KWci�2:�*&�$�<W �������ul�- p0/�� bc&���Z��nah`]��C��T��3Py!X�>܆�.��a���7��r�ln!�Dƌv�`U?�zr����v�Ƽli�5Ҙ�Ȗ��\7'GbbEWl��]â���K��((c���0�^���2]�hk��C]����I����N<�������V<��������}d�O��b���:�9�2��8=�k ���������� �J˯�}i�\��B�,a�R/m��\)�S��s�_��t�����H�4�sGƆ���O~�c��~0z�Z��6㶣��V_/M��O΢;�ؔ�S�~X!ϕI�t=x���3��B�G����������=�݉�� �p��j��sa��ݙ�y@��.���G�NEB�$�q<W�d��\��������2Gqww�������*��%5�Û�˞5�sY7&O��P�$�i6�qj�U�xc����ӷ���䏢��'y��o=��������R����_��_���v�vĝ��B�o���-�PN?��o~�=y졸�Γ��<+3Wb��3�vwtAov �-�&_��BXa��4=q5.�}+�2�C����i�N�6hI{6c���/� ��H-JB�>�͕l�=C]��ݱg��hU6�<3�tÐ@ShTgW?�4PV]�d-xa�E�u�-c6��M]wl���2�,�Ea��6��9�Fo��f�ŝ��T$J���d<�#������Ŀn��c!⧷9ö��5��31�]�$2'Hg��޾��nP��XD���م�4� L=5������lE��������Xi���=������bt�>�|h�޹p)�y�9\¹�ԗ-ms �Z#��n�����v�tw�ՙٸB^~�}�~0Z��f�s[����Cq��@:0#�Q�~cl��'�8��?����Q�oh��+��Ƣs%فe�D{�:"�5,]�t�w��'~��~��qϝ��b�g_M'
p��?��pxp���<zcߞ�8|h4cY�?0C#Ф���B�"��/H���ǱC��2Ң�՛��(<dz�<��"�.n+e^�Cɡd=T*���t�CeA�Jiw'~�\Jz�,Ӵ�P|t�T,�����}�N+��B�,����4���u�՝se>��Q�MfMK�t����Ѐ�za�>��[����p���K����%^z�Z����<��?�~���9�ҮX����|⭮x���1g�bt�h<���ot ��׋/<�?����(�lp-���$V�D�-�6�>��IWian&k��{cx�	��� ��q����9N�YO+��������OU=�gV�8���~�7覅ف��a`��V�j�4�1U�{zb���v����'vB�0R7Q�.�45�qZ���8�	�н����7��އ��8x�VLOL� ̫X	���5�Ǌk�F/����[��|�z	�����.S���Q���G{_�~�R� ]�]�	�h��� φ�e�bl�p<�������"V�W�VLbIt�E[/u6:�XO��R��t5f��ϳ6��ƭ���P����e�@�T S�115��-���]w��}�%�w�#�����3��}��E{�6@�6Q�(�ۏ�S?���X��K��ʺz�J������Z|�?����۱R�i|�k�穷����/>��GP C��P���(����p�������wh<��&?z��>��s���/<�ԛV�V�ni�= �JY��͎2��>R��ע�n�JN�ܦ�^��%��@6�X�JCCA(y�Tv��9��4*���⻫����Z��*��D��t]Ҽ�"�D`:{�<��3o�U�p�� �ͯ��x���cߑ�1�:���并�<���m�OT(H�-�~��w�x'��ē1M�e����,����D��e�^c-�Ɲ����������X�zBy4���w�h��vaFR�V� v����K�ҏ2h!�(�z`�'N�~,}n�w��;+��K173�Cn��l���,Ά���MZ�M���rY��nL�^I7
�\�����q�ɻ�?���q�cq �p+� ½A:26������x/��/��O�_�����h[ԃ.��v)?w9==��նP����B(l�j
N��b�B!�<�~��:�}�g8օ�0a#�	�������g6����c�1���jc�2:g�}��x,�������+��XB&P�o\��)Λ��ꍍ�X6�^�����R�9����?�(�����܇�����,����X��6܇V�*�݁�5���Vg�}	��?�z�}(������ȣ� vK�GK~__Y��_y9~��~/>��/�����NDs(���+(�坷߆����k������-�%i��b�����q���8p�@�sϽ1�r~�����_7��{`?|�i�Z'�8c@S>���\���-�m�.��V	�q�]���Q�5E��ʽ�6���?��T"*����βE+�G��ZVwR*�ȠÅVX ���E�]�˱9�W�cnbE����p���]G�0���7�ɕ��4�iRc����	��| ���KS���>��k��mGc`�+V�m%�Q"��_@���b���a^b^w�
�Cv�Qv��������������T������%N;G�ӷ���>�H�����5N?��Ci�s�Q��_Z��v�r�g�
����/bǤ#8ˤ��������3w�{|(y�#qי3q�ԉ8u˱8|do���P�����h0N��=���8q�4.I���{c���}�����4�ac�3��(?�G��
����nV,"g �ﬡ�W��.�\缺֞����^���7}Tf�l��%���@#�6"6&�}���Ú�qr�TW{�g��@��ܻ�����NUp� 7n8Ï��@�Cخ�UDg�⭷/bY��]wݏUv8g,��b���:�7���P<p�#q����C����'hT�G��@�~ۙ�29_�ڗh����f4�f��m�v3f�����:��G�Ǔ��~��[���h��Kq��;��+߅Fmq������;�S���;I��-�Ǒ=�be�h���KC�o�A�}�e��P�c�(K�WA|� ȩXbS�s���R�(�*���R	E�\�[�����{�+���`G�h�p��<��q�D����eTid�f�鑣M��ٹ�Z	A0���i�>w���e�*^�_�ߌ-���uwD��B�F,������F���~4|�^�r�l�����p
�x-^~�혤��$�u�݂�+[����g��߉���x��ȁ^;��� cc���)�3�
����`J�A/#E�3�?�ǎ��1Z�����<��9kX����bm܎!�����8~���(�[���{��4 
���¥��1���ͽwݝ��}%Z��'����<G�����"=z��Ĝ�s���4:�'�?�O�c�XG�����}�b{�b�~�����x�oS.�(Z')u7��D�Z�־m��R��ve*P��pۼ���Q�@������yg[�Lh~X][M�����u�G��^ĺj���
�ӱ]�̦3?aJF,0��*�jg�8{M���p���3�Q�
�C���s�L��0(6��<�.�����/���g`$�^���ߺ#�P��qw��݃�����q�#~�'�b��{q;��H��q�b8f�l�w_y'�~�%\�Ix�ָ���q�c��]����q^9��?4�BjR�UEx�N�>p"�{�x<����?��+4zs�5p0zGa�R��㮓�ǽ����CXs�ӏf�{�C��G����+S�(:P�X�(UD,�qm���uU���h��Ѭ�����M�	����c��idG�2���?��sG�|�b(�8��Q��)�yJ6B�;IU#��r�I�ė�ɣ�C&f�eG*�QG�M��66�7ԡ�e,��X�z6c�n����h�+Xw��+~��*N�8��qp�����{$:0�綰T�E��^Lt��=�ȧ�4��6b7����{������~�)��ѱ�@�����}=�R�q��E����]�����;1#���E�P&��T�=X?c�X �{��I,ײ8�(�����(�s�
�{3��4>���;N��c�|򓟌���O�'~�G㮻���B�=�`|�'>?��?��s�7r� N����'}��-'�6��~������x���1�O���������<�lZ*n�rB���v|g%����j�gQ��u��a�W�n�9�l�I˪�����(]ĵ\��$|F��d,�.�����\%�wPw���õs�i؎���pi>쳥�X$Ͳ�ٹ�����@������M!�.d����@���0�Ȟ�=����Q�K����ߍ˗�c��@[�+���-����G���c	���O����P<��C�C?�Q������B<| n9u2>��ħ>���я�@�?v V��b��, S�Wc~s:&�����R���z�V�����֓�b%J�2xl�w^�%=X�&0��)�I�^��-��G*��d��'$}�wQŘ@�	S�H_b�˼D# �.g��Z'V��dhS���OXq�ZOX�� 5����&��#���Xpa��<
d	����L�}y2׀,,,�c�y0��/�B|�G>�g">�я����8��yܓ9������y.*ۜ��[0�n=x$��cif!N�q{|��/bU�n8�p�B;����3V6!���5�޷�@�A��x���O}�����!���8r�.�-qǝ�i���4�3��ػoo����%{��b�i�k�9��ӧ���#q��q��?f��S�<u�wW�ŗ^�g�}&����!h�33��0� �����
������oG���Cđ#G�w��3qeu���Gѹ�q�9W"g�)�łt&�;�s�s����k���0",p����"�<��
u}��yw+���U�zm�����<7��,]�%�Zϡ�fV+��Jĕ��nm-EOÖO<-8@[��K�E����P�SD�O�����@ggɾ�ƛ��o~#Ο;c#��x�~�(�	��\����ݽ��cw�F�ĉc��u�����D���=r(��ߋ2ߋ�:��S'N�q�������b��p&�9�J�u��X��]EYN�;�+Ƈ�D��kS\c���#�}Y���(�\V	z��㵢Z��?T��HȰBgYC�S�p��F��&��[y�[�J$�A0k^�R��[[Ľ�e8ʰ���*��?�6hvn�����Kμ4�F3�x�|���� F9_fz����C��h��ġ=#1=u)���_�o=���<q����T�L�>>�S?�hiV�ע�?]}�ڏ�o�t�)B���`���U��#cV�a�w��fnT������"9@����'~��g��~����c�!��'���U0:���je�0��G��]�u\��8w�|2���)�W�^�^|!Wn:�h<��3�/}1Ν?>�Hs����Yā��9�H��^�?G���a���s��-XH�r��F��
�	���F���V��o��3Q���_*�)��4�q���W7;�A|X$?P�wX&H�f���K`i�
��N�f�����민��sq��Ŕiï��QoR?Nw'qG�ڱ0���Y��O�D�kl̜2�p�3u�kG",���lL^��=����?n���s�v���o�B��鍾^��6'����9�����z�/Ӿ[=�(�f�T���OW�}o\�1/�p���n;�'nݿ'N�ũ��8ԄQ�#(�>�&�Jo�<�F�@,/��<��swf[��i��?:4.Zݐ����
��Re�#i������s�v^y������ʺt�� w�Tp�;Ox�)�8�u�bFFGR��z�m�+�>����!a4[~4�|ci"�㧁�BAkc��¾�����?��l�������3V���o�;��!�!����g?���}�?F�ZT��qG�����B�T��I�SąMZ�(
;_{�l����4�5����C��o4�G�����S��${����ie��ݴ��ѤBU ��4w���}2����8>8�DO�7g��}�l��J�A���I��3wݕ��Y�����qF����bǕL�w���G0���R��{Ş�s�HW�Z��j=���B/*�:Y�pN6sQ����Yj��syG�L��R"E��ԭ��
��ߎ�;��ղI��P�>��,  ����g�����,󱹴����'��7^;��z����[���ճ��Z�m���sM��������bO�Ym��G��f,~��!m��J#�wL�D�����}�Ē[\ l��n�(Ws�<�7�Zpֱ���ы@�o�u;G��b�=R��r�/4���뱻W��<8 a�=�@��X���qG���>?���)�
�]J�gX�{�5@�z�3��M��[�(5���9s����r�[GZ?��jD*zZ�ِUG�D<�`�˯�{���5q��R����(�}v �zmr	G���qrPȴ�L�����k��I-��N�<�*gp� �3K탱�=s��=���}k��&��h�X�������(���QIs��˯ů�����?������7�_��g�{߻�q�����FE���u�3ϼ��ˬ`)�*QιN��YTrxI7�Y�m�B{{���/�BL�hd5�k-P&�H\��z��T�j����I?7�Q����|�cCQ,�����a�\NKQg�r�OaŁ�F[�������慙I����t5ߛ�tnnl��0��߂P��8~~��ΪGP�*��~���@��̦�5�#on	�����y�BӅ�;>�/�L������G��p���c�kW��|�l��.��G���q�m{�g�j�/��>��=���(���̎{��svp�B�c�V<g���CKq��i�oOt�w�ݸ-�q߽��~��)`a�zY) 7�~6��2<�ҎB��Al :�ܲ�%�G���:��#����qlA��pʾ�����M�\tTw #�-�V\�pWe.�G�ę�wa��
��i�ܳE����se;�ieq.ڵ�;����i�Go`� �)�lHT"�	v�[�:-�]ϼVYk�z���W�N�X��y����8��hm�����R���r�������V�ZM�:�У��-����P._�����q�wzBO,��O������7.�"�<�o<��#q��QL^�[���9�� ��'/�W��������x��o��^��~��\%��V�c��n?�t�I���kme5�rLc�.��\R>�)<9������KK�[?]�@���.���
����tI�?Q�N@�%�i���ٟ�~���~)����a��+�k�x�)�*,5�
me�ny3�zm�|d��ƹ*��.@�i��ܞw�"rb-���8v�0�,~�i�U
d�@�9�J��a�E�B��U�(.c����H4���������=���C(��VG[h �x��������/~��?�{4�c_��}��\i݁��!M���
OqR T0�}M�V&c���.�����ĩ����Џ`i~�Ch:������D�P�޵�N:�sX��ߕ�*�ܓ���g����gfbbb*ff�+��_�!Y��\�R� �h�H�Ƴ�b�g �qw�}��`�v�v,�ҟT������]����]X��4f=�.u��<����n�a��W�k۶�ع����Z���_I�4������6�*l?�1=U��'/�ky���?�5�����0nL~��Rh��W�4�E���ތ���.6C[�U]�������G>����λr��w��b���߿�_��߉���_�s��x�i��8���C`�@���w�ʼn�����v�inٹhY$���f�}[�l��2��+���^�˗��f1��,.���Nѫ����s<���O��+��`����5���%�j�^,�Eh��3�0���i�g�'��x��/��
t݁�ת\�[sYA�ś�]Mk��o���h|�r�Pd��9��ބٲ�<��ՠ�]mkl����bhR�둖�SyU8�{���O@��|W��ȋ�H�-��e�}C{����������O�&��։��oN/�/��ߍ�~�[qAy�����?��_���k?���}�%�ն�f=��*L�n�Ŏ��hi���BK��1[I�q�"'�^M%`q67R܍��o��~��~�������{>�{5�KJD������$�<w��+q6{���/S�b&qM��g��������.��M�Hf-; $@ۿ|�@C�94�o?w?�h���{�ĉ[qyp���:�4�驫�en��\iõ��]�]'�.�k�6�E�W,��X\���Ⱥ��!]�X��VU|����|��m���w�.����BU?U�D<Ri����H��Jrx��_�,�f���a����j�}j2�F������1�z����W����C\��_z"��{=�p_$��a"��W'��: �i�w�v��襥_��+��Ⱦ檓��<��EC!p>�2��~��e�~��]�6p�\>35������R�� �p��u, M�M���(����u�3�v&��`Z)�HXk3��K/�ٳg�n�|���Tl�6E�<-�B�?p8���c1<2���:�Q�	��0A�HNygf�Qf�9�e'���\L�L���k������';��F���Z��C�����IpD%��T��0֡B[+�U�#�]�&m���\Q}��""�װ �;��{�`�}e%��g����?*�Oy�c=��\?����������?|.fV[1z�t8y��!;���;3[qA���USrؙ��Rh�D�t�P����Xw��6��%�(^,���E�e����{�m�%��;�;��Zxb��4i�ys�\�l�KԹ�V	繹	,��(���nb��ԃw��3]��s�'������G���Ô����,_U*F�\���-�CA��usֱ�tGs��*�y�7*�My��U	�c�"�(�Ny��C�rT�(�z&�ztl4�T�6Z�����H������ѕ))<$�[��re�4����@��c͠�bb~.^ŊXp�R�#N�y"}��8��;��@?8h�~��Y�&���;�>��=��x�����=�����=?����｝V}�JYO弃���X�����6S��F�4�з}3ν�z�ѷ���{��g�{&f�f��CpI�m>�QܪOa�<ve?mP:*q?`n�;�������<��x��'����z<����K����<_���(�hc:�0�#�ѐ]��pILZ�7s��%�ץ8�;1.��9�����8w�t�m�Z�p*I'��$�
��.��̩xy!�D*
�3��^5b]Z����W�t�^u鞪��MoH4^z���ן�'�3~���n��מ��v�C�D7��5���S!]c��[��k�����/=O�x!�~�j<��t<�¥�-�~������g�G>�ݜ���9ҍ�>eO�ǳa�K�( �K��~����w��b���;ԧ�ng�5Pθݺ���86����l��g�ֲ�C~	���
;����xi��$��C~q[�v\ ]R�ewL_Qu���=g�b^s�D����
��F����@/��L������2&q$���uV)����w�2�4�.��#�I/�ļ�k�\vb���S�x��{Y�)Q�~L�
�+`�0�gfc�߆ B���nYѼ�����͎1�B�v ��0���L��������fg���3'���Ϡ��cp`(��?��S��k�pVcqm1.O���Μ�C��C}�q��q?�<������c������7޺_����C�t�g�\�v�ġ�鞣�_�ïa!\B!�?��
�V\�p>��p���/e?���;2�s7�;�J^S���#�硖-��z.暊e����J�{��oaQ�!�S��s/��ŋW����slĞ�{��ѣE���Ν;W�^A��#�7�"�:�읳��ҥ�XD)k�\��O<�L��V��������'E'®{�fO��:��f1̀�UL�b�������BӴ&<�$��w5M]�ŏ�m��Rz��W�)���^����F_~�ɾ��VNB�S�O!�c�ex艧^��?�||��/Ɨ�x1�}��s( q��\5���$�s}��H�rt_�c�B�o<��Ǣ�G:���~����E�z~~đ9?I1�������*�%�s1V��#_���9���n+4���ڹ�	��U�h�<l_{{W#��b�7#7y��Zҕ�41�;�#��wrr*���̋/�o��B[�o�α4�x�� kz"�k�tƋ/���M�����:�}Fo�u.���K��f��6lN�rj������u�m u\"(q��0�++(,l��w��[ǝ'����R\�|1��>3�B��2S~����k:�M�3�`ef�!�m�
F�ކ���������������>=�P�r�-1<6B�_����o�����p\�`_���[���s��3g�}QV݃��fO2���& �ѯ\�E�Vbý&h7g�r��N:sU���L,-��]��ķ�~3^}��x�ŗ��'��׿�V
�3�</��T*i\� .�P�J2�f��	}L݀����P�Ԛ� i�n�`h׎�F��5-�m��6I�,�}:�[o�/�
�=�8<s����Z<��'iY����~k����_��Wq��R(���N�ZV�Bv���0��k�)�I�"���\�R���r��~���D�^���嶞����lW�'�������7eQ��0e�u>4�i7�M,�W/����5?+R�eG��7�=;��q���C���F.d{���׵������7~�i���߶�^��_�_����-����C�bm���>j�9��v�k1f�S_*������_������Z���+[�5�Z�U�4u5�{��x��g�%����^�	��S���+o��XtW&fȷtк����J���7ip����6;*����_��`%yTgNVS^V����oJw��:�|^�)�Kc�|�B։��@~�H~�����-+Ǌt�ݷѐ��.o������%�
��� i�uSЙ��b�vlD��QO+TX{���}�2��T���{��F_ot�z�c�}�3߈�˿�.�Ggk0Vh����/<�j\xk6����8�F�Ǽ�W���`�\�O��i��D0iua(�&���q���9�>E��ƫ��U��<�w�--x*K�n�cs�^zg�Z��KN�YAP�R`�-�ۡ���?<:���v�2�:�n�-Q�/�nX2$����UJ_g��F?.���-ιsg���E�x���L��-`�����ō�ro\�s���"�|{W-.����ޑ����o���X"O�z6�m�d��JXe���A�"g�kW�j�h���"�?�|����:]��Ͳ�aEu�TU�2�&���cM���d�n��x$'D����i4�X�R���f��Mz�IJ[H�r��h�s�����@���_��ӊ��;���x�{��O�>|<~�~0G�ܑ��ų��+/R�3����Q�[_k��A]����l �Q�9l����6�J�v:����ƽ�7�T|��6P��ukqq�
�e�ją˗P�\/O�jsv����Ć�я��ŉo�uk�E�R)��{ϙ8~�H*f�����/�h5P��WZӀk��u�/�C�8���b����8��:-�� ��_.�ؗ�G�q7�?�4����Q��"INB���p.�;8�x�I�{❫�kX/�v�"6a#��|Fu�P�`�����Վ�����,]1��0o�A7�,*č\z:��{o��G�0�b���x�������'0gQѵAa�N�O�����=z0n��H�m�.mE��v^�|��w⏞|��n��: �L�w��/�O��E'�u%}����g��i*�Q�K��o�8��>���l�.�ǭi� ��?��J-|V9<B+�s+���SϾ�˚b���;���� �;�Y@���G���IP-�Ƃ���Ζ���Sv�5�H<��p#�燕6�k|l,n;q<\��EK�����Ŀ��/�Ժ��'��,i��{A�Ѯ2�����8*��H�A��W~X��7�a��f�|Z*+����4��:u���|��
�#]����j�	cMt���w۶(+�bTy7l�pϺ����~���?�h���������C �r����1=��DQ���1-�E}����8q�Xc�>��3J}k)��wt����~,���,��v��O�D>@ɡX
4x(�7'��z����x���]yb���'(^�]���^�^ή��"σ�B!���Q�V�P����t<��4*�zo����fH�ǝo�7"��?��X�r��t��Wm*��4�+���yg�Uu�)��ͥ� �g,_���O^� �A�91?���?p,�Z[��8�;�	�mR��J��y�Ph9�O7���D�u�D���k��[WQ"Cd:�1�Ri����[0�F2T_ϻb�;hv�"�!��c���P+V� �d�ݶ����)9��%�,��	���lC(A4\���7i���+:��%��-��/���?�c���v���&�+(����s�FaR�JT? �4K�9�Q�{�Ꞣ��s ����.�B+3�����s5h�wW�մ���8��sjuC���_���>z|��8��S��51����fsv��W�V/�2<)m9No'"f-;��;�)��`��_;��?�W�ԫ�c�F ���s^��=Dh��v,�l�C]X��L����c �Q)��6��wm��5,�5�\3ra��:�y���8�
sUE��n�؅rr�������舿�W*>���b�j
��o���۸p~�bo~An	^t��Ah�mТ%_Y&Z������{�Qh�n���F�ȷ���u���@*�lM+J@�+7��a�-�VP"��ҢKO7��+é,���{b}z!����c�6X�N��������u������U���:�ntD� ��Q�(˲f�c�Z3���ײײ���eI�$�"ER9�nt@�X9��{�����wou5PI������/��}���O\K}bua��ܽkh]>r,�=��դ��~���������l���������\Kw�K+Z�J��ك��y��2$��o����k�P�SY-�����F�6�e�M����<�g��B�0��ZpY��;��y>�ƇϜ9Cf�cz�)7��2�����[��8��[P�a�3����򼚢�Ɲ'C�C*1 �BM��yIn�Hv�iR����٭hï4���f7B�e�M�������RX�IiI�O��].�s��w�s+}��1�;�՞�Q,�=k��k͸c��n�>����`WLLհ�^�K�nmY�;���!0��'���Z��=�ĆMۢ��֝ S�Z�C�v���ӏ���Ԋ���2�n̢��\�8>��щk�Y]k�C��ş�ў}��\ocF�!�rUuW~k���1d^�+��
��|�b�9�`=�����@ ����W�P���mۃ��8���=�.��xi�q��X����p�/$yr��[�����ˀ�l���q�⹘��Q{+g�8�����+1˹{��ƌ�^�H���TL�v�\�#×c�֕����}�t]��8{[�"-K��ܨlks��G���u��nئ�qAgp�86�ޭ���n�k�ƹ�Gr�5��������[k�a*&F/ĥ'�'�>� ������M�ǎmkp��y+�����l{|/�u^3�Q ���!AПy	 L�(��4�����V��uZ���Fkܸ{Kܰ��ۢ�T�1��%�JE�F��:�33����#0��0�o���x����-c;ZޱM�0p�J9Ν>�GѸ����g\�o�RIs��nn�v�/5��gb1[��	-�L1��մ��.!�:s�%�C��Qy���
Ȧ��ч����
כaTD�ZĲ�i|AwH�[�qp�O�&I_���<�_�xGK��F(��p1~��Oa6{#
�u]M`.3�X>-%5��N? z㾽�u�&�. !�}r'5�[ ̩��
xn$��Ʊ\Ŵ��1�wmc���ι�[1�0��Y�:#]=�@̟� ���v�m[�Qzp��źD���E������J��V�24p�V7 ϥ3�4|�2h�,��l�]0��Dۈ��G�e�e ��i�7>������l�z�ŗ��'cDņ�kچ�l%=t'ms7��Y�(��]w�/��Z}�4���\(� q+���.�%�.�5���^���m¬еԲq���L,651B>���(�(ݬ��ɹf�s����XWcj~���!SŬ
];8�vl�M��3]�'����?���P�Ʊ2v��+�5m���
�Ex7K$��A�s��	 �n�xj������O�7>��щo�D����nE9� R��ԝ��x���І�qal5�� �Cgc����*�=�Fg[5Ο9On�o}y}�yjV��f��`���*�#�-�2ñ�>���������^4(�%��0�@�jNeV]״A>�.Z�
���Q)v��Sa� H��hv��֤�����8祕͡��1)}r\w\�4��P�sSc�7n��c��1����5�5U ��g��j

���be4������t)�A-�hLia7#����de�����v��� A�g���4�����c�����<7�R�	`���`9��7e:�[>A� ��`k�`�*$�T<��5��&`c��ۅ���������M O���)��p�oW?���}4~��>��q,ߚ�h
[�u�0�Uɞ&��o���b�0��!�;>#����{�LN:Y��ؖ���R'?}���7���(*U��"rZ�2
�|;����������k��p�'�b�c��P�Ȉ�i��0w�er�^DҠ��ҍ�P�ԯ�=*(��.�~�����O��'sM��#��=%ֳV<��� 2��D���z�>����4���s�e�-~�S�got4�cE�x�G���Uq�K�tQ��_<w.�>� �3#ˀ�S���Kibk���f�1�0o��]qA!12�K��9\�w}Lѷ�P.:"-������&�bm>לݥ�����cbz��I˼x*���/7�$W)�J̱6��Ok
F�jpsm���U��aL�i��E�J�zh��קp�ed[C����%��	˫�13r>�o�C@���u�ؐ
��Fެ4�֥s��\nN��6�ye�A�oR�Z!�c� hg#(o%#HP�>��W�D&�����S��y��i��5�`�(��<if�O��_(<�Bɯ��+��=���!��3�4鞪��V��-Z)\-�o�=x��DP`m۱��ׅ�).B�sz�{�o~�Wbh�Ŋk����f��:cZ�LKҘmh���	���ɉ�,���==ϯ��C�U�����"��O�,�6FJ�H*N��r8�I�l౸iߞ��o��w�D���v݁�-S,��)F��_b��m�ŷ=Fs;�y�ux�r���{@8hR:�����/��Qk��� d{Բ��4��AK������s��UKW�*���ů}��������T9�/��tm�H^�D0m<:s�d�>uˣ�./Ɵ���q��e���B5�.�\Ι��jg��s�����
�.\��Gu^Y�̳e�ƙw�s��
Ȕ���C�`��A��6Y)0��1�v@DKDa�s|[ i���R [�r�@�v4ٺ�J��?��Ο��3�p��(wt���%��X��ș���m�ɘ�|*\M�px>I|�ƖU�
��
����Vg���Vk��ρgZ!6�i�
 ��t�Ia-P0�LE����ӈ��g�j�;D��Q	D0X��$�>�}n�����"�FR�gi\
2�/���Ca�� �7���D��а9DEbS��)w�G��i���l.`y+�_�c&����q���������=.�w�2�Ma�"�X�Ν�^�ݴ}Gͭ7� �rC���n.�سaZs�(����/Ɨ��U\�gP�i�]^qRg�^���pq)��5����|2z���:�aK��o� <����֪�4;�Vg7`@�\@kxl,N�GA��p9ByE%a���K����^��5rQ#�N�Y����WZ���Ć;S��� ���V�S���3�Ȧޖ���O���(ßW�lʪt*�"�ˎh�3'N�?��<yy!��W���H7�U���a7�j��RG\8'�����]�b*�]b�ACິZ"��cS܇ K����;,����k���Yk�8D{&t}4
5� ��ꃶj���Nsb����Z���s�c~rB�����
���wtE��7��F
I*E[�J��}w�|L]:	p�0��Nu'cQ�wC6���$�B����(�LU2	��A����rj9����"$e7qZ"�ي��Uƿ���7�K
!UpL��xZ����NVu���5�,��H�B�o�U ������E. �	�aK�844%���r:�%��?��c6��~I!���cԏ��ŹB�r�Q��܎j	`��,��Lw2'�Q�l<�2A(��n���� ������`2љ��9����eT�tI>�}����i�6U����^���l�6N^��m"�U0ӕ����n\�*<�Ug������(���uF9e�i�H��� ח�muiJ;2��a��EE1��Wd��7���A��� iz��?�@|�}�H� �D2{hS���w���m0�9,��X��<o��_>�� c������L�j��U{�B�����<P�D��#�,��܌����������4���"Z��4#8�����G�-�@m�AO~�!��ݻ(�`�`���/`�h.A�\�Iw��R�i�'�.���+x�v�j�:z���w [��'��yDy�<Z���'z�b��[0$��J�
�ꂙ/���! �d#�kQh=��tBB
��j[�)X���k�NoO:���2V���=M���F���ڮ����?�r;E]-�<d�|�~�Ez����F�h�|�9�*x�`L��9+�O�r�*�Zv�v�'��	]Z� @^�@������z$�)������r�B�%%��� ��(��ݘ��)���!�|Am�^�Y�v��Cr	I/����R�0�����etȁ1��5����p��Tҏr5��"��N�s��U���<�ӔK�I�j�����mX�,Z�u����@��6Ge�pa6�g�x�E�w�J�.�{�s�f�.��Lv���������ښ�DV�P�=0&�O� ����f�pF��V��O?�B�LF/ �A�g,��a2zn��Ԗ�o�9���M��!E���3���Q��쮀��s�27�0cۊ����:m7���k5��U�����x[�wnqV�+}�7_�O�*Hl��3јs�9�|	�_�Qr��%Z\�	v��+��$�F7g�=J�M[Z�%���i-�}�h s�m^70t����}�
F��%�W�I���H��W�fYg������I�����ר�kc��҂X��zB�t���� ���§��7ϱ$n�޶<�C)����}1�T����-KG�Ǣ~�Ejލ�/bON�GC�Z���7����@�e#��h+!`��%�K]�v��6��Q�k��=�Է��ObZX�1G!ף�F��=���s�|- ���V�F_=(�ިtzދ;�-�(�2���"��yDPKX�ީ�;{�o��j��,����~��lL��t�|�P<M�~=4�[P����/l�� ה_E^��{�$�����P,6�:<۽x�������̕LWh(?~m�Z��i��3��r���-(9��[o�|���-�6�37K3�Ѵ8�{�Vp�:�%��l%�s�[֗�K0;���0�e���� �g��! w3/�́O2�̐��p��d�/��)PZ@�7�-QQ#��	$���ȷVV��0�^Z�G�m#:���u��;��?��jy�Z�]�籌�}������3�/7QZ򜂨4ܧ�~���������#c�kjZ�׭_˚�� e�ةy�i��qM�>����ʯ��?xE�#j�Yg�z�㣏�������;�����������D�i�p2V �v��s ?yhDTǉ8g06Jפ/�9�-]� {���l��Mȝ���k��<;Z���K��Z���D^i sF�Lp�q��3x֡�X3r��f#,t�P��ɋ��+�:5�~�5���u�j-/s�2i3��p�I�SO�N �Qo2�&#��5��}�j44���P��������	��S�	��f�5��.�4~����c3K�ܙ�/dp
�]�.̔\twzr*�4�Nd&-l�#��S��4��^-� �D22BQ�]�buV1C&���%nر.����7������� X�1'j�JT�D�ʚ�~����U��bm/�u���Yw��]7�rZ6�NZ �ԇ�1���|A��H4A�L����Sص4�����D/�r�5�)��<OX�F��#��|[?L��]��5��)�����P��$���ц^��_��m�N0(O�!�#�y6��K�%�j_S��@�g㎛����;�m�ӧ��>�Q),�Łݛ���n���C��O~(��!v���:;�����u���D%����˗py�T�*ߌJB/�V��ek !��㲴 f[Tq�<R��.�xH+�)O֍�2m~��U8���|F��[�g�g�֪| o䰆V@�d�Efr�a9�Ew;ێ���Ie��H��ح��[������o�JKU��{o�7��%��yq9�na�z4r�g(�����ehf������nٿ#�l �Q ��ļ�i�DԤF��+�X;a���t�y�b\r7;�4cͱ%$�i���ff�X���?�^��mQ�zn{��i��br��#���@mq:���C���<������=����a�樶6���8�����wq4idG���%����[�x�����I�Ʀ��	�����j�&������_AP�F
��#�aݜE�	w���Q��{�4��i�:8�e	��-#}֚������R�mGe@��P
y����AF,*�
�� ��	ғ�k�� B��7�5b�{����2�cDr�?�,C�[���~#>��_�*�ϼ H쵸����7�񩏿?v�����X�m(�Ih���{n���rs.�p���lR��3K֎��9�nR1�]�e �,B>I�B9�Tr
��O� ��� uA�GǴ@���
�M )��?�(����� ����j7I��|�XZ��oX_�ZO W��^��o����t�J�;3R��s� b( ���q�y|;(�|,�/���X\�1��"����h�{�žk�5���[A.��!�F�����v^r��|�y��T2L"9j��J�q�]�Ȫ�խ,
n����m���͍�v��Jr0���X�߻-�����x�=wǖ�Q��]��[7����틻n�1n?xCt��cl؝�҅q?�dG�r|�ů|����gN��a�c aő�ڪ|O��Y�� ga�-���i������P-���9D���Ř���Z��H2��GJ�j�"�\�3
�b"����� o���B�<3�9�f6] �m�!�1y!U�$�J\��B�X�☍��3$��W��?�y�����x�2Zf. Bވ6:�{n���?��x���sx����W^y3�fj�oצ��_�X����3�?��_��{�>���7�Ͼ�����_$wN\����[���x��c��G��8!Rp��)�O}����<Yoi�i�qްS23f2uR��Y5�^+~�8��um���IOi�P"��YG�Z�B!���d��!�7�=� �gQ�KUD'
�N �l$�oF�h���IO�[�w�
zdސ?��^C���`��"Z�?"�]4A��h���nD��=[ ���6/YKk�H�"����ŏ9�Ϝ���	�G[�q����"��@�����:�P�̤=	����X��5�L��
"'(,��ę!�	����;�����7	}��8r�\?y9N��DWcӖmq���b��M �HL�]�ڼ;�A�Ź�e��{n�r�G��7�:�&����|U�H��1p֬��	eJ+*�C�=� P l���T�=Van� �PkIG&�ғ�-֙c#"	  �YP��fT�`O{�z`g��͒����kc��5\�~E�y��v�l�m���̤��U(�����Uʥ���(Vq/��h�8�/7�te�@ڸ����X|��{c|x4�x���������t��_��G���0�C���y������\�K��<�������131۷l���/�o�u(�j�4��`��(w�Ӱ.�<E�?|ֲr]a�\��yq��&�9��<�h���`�M�]�n�xY��}�!�*��,�fmQ��V�3eM����/�a����i�r�z�[��e�y�'����y�"�`r�3����|�5���\"��?�Ch	i�j��z%�3n��׺Xŕ�f	�|$��e��&]���Ws\�|!�s��u>|>.�NǼH�Vm��v�sMoW6[���׉�5�Iq�!g9���& 8TV�i�M{�I`�)܎�5���7�6�m�/���ƿ��o�7�f<���x��7���^�i,�΁�1��7��wݴ=z0w篌���Xn�t�-�b��m��/ǳ?}%:�kbr�qXI0�yM�K��7LfA$[�EUK��uՆ?iCؒ��epR&38��.j�9���s��e�R���}��رy(6����/�Vp���b������~ �����Q,���;���x�7�{ Ļo��W�bd|$FpZ:�b��5�B:��+�K{G�pќ��o���s��{���[\�N>!M�q�!��]ͽ��3~�3�-@�;+q護r�]�V�}�=�Ş]�S`��x��g�K5��(q�lo�����1����쉣G��O_|ުP:@��I�o��;ж.\�?7E��$yK�����P{�!�'?���B���:̴9*����%�*L",���
�m�%X�h{�
=��C|�̦u��h��p)�tk�2f�~˲�t�_ɔ�<�y0_��rZ@�)���+~��_�B�I�-X�^�g
��2���jǝ�	x�:�v�Ɓ=[se�����Hp���͡TDL$�>45�m�>�_*���T,j� M��,� T���n[f�X�����[HQ�t."���{ �V��{�o�֯R�+151_��7��׎���i,��م�2>�:WF'����ܜ{��a_�����0�ذ~= �J:r
�*��B�A�r��ȭ��v�}C��f�95br�D��O]ma&����#}�&����rq�F���mn��[7������o��'����d������s��O}"0�L/��/��"��vKl�vCl޺=6lښ��Ƨ�b0+��|�%{Ұ�J�����4�]�`lL*E^�k��6�FDs�ݐe�s{��n���(z���[�n\���|�"��to�o�C��	:�M�����cWrQ 'έ��¡|���y��شi]�u�d<�����7�5�!.���&��^F��(�OM\<uU��+���u����G�W׈)7�Cqw$��9ݙ-g�7_!�嬰sȧ�|7�.��2�|�݂eօ��x�sMB��l4(�E��??�kū��D��1TZ"��]m��7�ά�Q��a�3����	"vK��m����D\҄j˥x��3������������`��#�4� bC��$����ߏ �?-!�HZ��=qߝ�EW���O���N'� �0*�C �kM�9g�ʥI��յܹ��vl�1���5vl����A��������<Y6�p����kT��̼G���32�bC��\Y�c(��A��Kd�5H]� x�@�;nEPw����7>���EWGK.�866��=?�|27~~�͓�{����o?�:g&ݿd-�k׬��Ck����X$�����n�]�|��K���� �8�v��s�L��՘�x��J��-H�
������-]�m۶E7�قU�s�V��5�������5п�=�:ch�R,�rNQ'yo�����=����M�׾��8|���S����'d�<��$�pL֕ݨ�:�g��
M�x�������)ՙ�W�<^����X�M����(mS�I��~���W�C���\�yy�g����)�'��Nz���:������:�fM�H'�+`��Z!>W-���m�b��M�<?�;Ӝ�êT4<l��7�b@f)�k ~(�g���X"TxMSRc�y"�j#�No~w�B�Q$I�Lv{j��%
�=:��$��d�ڹ��Ck����x\�t9��`f4����ťf�p&5�[GO�,�M�Po��y����_�}���kG��^���!*�pˣ���!a͏'���E���D?����bf��	-Z,%�c&TT�U38USST����'n?pC��T�������C�>��Cq����7�����?�m�Xl�3W���+q����l]��=�sˆ8�R<�ӗba��r���������d�A���׬䢢f7�ļ�G�s�Y�q�ku� V��˗c ٸa�Xg�]�)v�>����6.݃Ю��6c��;pc�9p0�{��xϣ����o����������7�_��1��{��7��|�|�@��k���|VZ�X&��|�^����\��~�w��O�_�}�5���"��;,��J�&�E�<����W���2�:}7B#���[0
:���;�����P[ #���F��[��4�xu�;�Wṵq.��xW��SkO�߿
"i�d��� 3�{�c���\�u�B\����Ax�����w�^$�Z���eS�F>�'%�+���� 0[6o����"�y�c
� ��ƧYZ�aZ���܆�����#'O�k����ϝ�]�����4S�-��h���y�Vs9 �Țc@̻rug�*7�̒m,dv�����:�M�Sx��m�ᳯ�Wۡ�c������x�]��Ϟ�[���'6����������D[�/�c�tF��-.�<��˱w��ضqA�o����^ (���k�,�J&���0�f󙷏����^.�jW,5g��ھ�_L�9�ˋ����BLM�S�uٌ��
yd��v�#�w~�<�|��x�7⯾����O��ѹ%��x^�7Ϣ�?�<-B��WP���4o�k��4�x�ڵ �1�*�1�|��fq�����1/f�u.�"����-�8�$Sh<�oS�KL� �F>�G�����/hb�����zBצ���I�_�m빞���pץ�.�����fA����1Ѓ����������ƦLv�\O�M�\�xn�9^ם��Ha�P�:���\�
"����(�>�+�u2������+��C?ݭ��۵'�1�Dw��8~�\�=?J�dۑ�X�0x�R�:� �R�q�X���ƺ�;����������ci���݊�v'yI�M���.3J�F�;�H��z2�tӺ ���B���˜��"����J���s�A@`}��,ž={c�]�wϾ�a箤��Gq��G.���l6l./�E��d����7��M�o;ϼ�V�E5�˸.Xg��|�3���������ẏx�����ר+���N��=��YJ�s���Ϝ��^;���񓧞�����+�� ��L-N]�׎����|$���?��W��?�q<��+�Ʊ�1�P�RW��[�7��t2�������b	�d�z�κ3	*c=%]���#����=�+����w3���t�
"Xh�&I�H>�E���w���0����n�w
K� �|'���M�烒蟹�LԟO
���`�D�z�H�%vm]7���9��E��8�$!'Š�ڰqU�|��WcM3<��������-6حF{�4M�;�_��p2���*.D�d�E�a�� T��� ^m��j1=>�s3Q��R�A����)��Mq��b9�����q���<F�Q��Ll���q��tubnC�V�������f��w���h��w�;O�[j��Ȃ����d��[8s�إ���kI�G�{{MJ<�D�g�峫8+�(Cʘ+�^;�����m{�������S.ר4^�������7��DDu�5���c�����#w��ߚ�}�[��ޟF��.��	"	���f
��M��C2��#���)��y�\��t:�
'���"��Z���:8���}1���� ���E�T���N�\�E�mk�\���������Uw�/fRO�S��^��B!�  @��d�"��ך���[u�=�';,�A@)�D�^ԙ�����6o{>�=i%� !�q�c�\�jwo�(�,J�Ņ`2�g
X
�]��.J&{�,O��L� ����;�`��e0��l���C���3�0������E��<��QL�s���u��/=ts�ڇ}X�.�@�m��-⦣L�DD)��HA�����ӉHS3+���s1<9C`e ����%��`3�oHK��׋�Q�E+`��ܗ��r��L37m� -ε�I���=�3w7��x���8�22����Ni+͋��s�)�ӻ!��
!�+���D������%Yqn�]��_i�E��Zj(-W�����\)~S��F���J����
m|�sM��#:�*I֝���.U�����ё��:���*]1��ͬ�ļ@�_=�;r�|;w!�9_Y���o���ۿw�vK.?��k��k��I?7�`wB�K�ʗ�*4{�dTh���[w� M�iXYʣ��`�dFMYp@\��ptƴ�Z���f&���)j��Q��& ��p�K7מ�����Ss�~F��q1f�|��n���Il%�KP5�I�*sU�S
�y��fXN��
!/b�NQ�����=��r��Nl��;��=2��=�}��� ���|�b��S��5RO2Ӓ�E��A�!s<P�_X�u��ƌ��G%D ��9IT��/
|G�+ƥ"�P�YtWy�oܼJ�w.��:N䶃7ĭ�6F��s���!��� ��H���˓���(��cěv�ڰj��� ei:ۯ�
_�<���Eb�`�)L���H|B9*�6;- V;�I��g]׵�w f��/�X����:���^]��O���"���˹ҷ#�QGw�s�)i����p�/�����/�I�7mI]ϽB��xF���<P5ǐ�y�{?I��������tug������Wތ�^z-�8GN����{1�y�,�Z킀�qÎ�q�-�縌�^>�Wߌ^;�r�h����9� ��SZs���g�y��d>S�� ϱ�>Zj/{Ѡc3���Mj'���.M^�~����R�߻#�����BY���賹�oca �����K�Znf$���sÆ�*Ubεv�v�t�5b��z-��㱸^)Kş!����z�/�����/N�+�;!��\>JPf�/�!�8�I��O}��ֿ�`��&�;���r���خɏ���~�n������w�����>I�����D�w����9��rgo%�2%%�*�d�T�f��9���fo9�'�6$���3�:�Cn�fϙ����șqs����� xw�^�IT�Z��jTT���\"�#\5�u�oQk�L��%\����0�3C+m�/���wG�f8i-8��[>��K �:�M�6����o�A6,j�R��Dh�� `3����H��p޽�M�t��m�����f##�q�8M<q�l:z"^{�p��4�sPf4'�P�_@��\��P~�Oa�I_.����ЈXsa� )�u�Z�k+��|�Zɣ!�Wa)[�&�o�z��T��*ɳ<�i�	C��t�Z�����{o�{�3���ػ}C4A�����6�� ��y7��W �̓�q�[�������E3���'s�\v� ��R��U��K�R����z�o�;���G��^3����Q����a�����'��1�<�&"� �?�\�}�j4)x���pm�W�2����U�K�E9�i�;��]����)��n>�"�Yt'yv���Q�;� k�� ���� ��Lz0��C���8z�x�Ǖ����W���_?���<xLC�u��ȕa��9���;���+p;NO�0ù�&l	�,��0eg�G��B l�FO��u�w��c�;cێ�q��x���r��2��L��� ��FO�b<x��غimz�5����[.ǒ[E`�M���X.p���>��~{!7֦ݢ@�@��'��D��I�5=%]���l�Q��_�׃���sS��y�ܤY�beQ"h�{��]w�_�D�L����>�;gr|�|��v�@���T3��z�KK��)����Wh�kc�q�!��ήp�7ǉ�7��J)զ�����/�c?.Ntv�ݕ����,�/\�/}�K��o|'�yJ���Lw�q{���c���1�K����,��_��Jw!PI�dy'�]��JV�.��O���Q��y:�l�/ی��F����呟eS(R��� /<!��;�s�<M�Ɖ=�d!�Fm;�9o������FN����^�+�]������Q��y�����p�(J�;-�t���ܫ�hn�}��ۿ�K�чwE'϶4��H��{�=ja��������c�(x�q��E��i�d��AM\Ɲ���]���<G��igֳ��ʂ��sc������t�����B��{o���{{|��;n�9F�G�#�^�d/�eڙ���0������O~��سm}��t�4���85�2��'C�C&�����j��$�@a�a͈	���p�>WF[�Lw�������dlhx�k����;��i�j"V�&c�@W�u��X�]��዁����2ϻ�L��V���%���Nh==T�|�
6�	��\�mƥu+yj�ZJA�?�3��捊{g����2Ӓ�p�� @ۈ�bmO9~�3�ٺ}���O_��~����+�blb,��*�q��ؽ{kl��T��[n�{�#~���������o>򅿌�|��1�8��޼w��ڼ.T��������-���5ǫ�&i�w� R��<l�7����v�������n�Ŵ��MDk$���l�{d�T���oH���������N0[��^�NA�|�]c��*��W�N�>Un��q�]����
�*�q�m��-=��;�.'�r�v
I 1n�Z�ҕ�199��w�[G/���W�h5A
qUp�ήI����d6������s�D��9ś�m��G)� 6���,��Ï>��]���>v2~��q���_)�c�qױ1�H���;vl��wn�o�!֭�C�:�w;�n��0KD	�V�i�Y�x�������g(��j�P!�5S�Ҥ�g#���|~х��(jXL��j�as܏�����|��x��7�������cqn6{tj3#Xq������~�Cq�]�����q�ĩ���0h���{��%W@#6VC��X4�g=�G#�O�w���ex�f���w����x��;�S{��Ξ����_�qbd>��:���m[�G�w��m�^����=q�B|��O�~���^�a��:�\6�DR��Z�W�V���`�g�g�96�u�������.�o�Rߧ~�:پQ���8�� 8�] i��p��Z�
�@R�j��j��erW����|_��7��1�����X�E~T卢[���?�g��SѰ���D��@��ԕ��"��S�T%��K�sR��<|:N���H��;I;�n�t=�w�G������!u1X��W����D�z�S����RB�n�������+�2�\|����g_���<�e�x�3��[��U{�j�� ��\\<w)�����1������o�3\��^�8�1��
nE)צ ���n�`޵Ɩl7�#���ء���LE�q`W��ݿ�����N�	§�MA�����wr���7lC�wQq��k�x��G0�{�ȡ7�ʅ3�a�#����\�������<����7�/��<�|T���ɬu�J�*��Y���� W�܀��O��X� n��cc*��~�|�VLه�)�����l����������R�ژ�J�x�d6oY�XW5,��lk�ı���O���GO>�|�˹X��j�V�e�������u☛�X�(�;��G�{r�֗��sKf��B���w�=��ME��
� bo���6�S'��?�n�D~7���P���w	~�� �i[�Y�����|0͂?d~�i�}�ȑ=YѰM$!GZ���q�7Ǝ��?"&��\�H�U>�����R:~*���+���֎H�Y,�������i���iܤ�bT�ta����Y||lm�@�brt,nBH����|���-���zM��qjd*����R��G`q\�y��D \p��\Zl�7^}=-�=�vG��W߈�_{+ڪ=Tr����^h+�����:��*�)����i	�˧i��B�*Y�� \a��,w2;�e�����
C�(��8���?�q���I���Zq������ ��ضc]�|�*�?~�3���/�֬�^9���?��w�F��,�e k-��� �<�#��`
�E�],b� 擜ןwlt�Me�p�. �� e�t�Cw�[7��^��'O�6�5ۧ(Oiy*����-X���ek=z6���ſ��/�s?}%&QL�����6ۧ��eΡ
���"�D����n����!�p/�_��E7��X��e�l0(�m4xR��
��l��~�lN��V���uC!���I;�> �j�Z�����l�-9��@�D�ϻM��P�3�9����۞����8�F�a��׋�]��_�GyOZL^�ΛiX"9A�Һ7��7l�r+�r)��ܓ0y2&�!/2c�@ 	�^�������
��,� H�p"��򮌑�}�3�i�rtm&u^�lݲ9��(La�����˹�Co� yi.zb��B��[�l�Lb [2���}��Wpc%�`�W$��k�/�����E9fx�5:�Pϭ��e�Ys{%{x��(N�6��uR��n�_-��.k��_Y�a]�߰>��O�����?�����������W�����J�,������~�W���w��R��l<w�l���ǿ��/�0.�.�(t�-!W����e�@gW�Ty��֐n�a#��������A<ggR&�����z'%�fE1;63�# 
���,�fDoZ����TT"���5��� _{�'Oė���q��1�=] t������Btو���T���~F�&�y��k�<����o�<�����z�Z6oe�Z֍o�����k>c��p^��O�k����_˛W������!��G�甫"4��x� ���F����璬�~�3���bq�z��Vx� \#ݍW���"��d��n<A��~����jq�=2�@��-��� ����h��57��]cn�a��T��r��L&Ȕxju�ށN�;�KҬbٔ��hqv�t�bۖ5�e�l�tlCp%�J��N�Wa��(C���\�O�S[��k0��v�BЌ����т�R-�з`�� 8��
e�R��jT��Q�� �F���x��7�?�I�8s9��-4��K�w:����b\��{�P��/� �������ѿ�/��鸲D�1-}�Qs�g�3V�M��V]��#�l,a5��Kl ��R�F�K��U\@��ͨcAک�6,���Z���=`6�4��V�n�b����x���>\����������@��Lt��b����������`mn�vƍ�7���wum����������6��V�^u�`��}����V����m�Ch�d���Î��=r9��C+ ��ǧ{.O؂�K^\��7�i�`�z�A0���*n2şN7�Y����m������-2�Q^l H���BC��-�u�����.eJ��"��Pk6)͵F�H~H��(��������ةq��(L��!����p�m�̴0EeP�l��QPSZ�45\��F7�Ѹ\r�U�5�1<��t��Plܰ��y���`�����Cm%�my:��h��c��<���q�M7ć����}��D��?/�y"z7�8��r�M*?�&�@׌����3�\��nI�5k����7���e��V�f@����[�u��&�VM�?{������<��h��W^�~�fm2����;�Pwgt�ޛ/����O?�r?v,._�������e�R"_v7�Z��3ls[���o�+����"�4��;;�]Ϳ���8 Ȏ��A�3��¸C}��?�ĕ+��cӖ�i�8p�M�w��X;4D�q����;v�}�o���(�8�o<��~glݾ3F�&���K��X�T���u�&�z/
jQG�Í�pR\�/��+��gE�x8�z�s����P�n;׆�=�3]�O����gB��p���ܳ��x��L��ez��!�<�B�,����uy�oM�g��-�)�]���ƽz�����}�au�v;+6�<��d-�;&�_"��t��9^p��8r�|��8�x��\+�h���� �͈�e��A!��3�uɑ�d����ȶ)����t�+������\&���7��1y�\���peWz_�N���js��<�?p{|���{o�[7!�x�c�ů}?�^��6w�=�jMx�s����Z`�����.�2y\�\.���|7{^mX���#�tr��<R���������\k����q��	R��5�����θ��[����������o��W�ĸG�x�F=��Ў�͵8���S���^<���F��l���/��R-S. ;p��X̠u�J=�=���m� s�:sА�.��~�����(���Ex����Z%�2�ܖ��JGota�۰9�<{��Y���X�-�'�}t�b�X����F�U�w!����� ��)j>��iiR�.4��-�y̞�|�)��o���V����~�L��m���,ٞS��|�c��o���|�'��-����AĬg
�	�T$cz~�����I��8�}q뾭i�����yJy�H�,  ����iO?�,�v��BK�շ��'^8��8��S�[l�{{z��9����jD���Q�e��P�¤s%�*��$���+aWp6|�x�ך;��������(���
q��c�O��G�T���K2�P����vEg��_'c�v���� ��Ӹ=1���^�
��"Hr�cAE+_���*F�Q�ќUsf���1_�J��3M��O��&i�F&�|�h����?z�-152���R�@�[�&{�+�6�C}�b�%N��KS�1<VL2\�qs;}6����ĥ�٨�T 9{� �#��̫s-��Bjl�Ҳ5Fe:hN&�P���XZ��EW��R{G���<�k��������a�M �m9�o��=G���P�~��,�M�Oa���v����s �" ����ƓO>�.��*�.�9�Z�ܣ�s.J!x�{QZ�I�`ђ����+Me�yU�I��L�!�[W�"?j\�]k?����R.XZz-�+��f�<ġe��h���,��3�����rH<@~��;K�u6��Su$浼��!�f�\G�-�t,�D�婃��6�u�ق�j�u�~����'t]����.�%(�^�7�,#|���ug�y��h/w��|s��7��
"��Ն��2X]D���3y!�]��Mq� �u�n��]�Ա��:?1�yv�Z�~����{[6ƣ�+��`��t�¬FG;��Ԃ���\���
�T�E����^x����O~O=�FL/6������t�;������P2W��X��f����,��֐�Ȼ��g)��/�`6A�4$��R
����t ���+�x<~�W>� <W2i�@��^�
����pa��|hbr���:�O�����q���X.uQ�%"և�����6d��z�s� �M�>n��]�f,��Ź�����F��n��90���|� �{׮�"*�l�wYcZ��Ύ���^,�@���G�bjj*�gfRQ���؝X��R[^B�ղ���:ZHK���2=�W̦%�DD%�Or.��⮂�ץ��K�H�D��c�'�����G}���N�iy--�A���^����ޜ��@�t���Gr���{	"���	�S����)������ئ����"k:��������b�iq�	��%n�@"��,��� ����5,���m��o>����%BE�|M�3|�����õ%vG�F����9r軲����D��krK�;cd4{1��s�W{B_����L�,��m���溽,k���~[��x�+Ŷ-�c|l*N�<�o�y��ɘ�AK��OnY����6/!�Қ��lΰ�=paބ��V�"���؏���w��% �����/�������QW��l����<���nP��[+�S�.^ș���k�[�
��i���!-��g�c� ޕp1'�´�5��V�1Z�X;��`� ҇���'���B�QN���l�ji�Rh�\����g棌�Q��q����(�D�v��;�&������#{ut�کwG�:g��ɓ135��6]U�M�ᛯ����u5ܴZ� -雨��U��e���5��s��n�PF'��3��6�I�����z�QO֫�ȹRu�X�l�Y�+�Z��e7�o��:��k`0&�"�8�E�&�hZv-l�:��r��u��)��(�t1oy�=�@���
���^�.��`���h"F�I?�m �J�Sڴۢ��?᭹9��h���b|��ů~�^ ze#7�E�������"�4'�5	���k�A���?Dވ��1R� ��7@D�դ\�3̻� ��*��"i��|
ە�]���v�5_�+��C6布��	|��c!�A�JkZ�t�\�`1�ПJ3�]X+����l\l��L/�߷4k~���$��t�c5b��?�b���Id+! T>`�BI�i2Y1ƀ�!,���P����rVs+�D%�G�
����Li�5њ����Z�ID���~_��y���M2'�ߊ�����5ʘ��ib��쒓9V��*�O��Q�Y6-�@��Rc�e��<.F�n*�_�v%,H��V� �
p�v"=kbpw�a>����^�_u�T1�N;��ƴ��
��� ��؛4�c.��@�ӥ1�ԑB��﹥��(5+�1���V��9]�XE.u�.�⎴K��!���A��+�b�_��+��� �}v�C�r��T��gP��mV��]*�ܕ�r��.^����Y�"CWC��"4�}���	"E9�"T=����GbZ'NjՊӊl��襺Qț �u�����GD/����\�|M,�ƇM����J�U�XW���2���K#\s-�����N#�,��\f�+��udI�J����yy-X>M�U�l_�t���a�ڬ�D{c`p}�H8��Y���C�S��f�ʬ,�Ԛ�+ ��`�t��\d����@�ǉ]{�P�aû�
��֜�¿4���nm�a�i��3Tj+F7���2��?n���Mi�ĺ�ԯ`e�&��R��9;����gm�\�hI�DJ�2#��%�"?
ྵ.��F,�`Y,�dv~�M�@s��f���3
�G�o��m��z:Kэ�Yrf0��*����cѲ8���JK�w:i��Zs�􏥙�hs̉-�fh�B�%����2_�`yꘕ�Ūm8J�RV�^P�2U�?q"�

��7@G��[Hp2�e��ؠ�L�6�g+��F>[��Vݳ�be>�3�[���pX�"e�\��(5�W{y��W�^>��5�k�s+�ei� hgૹ����� �U�JY"(E�I�"2TԳ/%Mx��"�<�'�4�n9�z*�޳}�6���΢����k��s��w{8��Z"��0�<_[��G���K1��}>�[�݁�dh}�z��E��M��"cS��\�����y����&���!0,�U�ӭ◷�b�XQ�T�*���R��v,�r�@0Me�����0s+��bG�F�e��y6hl��ؐ��j���S!e^�¥&����*����j!�wtK�V��8|s���&�k��.����T�'w���4-O�ˈEV��L�37A,#���Y�*�����iқ��ٱ�K;���?y�n�:�g9�z�u�i�	�A��`���$�nH�׆�t"pz |k�Lm~���"vwĮߢ�W�~(k;��XT�� Q����r,L�'Ui��g7�6=�ת�Bڜ���yȃ�� ��b ��Q�E�x��ͷ���pn��_��Vps]�\�h����G>�7e\��?�~k&_-	<ǽU�	$A=�\[�y��� ��HWms%>-��Ս��*N�8�I��P/b����u����m��Yc>`���w_�� <�3�>��s��m-v DNQv��gǆص� ��ó��>/�L��(�Mq���8w�"Z�3&�ُpe��ßƕ9kaq�&*Cw�ޙ�/!���8Vbn�Asr+�B�fi'歽4�cØ�<��ۋV�_�uсY_�����ZmճmCFA��*��<�F[�	mq-���gZ��ua	G�f�[
=�^m*f��ff�YX/͸^��M�$�ܠ��^���\*;Ln]�4��j4���1L����l�@7��Ѫ��2��v�+���ʂ0�Jq�������
�5\�9�k{�*U`�^��c���'�E��l��mjn9�{�]j���}\6�%��Y����S?�����D�WI8خM;[���q`�`l�U,����Q�$�E(m�q���2��=,)���2��V��a�Z�sg/���A���O�N���ڨv���L>y.�]j��J��T�mC2��j)ZO+�n�ᄫ]���^Z�����N�a�?��b��K��ݮ�����Οm1je��̍��[n4�s�|^M���'%�V�q��*�Z�jfޱ���p�{	빶�uMu��>G��s�:���zhԍ�F�yT!(��F�z��0!��,|͝�I���4��������\�K��n,���3>��������R�Z���� b�;>N�8�U*�5~���	"��h܅ܼxy�j� �0)�9�J�:x��N�d��o�H��H��ёX����x����C���}q��%���q�Q��E����>6 �(����Q�]�j��$��x��Ɉ�ӧ/�O�o� v��WbZ��f1v��8�9h)�WP�uc�e������٫��gۺ��c�
���2��!m�]J�@k]Ki�B{`\��|w��W��k��K6vj�H��n�5�@�>?���3��[gb��m$*�H��O�Oh0Z�TR�y-���U0�3��`i������Cq��mXM�0%s�L� ������SS+���]D��b����Ҋ����}�}1��:=�%�2r���<V�I�=�_�/�շ�g^�Ό��]��{��7
�s$)��� ,�ൢ��6t�)���5��Q���ܧ��1�g�" A]ca,����g��o)-�����pɅ�˵%�n����k��w	ô� �ȇ|�ȩ����q�2n^G�E���J�z����6�FȢ׏�*�P����6�$f26e�M�R���6�z��zt�G�O������O���{�0�i�D���k�/_��G�C�r�-��?|>���K1���ᴌvXĴŊ����ŋ)p&U�H)�xD� 3��7� mp+�ڧ/_@k��g>�X����D����Vp��p@|�;��i�#D֙���!m+W�w6�� ��P��!�+���2)it�?3��7~�WߋKc��3N2C�(xN���W��ʱba<�nAd��E��� B��G�_�6s��G���#	*��kz:p|\w"{��!��4�� ұ��%w�w+'O!h�f�3����lT�ݱPk�?�·�Ͽ����ak���"�L��w�?�i�7Y����G�
����� �޿/>�ˏG_:/�`v&siYiˑ�Y���+��h]�}D�l��.�W+��.D{�PH��s�X0_�a�Ͽ��/�?���s�Q�(�=�Q>�P�46d�e����J��2�qmf"��`�����&�z�1?����d[����[�ĺ�F6���I���A�i���9\nv���ҙ��E^"N�l�sr*�o�G����&����2�!��f�4o��v5�<䳢>)>� �]�;�O��i�z=��g@$�������;�㺏{ow?VH�w���]�~����n�M�lpwl�s���RZ�����ݝ]��\2VK /�~]C�3T0_�9-X����̹�Ǝ~\�9y�+�f�<xO|�����5�s�D�����n���V�ZE���}�Ub�o֭��-���19�O���G�1���c6�8�%��\a{r�BWd�A8�ygl�>+���J.��Y��թ�h�+0�������v��Uw�; �]�D�*�2�F�L���g��TЗ��՘^��h��r��X��� ޕ� �G���Xn[G^b�y j��X�X��ۺb��˝ф&_���K1�:s��4Y��;7��,X<��ȷ�ii�`�8{�Fg{�ؘ�����
�����K���r!���!@͸-+��Xi]Q�	,��舙��o�K����������l�rm��Ρ�8���m�Q�̕�ȅy�1(�cq��X1�6n&� և�Y�W��\�2A�G=����
	C���pRfZ-i1w!����N�7�-��jo\��鱁8z�5^<:/��kĥx��T�rb6�:��/����M�q5�8S��N/p6�s2^?:G�,���R�i���1��3X`�mp.���5�.
X�M���(S��8�O��� �u>Pk3�jK���j�f�B���ԧ�փ�kx(wG#<�Y��:���=������CC�r��J�F������<1-:_%C^���^|�#H��m���~�b�.��hk'�� �,ώ�J��z4Z"�4̑	���2j=��f-��,MF�^��}�#��)����큀oӏt����Dh�$��ik�<���\6p�l�#�$�KS�E\,��f�{0g���h�˹:���x������|5&Ѿ�Rs�.ӷ
4#�������3hջ�kr�!*U��s�^MK��Sm����{�c�ߍkP��Όū�Of�����>�@��鴤t�f����0%4�=�4�\Bt�a!���vn߼!�ڻ-�w��\��o����ǿ�gqq�/�KCdp�C�Ne��clh-����]0 ��2T��Ų��{����C��in2^z�l���42����7���	ܒ�e�h�`MS�c�6�*ņ5���J���:�
�pcu��ؿwO|���}��ޯ�������}n��\LJ�|ʰB�a{�����6~Rg��e�o��˱8=w�������=����������	-�E�k
�
,:,^��qv+@�k�*�HYkE���ۜ��i�K����܊64�����A|��ף�oJp)�P,�Aa5'�pn�X��zȞK DKo	��M�X�LK�?5@'ғv$\I/��
�r�~���`5)w�4}��(��������J�2Z��r���� *7�".���/� ��@����S���b9V�YH�/�I۱RFGFRX�
����&��3������F���ZC���{�#~�3�-��"��_X�W�8�L�ɳW��W�uh�E%^� ���l��F�n|5��=�)61�s9N�������_�`t�OFŁY�s���?��}���j�C��/�E��}kgTAa��>�d��)S��	"-����\�ȯ|���̇���/���O�8�}�Pj��'�� �H��r���g;��+��e/_�􇱱���%m9�`��u�w~��qρQZ��o}�����帴���}d��@��F;b$i2H�2'�*,�_h&����?����7>�xl^��Ο����'񓗎m�nՋi��UDfc��o6���I��,��~���1��Y�N�C!�l��������ߌ�o��8��o���3 �e}�ܣ�Օ4�0/��:�8��Q��/4\��������_�_�ml[�/�?��_��31���ԁV��N�%�t����'�nҥ��s���D��e,<ޢ����m7���Ožݛ����?����ӯG[���m[lY 0�	`kڊ������z��@&��kkP$ DT�� _�����Jw��wu�"RИ��lYS�{n��~���Ť<���p݈��$N�@c����P4�p���6�dF���i�4�>{M���&2�{�*���^�W^y��?^
wX����������$������x.~����x"����Ǐ�|.��ď�/�����W������;?z"��ē�>o~+.\:���OLMƑc��{?�Q.����s5Pw�Tj��2U
S��k��6�l��ѐ�2���:�`��4x,!<���sH����Ѥ��es�" >7�"K�KǙ��"C�l!w"�{��b����6W��%5U�����]W�����&�� 	�i9���:�A�{Em,_���� �XV��{������d�?)"�9�E�CV�wn�[Y����_�M-N�+QF��f�L�q&rW�t ��116��q��~ α�AU�H��b�F0��T�Uc���2+�뒐N���ox�
��^h�S¥%6&R�JU��o���{�s���m.�e�wn�
X%s�wh�%+xW7؞5�G���G2�`��y�/䜵P�+���D]�l�Iz�k��`cr6Ï٤!����������Dj�ֈ�γ�Q�_=g)�E���t)�b�6��I+3�Q)�72����S4�ԯ{l���0�2�ѕ��@�
�x�ͷ�#X"�Ga �r{P�����2�E��� s�]��9\�9�1�}\Ш�k��k����Ѻ�.��щQ��0U%� ��8��{KK��,~�t D0Q�ж��nR�c��꿊KW����:pozf63+f��V�sɿû�|� �8��s'q9�։�jE�U�{��U��4N��(h��ZZ䧍�����|{�'�x�!��_���v�ޮΨ"���k�0�Z��������ub��Yͧ���g�z��L��b�s�'-W8[��0ޞK)V* ���,%�����vy�5�g����tKr�:��0������uqu���N^��Z�)F�ۯ4�?�G=���.��etDq��]��f[���l6�;6fuq!�-���ٞ�O(<L[D92��I�������?AyϱR�Y�)�(��(#ԁ� M��_f֘��
�#������$Yg@�XdJ��J�R�Y�<+��,/�ak�~݆ض}���=l,���x21� Z��6+���S9:�����e�2A���n�ߟtl�wģ�`E���>�}��|�z���V�:;�<�PsT��V�d�&����.JV/۵����(�I5� �\��&ii�8��DGK��)�ܟ)�W&(�8�5�uʻ�-_���yܰY�?��+%���-Z��ə��9ۈ(�q���+�|g�P>k�&���mݳ�'J�e��:�Ǯ9GfNA�h]�����)�E��dTF��8����m]�A\���@�&�i��jA���y"�E���rL���!��y��V��Yai\a�.�Phm�\4�;����$�{F/	�<�#G��ɓ=j0T'y-�t��NG�y:��I;�P�Z�:j�|m�.ۚmhv��2&��I~l�uc6;#����f��bnl"�3#cđ����%��R�:)Z+��@Tԏ�ΆS.hi�d}z�z�:��#i)�����Y��P(�"(�Z��P�H�le%ef�H̡�7>&8�`@"ɬ�G�Hj�kb�F~��G`����VN4��D×/R)��2�¹5�3��TL�燩��h�ĳ�m����2�HLbK�������i�-!�+r;�X"�DN�nCs�utE�y3���7=}фf�{�0yۅ�Ģ\�����6�3i��2�Y�ۗcM{lX�A�Į��yc�]rw1:��]�4������_��{y~MOkT[І�4?I���eL�R����V�{9�0�Q������F�Ve@�y$�0?��	���Q��MֱҨ'E�b%��k���x�;�wĶ5��ر�*˱��q��[�mC���W`i:�8�����b�C������!-��ˎ\�n���N��zTS������1-K��Exk�fia�g���m��6"�Foy�k�i>�˵�������[^�.�ܙ���':�D�D^DJ����	^%
z�+�x+V���$�D��TFGcn
��X  �1��c_��Bή�z���Mrp�T &9i]X)D�y�n16 @�6�r�������/����H�L��5�'�Q��e?�G&��sn�AM03����5���a�ձq�,Z2��c×10�b� ����K�۹ݕ��8����u*z����m�b����rt�ע��� n��ƞ��	\5�vf��FY p�u�GsGo����U|v��u�����xH�j0�;c��ؠ�׊�-�tW��G�<�@ܳ9��X=pS|��Ɓ}�R [V�zh�N�[c2:�������|�����7�W?��X��˳�0r�X�Q�[��?�R�$�YZ�yK���d��d5c�Y����V�5�]�ӳ.>UKP�-`5-M�`OK�y�8�k}��i�=�:b��.@�;�U��������(-��@x+|�-6qg��	ttڍ���==ݸ�̿|�U��<����(��OsKrw�}��H'��k{�6���k����A,G;�uce� %h��8F�_���A>y�:许i=�A�tWWb����Z*�
�
ej���Q�gM�ۦ0�1���T��ц{�L��j��� b�'��t Ε��[�t�,'�ьb*,��Ǭ�w	�{�jw.�`��+�ǲ�򼈒V�5$r���W�P���|L3 �����rH�i0��$���J$ˋ?S�kr�6�JV���L�bݚ�شn���
3��h��K0f~�r�,]��2q�k+W0K'��2E�G	lo�10��W�8MT���vs%g�jM�N1�/���\�s�HF���v���89�?	Ky��6j�5������v�ۦp���'>������5���Ř��}�غyM���ĸt0eogK��;*M1��ٞm[����M��a��f0�@m`���u�[k�
m�U���]�֖���;@�,��T��G\Ct����5�qDg���\�j�U��%�_)����H�N]NЩR�A$t���|��
 �*7^ʕ@H��:������@� ru{�nl$\�F�.��`�u�#�8��a
{������w�[c玡X��3�z�bӆ�����q߽7Ń���sK<p���O| ���=��A��/�3X<�k.ڼ��I�N�GVg�8$�p{�"���fvrz�J�φ}y�2�d���.�u�u{�����V�������W�#�M�����R4��E�r�+YmE���52o���NT״,���2R8+XɌ��;��Ko��1A�������#�1����-������aH�_Og[<����+��P|�ǧ>�h|���_������������o�bo���-���m�sG�q���,G[;ڣ�#F�Mǈ��6�����nX��?��AIΧX�^��
��]���0� �Z���ы�o�j�3��s���?6�߈���/���c%M���ظ~M�ܺ+ek�غ>z��9�kfj׍F�,˱@: ^TG;�G̗�֬Y�`��C2����F��f������T� �[�RxDAl��YGt��J�u��q�w�v�'O��Gbl�"�`�f�-�e�-���=}�1�v(�l�k׮�q!QN�7��2&p	�
g�R����
�i �m"Z�ҙR��M�~.m�G�
XZj֭�w+5ܔ�J�ٿ#�+ � Xs:��<���m�[o?��J툊���Ŷ����q��=9>�]���5�0'h�`�8��w^4u�^�{-[���Mن��% �63��9
�^g�&-bk�*�~,�}�����%C�=ipo��I{R-����/r���Y��2`&c��\�K����3���B�S�}���8�e�߹s��ȑùN�]o��ܙvMu��;}������c�~8x����|���=��w�s_�y�=q�w���9���'�G~)��7��*i�"s� S9�ܞ�n�}v|<`b��m�&)<�x�%�,�eO�/Υ���I��4��X
���\9t2F��r�0�3'���ͭ���0�&���UL�*.�����9��ԙ�15�iWJ������zX_oo��NDK�s��:�5��{� CT����:Ù��̤5;���,���+��Ν=�sl��_�7j"�ZZ�x�NF\��)?߁U`W� ��Vy�E��������<V@��r�"��6�����zz��u�c�on߱-��Cs���v!z-�??����Yԁ2�+�����|~%��,�ĉ�ٓ��%רqm�9����l�<��n�rd�<4X�^Wp;�=�X�Js&��
Pp�	�HtkV�����:�^׋�ĵ��������oAb)�uO�s��l��
Y�:)�V�L���	e�q��[q,������}��y5Ϧ��i~��3��T�Q�Z#�\�e�{!f�qG����\m@sw�ĕ��(Uzc����ջ�J(��Gk7�H/Z�5Ξ��s���6|��ٹ��%k=0� (�Ne,�r2�������n��|��
m����^B����F�,T���R�� �:R7�Bk��꺻���S�/#���o�J���])0ZE��ݚ==�9Q���5�,�i����L�b�\OAp���?®V[BCh�,�B��To� �F~Q�P
 .kI��f5~�2 5��7�Zh�7�x#�'�q����?��Y�87d�E�3g� 6g�� ���̀�`�ҊO�{5�h:Nx�y.n��[��y N�l�%�u���r�p�.th6�~(6n� O�;b�^�p:N�<B�5x3�A}�� m/^,��z��r��Cyߌ'~�d<���T��q1-�N���0Q��B�ڻ����I�ew��*n|�o;��yZ����s�C�L�/�,�=���d7iq@&fME�N�_����kF��#{h�M�����R���U������x�D�����hF��V����\k���p�L=���f���9����`*��Dt��f@�ę�⫇�Cg�GO�WƗ�wh�3�C���à�����#G����sO��
BZ�1�ъ�����M������io�^*����p�y1���:b�ȫ%2&�-RQ���`h���_�kЫ%7�z�ŗ⅗^�l�с{�7ؗ��]
RШvV���>hl4��* 2;?y����3?�3����-L����^�[-����L3��sX0CZ#�1~Q��p�E���ZLs��c7Wc;������[s-�2�v�b��E�sV ����8f�`>�v\�
�٣dL��KP7�I)y�`0��}
Ǥ7Q�:[Mx���--]� ���:�(��2�ag���Q��&�Z\��#��oGܮ�ߵ��i��l��r�b=|$w&�����:r	'�:E�\&�1L�=��jg�&���<���7� �t��z�#����fʾ�U���V�퐮�u���ju_'6��݂`p�-x6i�9=W��Z��>*ҽ
"y�^V4�|�� �b�>G�V���;���g�~�0
���h�P޵ik.��Gr��xW������'����E���ξhA��01/#`�r[�Y�?u�t9~$�ǆ�8.]Ќ�s��d0˒� D�篐�%Lp���aw��a��0�uԿHsR���S2�#	�̵!ʁdc�-ZT>#x��*����RB[k��3�S15���M��(a�� �cgO�O^x&.`z�1�˕6�-.�	X+iY���׺+��PT8�c��]�\�T�.x$��<��a�!����r��Yk5z��j¹L���v���bZ>�0�A��A��ё˸s�Q��Uܝh-s
T�mmE7�#�P?�%��,��d�:-s`��z����?c��~vnwv$��XNٰ�®U�2y�=4_S���C�N,� ��Q+rdt��j�v��U�c5L�s(�	ܻ),
}�Uױ7.�j/��A:�n�h�O˖����3"��!�[�̏��Һ�Ź�!�(gc�Z��$�/��ko&��Nq��m�К��ʩ-�y6�A$�B
�P��S�0)c+z������x�ߩ} mG:��h���X$�
��#�:ˑ̬��s�������015��	d��hF��3'O������/Ncm���(� �>����2���?U�Y�d^@k���&n�9g���58r��0�|�ʞ�[+1s� d.Qׅ��V,�m�4Xi¬wt��4ܡ������<�G�;d�gІ<[.�:?Ǳ%�)CKK{�O��, ��0��nZ���Q?��Z�������,Uc��ڼ�_ڣ��+�e'p-.,�̤�8U,*h�T�/G���[��͠0{�׈
�@Q(��sTq��s%t��y,(��O�Ri�.�b(\#WFqM�bn�	��gJ�/�n�0�uYj���̻ �Y�3�i����p�*hk��	���-6/@S���_Yh��s��tZTu���h|U"�e�`n�r9
U���s��&�|���h�Z��K���pp;��*�����?�]�nɲ�\l�	��ƥ+#(�#����Ċ�	@|�rt��W]���.�x�e1���ś������W�����N!�-mQ"ͦj傗 5�(L k�l��Um+�"l�K�Jz���;�|,�H��nS���o�l/Uu'/mdZ�|��a�%�J�.x(���M�w��7-�m
py����'�Q~�s�K�£��д��Ks35��u?l��r4��j��E򭨨�DZ�T�~����u���8��Fù����:p�w�?w�r\<?#Sܷ=@Am�G�޾5	Ds�ip\�$߮e2>6��ҥ����E�aR<13C��(f��ڋ�r����<c�!IX �@b�����%��^�"qg�ΪmV��,�D�.κ�~1��}|q��e\�`�m� K��$.�� �wW*93�U�d�EUP2.R�v|o�X���i�֙��{W#�{N�+,&~Qw9t���z�N�bb|2'F��N�4t\X��U�.�\�c'�ơ�o�Y,�i�����\U�YY�e������}X2ݙ�[I�/��}�<Ȏ�(�cV nı�VnY)��gΈ%ZE2��=w"�X�$d����[6n�
����no-s�f��yH��Ԗ��d_���W�r]��y���GǮ�,8��1.� i'��V��q�[@ac�KR]���7�	��<�r��1�k Х :+X@=��K
,�ԗl+�	��;Jq�;�r��H�U��_��;�ۿ���w$28vg�M�Y�/����LĊIF*�bnACS�v���(���C=тQ�K-�5i��?;���OO�'b3��������Os�r\�r&.^<��/��b>�9\9����2mc��(�b.:@��4��|�;��]����5 G���J��c9c�IX�B%\W����o�ؐy��Onj���h$C�X@(f(�
����q��,${!��<W�wH�ti%q�tU�q"f��ĕK1=>~-D_O'Q���q�@ЁLQZN�����gs��y���z|��u�,�쪷KrQ�9A>(!��$�6ɬW��L����Q��Ӓ����18�O D \�."�n)���]D:R��^�}���<�WQ�o��2�\�7"K���$V���;�
�<��T4t2�=B�1��d,όG�k�b���p%�]
D�ev�J��;W��������Q�r��-������_�6�]��q��.�c���Rn��J�s c	 )żKZ���j0;�[�X�13X�6Gy�����jw4-b�PTݚVO���=UjKK�������ezb�	릕����-��:A>�2(^��N\�~�RC!�֖�.����\�JY��d ��Pt[j�i��ۍ]:�����r,��V�����g&�c��GpItw�Q�⹄��

:� svq-x%�/��J̝� �`㚯5|��9W]C�g�)�>;��ۈ����r9��ts09��gͺ�亄fh����q��.X����ڸ��@�GC18*��K縄,��y���@�>%�ܜ܁I��C����p�b��x�B��7`�B~��١ն?����0��e[(;�o Ӛw�YJ�H���z�`�(��)G:X/�F�h���X�j�˥p�W{���2�n� ��n4sO�T��i�>�ޖ{�5�ׇۀɮk[�z�RuV�+�%�d>��xO�N�У�=r\����J�l�ҝr��uQ��\�\�i����s���i<��0;A]�������F�v�\��p(a��pE�`�������觜T.&�:�e}
z��6�'06&]6�����`��,�c~o-cE��N��� ]V�grE|�!ڴ: ��ɑ����m(���
߲+��h���T�p�X��k�\1�4�zQ�7������<!8��z���]�\��F������|� �:�x���p7-���s\���[`���Oz�b��E x1�ff�����|�7;�� e�a:�4S1?=� #D\����^���`&RmM��ݺ�E>!fg��ewۗ��]�<�JZ�wZ0�۠���b,���S�*#�&�B/`�9�vvM�y�v�AG݃%�Ӱ+6���7ƞ];��bӺ�1�?֬��C�k�طk;ׇ�cu��b�!͙�K��q%��S�V�$}j�z�\�)�����F�iXT�v���C�"Q6Z���`_�ر=Ǌ��c�q�=Ļ�֛o�;n���q�q��7ǽ����sW�z��w��=̳7G��r�;�^�ޮˊ+�^�0���\��\el��ge�t�@�Hݱ��p}�&��@oç!Up��z���l�w�q[<p�}qǭw��{b��=�o��غi{l^�)�n�{wo�1���������}8���Xp��|�+R�¦5�e�鐲cf��&,�&�ؕ�.7���{,բw��6�ŚA\�lm��^`�r�Д�� �k�SO��ǹ�o55;m_
�OC��:A/B,Е����E����<�
��Z�
��ğ�@�Z2'�;�Ԯ QS�{�	
����1n���.���N��+��^��rťY�����Qk׭��k�s�k�� .D�]��M����X�����4-�D+�At<�k~�⼳/��)�-�*��[;�`� Kns01�ր[\85߅�㤗�Wh�ٮS�R���()|��㛃�}�ӛa�5ĵ�m��qc�|���i���kˍ�����;���ŝ��?�P<x��0�.��#i���p�%���[S��A٧Oe%ݭ�FXϹ��/�2�`^�3Q$.>l# \����a��g��ػg��p��#��p;�8��v�`lZ�=�n��k7���;c�� ���@��tW�[]v�ej��jv�S����}%��If�)�׌�������'ϝ���O���\��S���K��{��C��Іm�q��;b`ݶش}_l�y 6l��6�[v썝�n�=o�7�ŚZ�֮I+�
�v�eK>���C@�՝њWk�&�`}���td�!����ޖx����}8>����#���v".ft1�+��:�%5�9�ZVa����dê|)�8���E�\k��|�z������t���,�r��P  ��a����l�u����P �`�[��^�����^�KZ!��]���O��.�̿l�w�Ħr	=�f0v����������b��i�Z�P�ܾ9��7���wo�훆b���3^[�l)�r'~*,u:pg039�����1�ղ8�;������mT�.� �Y�G�6�U�[��(:�a�Z+��
"��:T�����5k����m���Z:��cm��݂��f\��v�����F6G_Oё���ɷ��ϓ���-��bE�p��@G=5&o���w5r�:QްY���)��H��8w�Q�=�}ܣ����l4lC`�M��꼔^��2�8f�ju܋pU�mG�M$K��-*y�aZ��n��^>���,��!��ƨT3j�J	,]J�%-Ǉ4���M�<2�<�R6�ۓqix,K��f��S��q��(��ͯ���9�����h��{ ���n����~i�G: 1���{a՟u��V��ll ���ԓS*�VI��u9v�؀E��v ���{�s�������T���?��k���)vT�ef8�U�(͊�B� ����YFA�ż�B�u�n�J�A�I_��SȶAv���%�7�C���V�ب&��;c%�L�p��5��
&��w�ZF�7Mh��u� 4�Van��\!�*� ��8A׮�m�vDo� ���оM%|�~rh}t"hV܎�;��{�����q�m�f��&k���V���G[�c	 �!���������獅+ #�� �f+B� ��[��γFhP��k�Tcbv�rp�p��\S��-ƅ󓀗܁p���������R��ⱸ|~6Ʈ,Ʊ���_��~�RLNa��ku�Ba�����ܮ�X@�ΏNⰵ�����ց�������~��"�Tf�2u.#�`/�.���,L_�1�eO� eê�������i/�u��`�F�
a|:������Z�킯ťK#q��0�A��=h&&��칋S����lS6�e����;[}��צ��6)�����Z�Α:|����}k �������+��A�O�9�4Ͽ�j�O�~R�`4Jm	O������WߌW^+�|��x��g��ѣq���| �����Պ�{>���x��Qʈ%��>;=Inq�(�;(�u�Kj.�*��`�F�w�c�lFVZ��3�>��rg|蓟�������������_���k~<n�����c�lt���+��H���m�	�ܻ���lC�!-T�6:���R>[�#̠�;� .�gۈ�,�� �B���z���<���ګo���T�g_>��?�K�dSz��5�Xm���̢��yO�\��-��Dl�pHu;�wPQ����tS�G�;��,���O���f��t'���r������[ ��@��Mz*����i��)�����A��?N�:_��I5�q^}����������[��g_��7HP�\�=�NJ%�B 	�9v��mp� jma�Mr������W>�K��7���S���/ġ��%�/���e�C�[���|�hh���XG~[`���+Qks�v\�}�q�n�	�]�I�v��G>��x�����G�����ġcЖ}��AL�@��-%�`��5��5逻64Yw%��q��x�g���Ɇ��%�e���<0.�hM8q���]�ͮu6J���Ή�\f��D{���o�����c��[o���9���'�/��5E.jX/�V� �S.�=|ڳ۸�D���%��k���!V�5��鏼�t1~��P/��>��G�F����ɵCk���j��ɍ�J���m����a�F����(��Z��)śG��104�����~��m ~_�.A�rG��M]CY�1-�W�������~���<��x>~��sс�\�aS���]���ޞh��ɸ8v%.�\�'��i<���q��4߂�ZSXLsШF}L���2����Q�n'_CC�I��^����ݔ��]��-#{[���w>�H��ԝ3U��� m��m45͓j"	A�ry8�-tqx2�<z����Hf l���4}�	�{�?�`�$��ցP�gy;-�d���M�50I����q�С(�;:�	�o�{��O���	wȟ�	��������澍�ήn~c2C�I����^�Y���-;r�W&bl>���b|���ċh�%,�S{�#�NCHs�� n�L����SJ�N�Cm'R�E�5��6s�q�ⅸx�|NV����.�3���)�yq*'9�ufv"'�/L��Fg��`�%*Y�s}V�hy�NFz��_��f��~��|鍷0?{�\­ ��H�\�h>����}��M�h޷�A�+Ywo�ʕx�����^ÚX�5����h_��.��G�řӧ��}��܅s�v�ٳ��'c�����NA����e�zt��,w;��Y�+WF㍷���o>ԟ��G�yr�S�F���R�A�����<�#����f��x+��8}�x����~�^��#	���q<u�8�t"�/�ϡ��ԛ#t�T��%�+��7zz��Q��/����3� ��1:�$5�a��'g����U1ʶ-���U�V�x<vo�O<�t|��߉������Ͻ�k�Fkʬ#��T��=�w���Ė��Q����N��(*\�ʬL,a�_���U�=#L�h�ԍ`�׎m�6��;n���vh�u������S�B4]�(���L��8y�J�z�DL`�
"����e�j�f���̱��1��<�l�ʫ9���y>\s]��N}�ԉ8|�H.e�Y�*�lfb*A�����	��/����2��72'��viZ?q*^��*��7m�3�/��rG�g1[��<���B'�
�P]D�O�BH�\t�9=��Pu"BT�D\��y"���G�˗�������N�X�r>���o������Wa:��i^ƒC���(�����ɘ�n>ג�gG��o���] \�щ��D�e�������,�r4c=B�L���Auv�c����hԋ.`�O���C ��Ụ�: K�g�Úu�18���1��p�?Ag`�?�
� ���Y�oܜ��a��oSq�̙8w�bL�w��§I.�]��3�كֆFwׁt#u�P�Y�cv��`���<+1i5ֆ���%��݈4ph��\6�wa1�DoO�DG�!��w&=�P
N�t{��pq9\�zaq%F��)G��	�+��דg�Zt��ab�H(���x܋�}˺���O��W���㸅�/ŉc'�ɟ�?�w_��Ϟ�Bz�ww���7߄+G�tp���LYG'�ɂ"z2���k��� ����nM�(AG�_ikA	��;��.@��8����;k���[��""SMK�?����ű8r
T��ՕQ;�B�4,�bViA-q��zm%���sU�v�ٓ�{� ����<ϴ�4�+R-�}������	��+�a��@�B�{}�?[���9<2GА���f�|�A~�Ģ��&���V}+氽)�� �=E�j>�ϵ��&{�R�e�.y1�k�+"-4M�a��jK\�|6�`���R�jGk�?�+��;7�к�ؾ}s�~�p�m���	w�\"o��atUC�}0�J����4tl/z��ciF�b6�\$؉\F�n��X��t$������2�g�֖�i�c2u&��M֣����m۶�'?���{�-��������g����w��8�|J*���D��u�jd���8E��c�U�k�Ñ~7�P����y�Zw)q�~,��@��%�x��̞{:��Ӌ�Lk�q-S.D�]{枻o�����F4������nE8�;�]�t)Aa�����m {�d�plj&�9mö��"sxț=*��'��@sd&�/ƍvR����Q�^3V��C�]6t>3<����u��g/�ŕ��k	��y�ضcK����8r� ����D��r�Qw�^E�N��^\�r r�-�����`~��e��lo!���L
���.\�9�D%.�N�����=�*@B%i�
"6��%��["H�n
2s��\w�j+��B�"�:����z��u7}���&b��ٸp��ܹ��r�T\:�鉩|7�em��K.�5�n݆t�9�3i���*����5���e<�,�Q�ȲI �-�/S�%�
5�"�D��s�28�����`v@�.z�����u�Y�!����G>7�|�3�xs��s#B�.nع7��>�k0��O+��<���ڥ vbJO�a-��s)]<#��Q���6'Z��Z	z��r0�6�29`�y���
�c�z�Lk�x����,���{������8u�l�]��:o�g�}�v��%\E�b���A��Z"h�%�m4V�u#��2�m W�q�n{�!G��-�VW�i�"�~lTwv��{z��HZ�q6��ɐ����Y��hq�v>�< Yt(�������'qhV��wf/���MX�S|c�:���^�2 !m�&�h� Byey-�ޕS,,O�����{wo��^=��9��+�lԦ&EN�O�\_�a|_:t<~��!�8q�J��4��{x���M��$��: ҈^m�%��t D�t�}���ζ�����A{1C�.���Y�F�}6�6����(H�H_��3�n#*CE��-��#���+���#ΦY��j�����+���������2�:�5r������:31;��+�89�[b���<��CiG.�G�c8�#a���K;�ֆ�&���'YaR��R�}q�Y�h!�'����)����C��P�Zkk�cf������SO>Oeu" ���w~�����#�lޕL�f7"b���t>�eq����ZR��GXj �2�%���m5��f��5H]�����N;o�����e�<`�,S��c9a/���/.�Ң4��B_���⯾���_��W���v���?�^|9��8}�v$��.�=��K�|�URr�\��*����οqPz�q�rcw�>�'Pv�F-�D�aq	�*'����SƲ��r��F�έ��M츜{]�9�y^�O�ޝ��|����B�3I@l�;��+���-	ii��f��mZ�"�)fIw����SVD<��\���1��G����E�]�v�|�-�ř��x��J|�''��z)NS/=�����R��A@���roT����)�9Ta2���w�bz���atd,\�J���Iܙ1:�PQNn�=v-*('8�완[X"֫��P�;&��!�C�[b�{a���Il���N�R�$��p,�\�}����t&�@?�%�Z�]���
hӨ�<7���k�o��R��h��M�
�O-�S��$8�������$�"�Qzp��:rK���̘���S
D��I�B:+�o�/��C3�&+��B銑+�����n�<q<ۋN�8_��7���|�5N�?'N'-h�	�ލ�� :T㦭1��l7�]��E�܄�F�ep5��C�2ZE�(um��-W]C�QF!:񱶠U� *�E�]��ARk�Q���Oa{�]~p7���7�ܱC171�ϟ�3�;M��1�Uh�4�T�T�^,�F�����h�]�B��>�PpѹU����	�d�}����\P�V��\(�K\���7�+i�j�Hr�x�3�5��\K�\$iи�;���Htv��Se,Ⱦ�༳�/v����š7�²rmޕذ~Ж�� -j�S�א���W����~�P1[@::���`m(��g��8o���3��;��Kyu�9A��"e�T]lKz��!ovm�v����Dg;/R�d� ����3IW�7���HwFyp[�k�a�'�ywt:H.{rH[�&MH���p����"�ZȠEa�kZ�L�LF���x[�^�"M��9�x�;j wyC�!(B��'5I��no�\is_!.a5`}��sfy>�`�T7h��Eu��mm��T���M
�ݷMmh0''�M��K'��!�$ x�B��9׬ ˕��{�z{p��&�;�f���[�oҎ��a���x�W����f��\�x1�{�x��O
ch��x�W��B7��Vv���92��1�f w�7�o�[AQa6�_n� ��Y~D���U ��GL4y��hͱ0G�,�,�+<Iy��� ���
s�8W~s��
V�⦽���=��[n�{�+���twa��k��޵���;�Yw��U>�jUA���l�iW�ۢ��.Q�ʉ��͊ 3�
���D�H�t��%.DUh�V��}-�[�qY�L��C���?�9���w�/�����o|7�|�ٸB�6n�pl�hy�_ ,\.��
V�=�!2��(�֊)x��(V!ϱ����5�.�x�Ƿ������@�Fa�s~):�'�q\H��>ma�Æ�y;:(�*n�V�!Wr������er����z�����r��|��r�����6ҥ,K �|oc�=b�ܠ�)�%4�4�]rU�k�������f�?|���'����*�Q�t� ���_�ͦ(_�]h�JH��Tp#�R�tp����R���2ͬ��gͣ.v�Z�M�Vy��XM���uBѥK~2��<i@̶2�_��)��e��
w�K��z5\������늇y8�����M7�7�rK|�?���'b���9���.씿��+6m�}}}9^!g�B�L������t�k���BQW?���oC���2�
�]H�tM2-J(�\�^T��3�?��������ۿ�����������o���E������رktT�����h\='N�o��B��kz��_� �m�i��j� [�O�F��|_�Í�a���%��(w�̑�ZP
�̳Xپ��"�sXFS��S9���28���u��x�����P���q�=��֭�c��dT�����v�Y���� �m��Ts�6�/9�A���M_ŭZׄ��I�����Tt]J��A~�k�؍�q?�@��Br>�~9�A+ɮ�E���X@I���%��0��z�[hȱ��y6UX���AfZ8��t�+��gs�0�m�BÖ(�/B
�	���kF6���.�)���"����|@/�J#[�;�(�W4u��,R��d,���JH�"+Â�G��>6�PL��KT���x�ώ���_u��	���Ey}g�Ʊ~nY� U�N ����2��.��U���y����_�\������| n��ָ�^����?{ߣyM?��8�OY���6���Sԙ�9Iqjp��LQd�z���_�Yzߐ�Z��%��q�ȫc(l�qM
��(lp�R�Ar��-�����g/\���;�/�տ��/�E���'p׺{�r���1,Lc	 ����^�����j�<�-�� ,ۣ��i�c��z�%�ha)s��nRh��\�!�O��iZ ��v`���6��L���lZ��X��<�t|�_˅�m��R
��G�y����/|!�;=��ۻ}�i��-٫s��l�_3Е>��f�V�n�Y]$�0A��,�nta�V:r,� J)�&���F}�F�CVf�iq���vs��o�:p�z%�*-X(0,�% ����9^j�� ����P0��v��A~򺲟����J1��"�1hNf�ha�	%B�,�D�����+�������b�����5�9����qg6_F��o$�yϿ��s.�<��و
�	+�$,M3L4�ė(ٵ�����6�]Cެ��ɗ���N�''�aB;x~���B�k�$Z�c�ơؽ�,�R���������{?�~�u�-���Xhb��5MZ�����!@
Q	��ֆ���Q�(,���P�b�O����l���|��
{��Z"Z���$;s��Y]&�}k��4���Z�6:�;�� ��4���&(@��ZQ=Dgsw ]h�jO.m9�)WQw�5w{�������l�̫Kv[@���-'-L�xav8��+U��l������g�������V���a��?�g�������~?��O�]<������N�pI�M�ŭ7�8 NB����j��R�'�� '6���}�"�Z�*b���n����a���o�����ǯ}�bۺ,��pC�J��8��>�A�B,�����h[��C�ط}M�:����n|�?��"���3��G�n/\v�d8J7�5�3/7L1�����T�y�4>>�=s~%3���%[l!����n�dc#iiZ���'  ��IDATݩj)n��T������PKtw"e���r̍G��\�i<�ה��ҿ��������s���qy|6�'�b݆m\+����Õ�sJ��  �����JbWCq��H�O�m�P������"#xEMh7�݈��ZR�_��C��s���O!�ݽ�cǮ���p��Z�,~�#i��]o�")��955�W.Ü��5�0�j��s@��BG�\hX�Y�F�-��M�����&s�&�[N-��3��2?��2������}1�v(��ͽp��3gO�SO=��������+�YW�o�3XW����!ͱ h�����Ȳω\���]�e���8����%�'���f�}�$�-13=�;˹�BE`�\��Y @쿬M�JW�p�[�����>��7Hy����;�5���L7��T��v�MWt۶m(��TP�c|̲�}6	@x����"�����.�U��޼�+n;�;y������;n��vm���ؖs,����(�rT��ea"zHf��޸i϶���?���uS����lOK��?��|]p���2�^@N����y�	��}���ھh`�r�:����-_�sT�p{��4<�9U���o�"8r=�w��פa�Bc\D`�E*W���_��L����A(ȥhA0`̍}�щ�ZzrB�
�K�Y)�n��*����[l�i�-�v���8r�Z|�:�Ғx�_��(\D���I��/��片H��,�ϢQ:�T����)�$.�cc�&��z٨�qn�����B<� �[����C�ꫯ����;R����+:�Y{���ZŦ�C���e1yu'/�V4~�|ș���w��<+���3j7��˱}��t	\�I�֡�e�Ľr�⚥-XzsX���+���k�œO=E9^�ӧO��F�K�:�_G�:Q"M�H�m::���{��m�+��.#�|�f{Ԩ'*¼�/���Ɣ{b���o��TF�J(#��/�z���➻n���i<'�-� |��D-P/�1 �=���ƃ>��zk�t��q���8x�MqӍIk%W.s|��b;����b���ы�56z��{�3����3hp-lAD���9^�6;�-eZ����;7�o����ч�6B����	��={w�M7�C����ĕ�}�@��=w�'>�H��M���)�����Pt1"� �_Ͽdl��|��fuc�U;�#�[w�Z�k�v�3nٳ��E�1�����80
"j��Ӵ��l����'��_��7��I��6t�z����;v�e)���W��0IW��mD�;�LY����]�lmOlA�Z�Z7_nS[Vb�H7���}t�Ɯ�D���sZE��E��1�{ ��(��NM�����w%�e�eNP��2�"!ٯ=�9�.3D�i��9��y��;b��1r�RLNͧ�����em�b1����#[ ���#*��_ʮBӞB@m�u�v�m���ށtFGGr�O���m�����
�v���"�6�tmHz�
�c,\��G�������.&��n�W.��Iv�m�G{olپ=N��zz��W�n��;0����2 ���n��������7���C��8��r�rK9�_{�dz��]_6{�a�v���p�*�& [������W~��qǭҪ:{�DnåZ��.��݉�ՙu�z�S3Siu8����3����M�~����n��A��%�����;n�-֯]���t�����P� ڝ��^��rʓ4_A���������O=�T<��+q�̥|�����/źuC��~��b�޽�����?�vn��J9~��k��N�q�4� �TH�Q�ֵ�-u���5]��*�W�i��_��/�m���)�� �ȫ�l����՝I�Ct?������1�5(��C���U�-5�m�D�Т�DK��h*�Q�tL�)�Z0}fj2�>>������E����d�sz��=��pʘ���
��S "�J}N��Fs{�`�,7;8�M��.^��������\<��Gs�۩S�r����d`j	�e��B�~���4���<�/�6����+����������ޤ��R6c
�ｏǍ�o&߭X`��i󖜩��޷oO�
�O�[q������B:�z��}���8�ow|�C���M���~��Ũ��P�z6=�i#�Wo��fے[61�ܿ+>���ġ7_ý:�V�mf�e"�'w�v{<��#q��?��s�9���ؾu[T+'�;� >t81���bhiy:;c����#!{�܅�x��bA��(hv�7z�deƁ�hz�!���'O��2vu�ŧ?�h>ϟ$������.���������o�/�/��e~3�?~�h���-&<��{�y�V�_�_z9^{����-�7f��7���D���bPZ�|�\a-�6�U��uA�~���cז��ɓO�׾�-��r�u�l��kb��`����j,Ŏ�|S��щ�x�c�o�(��ݧ��+����m�M�A~(�B�e���9N��Z,�����ђu-ם���=��nW��ye@w�t
��l&�`��hCkv�PaZ�4��Ǉ�md�y%\/[��ϥ�5~�n�l}���=  q~��Bw�z06����K1�{���i<�3��5	�̂���K�X:��W��p�M����<v�&���O������ܱ�tO���[ZLP����ӌ��Y6+]��+ &3@������Ł��I6�[�yy-z7;��a���3�9.���w����F��n�s��}({�1�x ��]��AV�]xjM��fZ�����4ݲq]����yf���"����w
�S�q;8߶eK�ޱ=��ߝ����"�onC���{bl$�{���ڗ�?����<�>�t��}�p'"X�
����5ہ�ٷ�7��f,�N��:pXx$.x6�<����?���2�h���f������"�Ԉ.������%�
��\���}m�pR��ub���������89�{��"|&�����s���+#�/�ﴼ��L��Y�g�^ �;^�C�,��Vc�ڍ(����2#�&Q����m���g�_�N���1ҭ���5�=��d���b��������^�SW�b��K\���uQ��2}���TɞW蕲��{�<c��:�r�k{f	"׆d0��P�����4��C~��L��6 �~�F>q��ʼ���.t|^�gh�+}�b�X�͢��ShVԈ:�+���a���,<��ua\@\d􄝨$*�|�?�Ĵi���G�첄aj��0�e#� ��%���ZY��<���eK���B�A���g�@��)/0:�����k�sQb �
Ck1�\���=_��_������7���w�q���s�w��_x�9�t�>�O7(�=��D(��fL��̟:X`7�|�j��.2����(�N�DX F�ϴ���i�;j�1/�ϭ���o�7��ո�&��p���8���_�y���+����~���=��:)Q�]XT_���Z�`���J�E�2�Qv2�#Q��F	T�l4xְK\\>�U��� \"���3�W��Fb�֘,l�uۏb�������Z�N�49�{�$ٱsW�e�����vX�4O�Q{7�y&��S6�ߕ�c Y�[�g�Fy.aU��:pߪq��8���pk��=z:��O�B�B<��Kq��e�!��ҕ=��Xi��,,B#��~AH~��ʲ�z�?y4x͞�%x:W7k�MCy�"�QAoX"�����
[�C���V�WO&���̜ɀE��h��Tx(�@��O�����+C��r�a�iޝ"�C�y\�Zs�-��jk� *3X%�5�Q9�jJ*��ŭ)�5�؄�9��J>`V�9S����u!�#�KyB�Qs�Q�,��e�,0EҦ����Tq�rJ2 �b�0�`_Ot#��Ϟ��}�Kq�������;�q���x��'⅟>�=�T������tו�:LZ�m����Z/�WBC�� jM&.�ixg���w��3��`�ٟj'!IGt��u-���� ��X�\9��]e�i]H���T���'0�Ǐ�I�Kс{* ɜj��7�59\C����-�OP滹#�Y������Q�q��Mr�����@�P�v�Pm�Ӣ�>���jW����(�X�j���L�����t���<t�{z��0���}�18�6���I����6�S��J�F_�h�ن��.�{�@�z:���U�e��޶2[����m[h�&g╗_��|�X'�b�-�ھ��P�Q��)\�*�m�)���/��l��U�^�mmX**���׀H���^M[OH�$4���
&����:�m�M!�?�3�Aϴ�(ZT��Ta��<�8��y(U���Mch�X�}[lۿ?v��xk�$n�wcl�|��رw_���u��]�16f���tD���hB����*�D�"��.���t�AKQ�Zb6��x	�ZM���6Щ��/_�m AnG[��v��n��[6���C�rE���w���#���w֭�������?�������,������5ϛ��TV�7����DRef����}З��!�(8�#GQ$A
$�!	��A{WU]&�dVVz�����־罗Y�݄�}�~���Z���v�/�O�ԧ��d�����3�S
G�ldC�T�������N^9��n��l���	b�r{?�4�uDɵM�0�+^5&0��;gΜ�Tt����3��}�=y�2}�3\?�����p����ţ���?�t�W�\���� ��\�73�I:gH�qԥs��-��СE�>m�i�#TL�S��'@�!����ׅoPY����51�1u5�>����׏ć>���l<���q��sq
�;O��wf�O��?�lL�I P��!�8ʦvӆ�,�pyG���U�q�ɺ�UJ����O���}���/��G����9>���i��R�sgNħ����ُ�g_x<�9=Ϟ��<u0�O��-ߤ����`:ZKs�y�y�s��ʬq�5�5r^q�F�v牤v �[������@�V K��;7bja�FC���ګ���LU�7�G)l#::S��K�.�&��p@b4�Μ<O�?�tو�7�������8{�d|���#��GO�?�=#���b����qb,:�O��Ө���i�z��]��/��훨�#�x������h\�r=���@�k����E��"ͳ<g]%�	���ZަQS��@$l���ȉ��Ь��r���4��t=v� r4�s@�?�عx��s��T<�>�	�ȣ����N�7r�����q4��9�'M����ߌ�޺k.�3�:�s�.����H�<j4���O��O�K	y��W���I���%�o�<z�,D�x<��y��x��3O?Od�N�O������mNǙG�Ɓ����>L�u��h4���a��~�W޼�}��� X6Ј6W�bӴ�U��6AyC��!�ҡj�E`�}�}O���K�nN��n����-�`v>����sߐ�GuF?��=���>���x;~,��eg�ݩ�1D�R0�<q<N=������_��gJ����FKi�m�V�� �������4��Z�!4��Ν�O~��Źx��jQ���;8�z?J۟��;�?~,^x�t|���K����.�<<�F*�r��<�>��K�.t\F�a�I;��ڱ�V�T>e��`���%9Ձ΋ᘎ���`�t9O�+{�e-�wn�K9��܅w{B�Uf2#���7��h�����avtm9�V` ?'�UG���r;f��Wa�MPy|b?��Y�=���y�F��U�~�=�#�URs`,���c�g8�ƎǉG���J�s8rtt8����z8y�}.���Ju���+إ6�~�ǔ���~X\��~�l��w5&��2���R�t�H΍��u��_cSUw?�n����������2Ə�0�A����N��R���a41L�-�؅VSwwDLsh��d�j���l�I[pwp��o�u吢ҏ�8���=/32l�V�ң
���I����Ð54�nLO��S�o6G	�Ȥ&���3Oőc���10q8zǣgh_4'�Fm�P4FC#��<�Ѥl5�6���ĝ��0ݝ�WG���&LYk�D�)�=����Lv���B��_��6�z&p� .M?G)M���o/g�b;�X�{�y�OޛC��
�u�b����b�Бh"��P�ǁ��1R-[UPO2�3T� ���7��6�d�^wv��6hW�[�C�!_��.����Kqq�?��'c�яơ�>�����ӱ�us~"�7�c�w,��ǭ�cѽ���;�t��P�<��h�L�u ���/� F�+��i��$Ss
z\eul�)�S6��Z�k˄� ���f�3���q"U��ɵ*� �i�${�i��8�'�-�<_�\��G��f}0(�H@ ǥ� �6��u�K؆�D�ҚY�;�&Bb[�� x���v'����Ѱk{"��2�.B�[�q��@	��R=�,r�Q��1��7��A>zz����T�\F���$2Q��0��EZ�<t�P�uj�4�]��Y�=���r73*�]�0��<���0��z�z�Q����"�Q����j[0��09�����@	�����
u���䃣�1�kn�U`�T�쥽s�1�
|�	�)םrz�\J�a�E�2�!0?t�r�@��89L�r꘍C��Ȃ�]^˽xgW7c���YƍXnuǲ�į�r��K0�%��M�30������xl��P����Hl;��ϧ��f�ӎ4`�ݲ�w�ĩ��	4�T�~@�|e���r{;� ���!�c��h���
�l��v���u��Ϫ.�ב�k9����`sށ��'ݹnn&��[h~��K�5)s�ȿ�%�i�9
�
�U4����V����ߊ��?�j�Ͽ���g����_�^������������K���ߋ��_�Q����������������_���o|!��������ߍ�߉�y���F�:j��5�K���{\u)�&���@d!ۦ��k�T�d`�P8CT	ٙU�xU�>l��@��z�ƣ4aD-��QH�U���=3b|&h_�f���WO��k�Td��i4���j;�0�+�B���ڹW�y+���B�u�j��2��--��O���m�Z��;��׃;�-.-���9�a��V�Ί�.�Q�3�y�S��xߥ\jpڐn�ﻚR�w���^"_�x�,nG�}�Yz�����ׯ����X^p7��q��[���o���α��}fΝ�zj6�ҟ�{�@�;�鸒WN�@��yT�U2Z_�M�6����s��p�����++�q��x���x�������)�;��u��͸���;W���1y�NN��}�V\�z3w?��rζ昙Jo9�k�X��v��W^����]P�W?��I�뢺U����ګoťKWi�٘�Y��7���.�ŷߍw(û���u�g0�R>��\��V���[��:¡+�N��0o�*�w@�g���':��w��>���&R�v޽|%��կ��|�����������o8������������/�����o������wⷿ���/~=~��_�����}�������!PF<?�v�#����/���NpiuyYZ�I��:Y���%L�����X�P�J<2��m�@�S".H�y�f^ 1@i<w+��&'�%��p�W~	?�܊ּ�x���p�c�I���6Dy7����C�p�^��u;���)�#̫���G_α{��tWlAġ_�<�1�3��� �.�O�x�'�S�r,���a��=<���y�
�(	�=�J��������K/�K/� ޸p!��t�{���^�
3�S^�x1nݸ�.����7�K_��x���.[��,� ӳ��������h��5J^���\vv�%�Ҳ��s�����!�A�̏(��~��⥋�"eq���c����c-�R�Ʃ��0�߹u��ݻ�q��$� P}��������e;�8읉�u�vB{��*��8�)� ��c|܍��g���Nϙ�ܑ�/���Ñ4�L�����M@ϭB��!����K�.�ۗ/���B8|4&0o��j1I�/���H�^��@�vx̾�D�m=;W��FF�s�C�=C],C?�����b�cn������E�Xꬍ9�a+hLj���s��WbE��#����!.i�C#=x������K�_�f��O:�%W�~�n��͌HƷ�]#a��y&�z�s�s�rl$f�43�s07�1�p��Uj�p�hzw�v��i6�_s$�yn���;o��kW.�[o�o�y!�����ݻq����/C�/�l���AR�;�34 jk�`:|8:��)ä0��M��u�N���Њ�*_��o���Z*����cq��I�C��t֝ڈ����w�����~5~��KF�>�d|�}��?�||�S�'?�9aP��S�0�O�PWK+��Ƥi�h�sP0~�c�ޛ玫�l�l3'�yL�o��h@� ����]�]��nw~�_�p�`�q�Fvߑ���pG�����7>����}c�w����خ7�c���q��d.����A�M�	�r���r{�x�WQ ���w˕���s�_�sϖ;���m��w9�H<������s9�|tl8G������=�_Cc#�a<�Vcrz)���o��	�s3�	L��M��� ��^5��.`xO����v�ǰ
 ��;Ll���,��hZ�?n��nm�H���
ڏ_��{O��Xp�iR��.#GG+����[`���v`��H�ڡ4\�v:/D��D_#(Ҁ�;L���lh �\d��	c�/�@�@O�o���\	*�M譼z�9���#iƴ�XU��c���6�ko���Ƶ�����Ӽ�,�\~�j5�K����Cغ0�j�q��qڀ�;�XUZ��R����t>ӗ y�*z��A��Rq� 	D"��ؗ+nU���e`��k �g�޺��?y��ƌ���vr��8�C�����N��u{�#e��𴑛O:�����R�p��-�����=�R���Ka�y� �M�h��_�;5_���*c0�S�G9���6��6+���as6��ƣm`�.�imf�`@<H����V�W��G�R4�mZ~��2余��#�~�EA�Ƴ��B�rx�~L������$�d�{b �?J���$496G������R+޽��6��60�g�A��~�oӣ���jMyF�$G[ 5�칚}�
z�����a�w�{T$1� hԠ�K
Ν.!�� v�_t����[V�C]�޺.<�dT ��[�)�}	��+Z���w���I��;���!��BB��	��-�6KE�&jF�8r�a��-c$�i�Z��eG��}���؍���H��p�1A��D><��h�}9��+(�����l���qN���h00���� �م*�4�4�v�m��J��Kge�*��ڳ2��&�\_�[��;ޯ�937O��Ɖ���є�i�
�������̙3�%�͛K�1�Y���]ZΣG� ���N�sHQs�:s^Bi����f����pU�
@v��AfU2���v<�m�k	�\+�5���\�Ei�F�M�1I���e�~��]״�������m�k5z�H�fo�jQ������"��{��X�S[K�#}V����{^���{�\%+�x,��"}��O
`Qkt��`-�' ��uQ c�5��~F�9+��^�o�Me_���RL�P�ˏ��}�����S2�/͗�>sN���!���u`AC�)ϡO��{���
%J���& �>.��h'.Ju�W:�ڍ�<�%���JWtm��VSs���t�� gY��G���/�d����	�/��>MP�V&Tm�-6�HI|\��&˛�L%�P@3Bx�}����x̵��~��)���W�>��#���駟���M�<y�l.>�L�ՖN�t��8� �)����μ�i� *(&��ƙ32i�cu�b�\2�e�e@u�ԝ��_�r��i�����~������Tݷo�>}&Μ=1����G��s�?�}���a"�HMg��4n�~�ޯcK�:�����̖*n�lz��w|�)ad4�S�oa<�Z����D� �����p�ʯ��s	N����Q�i[?k�����Ӷ���PS��������gY�3�ؔ�T�N�q�y ӕ����`�g��7qD��܂��7i���##��u~D��� �٬Ob�-z�h�}ٯ2>>#;g�NM����4�v���M�����vY�C��
��	i[��}^E���'w�WXg{�f\����/���ބ\MK��m�9�W4_���::�haI�p�$"���y�T�.��3OK�z	�U}gp>@J�F���ҫ(�tl���Q́8hP���C��T����Y��ɘ$3T-ns��;~U3,_�� �4u��@bښ2��#G�IG���e�~~Q),j���V-!��5�ʉZ��/8a�J��H���`e�(�ŚKb�2���{Vh�Rᔙ�U��/��}`����w���;�����"�;E��� r���8v�8�:�?AU�����?�����5��:L0s�����y�	���PBX�>��u_�~g�5Q*¨|^w�[���tF�4���3��l�����zsf|b4�eR3@
����_B!��[�Ø-�� H+H:C�}kZ�gG���Vj�����3�<vn��p>�</�)��j6�F�If���b6�_��ԩq� �p3���P�T�-L>���p;y�4��tΰ���;�j�h7�"�RH:�\*�3���疊������Q�c��1��JY$�[�J0���Ʌ�*{N�̎r*`p�@�؋�/����au�u&����']Q��4��5쒰>�nn�I^=p���q�x��W�k�8ܛ�ƀK$"B�:��n�H�<�dʰ�HU��\`(�i�֖s�����1:��0"9r����|8���ko�k���;]Qo��?4���hQ8����܍[��MUΜ=�ڋ����T�fú�L.,CBZY�o��a�:�M��ܰ0�k��$���0�;w�틗ca��\7Z�!��;$m�Y�7�&��2�q`̹/���mB�h&N���;p$Ν{
��W_��_�_[%n��L	>w?�;Q�}\�m�{�� �o��C�\�FS��	��Jo���3�R�2]���&K�J5���A�:0�,δ�F���1K������^j��R�(���e�>��c�Y��iU�^� a��8���3�2���j�_0������3�� ����qDj�6�1x��Ն k��1�>���S�=��w��q���v.�k��w~�K ���P~�&��ӡ'�.`Q.ӕR��Qb�4�i�����9y��c��6��x~��Zȵ?��38`�4b?Ω<�O*������{H���a5US�W�6D�)%$��B\0�1��$4����LoS���T� �Ŵq%f+7�AZ9o��:��ݳoߺ� ���w����d'$���о��D����'���g8�ǩ��0������ǎR&���p�F�gTe�HΉ������jJ��E�y� U���m^�Bu�U��BM�)4����p/AL��L�Ch~����a�&ZF}`I=�`��, s0[7Z�#�>G��,_�C��0����Dk�Tt�AQc�`���9�[��އ���A�ܑ�Z�/#s�K0Ow�N������~7���oǛ��ay5�7�|;^}���t�J�����h�	��I� ܄@����<R�EBh{1�+5�e�w�\9J�G��jF�W�R�h �:���Ņ�K��}4R�&�`?z�x<x����hև��&٢.��C#�〢��ǵXn�����K�}f�f�xwV��c>+��_J��xʱ,44r맀�炈�}^֣�B�t�N]H�;���΃��\�D{���Q*J[�).A$��{�ㆄ_�=�J��ۓ��Y&Ϩr�G2��e��^.��C�<&�����B������Yi��H������1D�P���0��d��W����$L׈}�I�C&��8�{s9q�Y��ھ}=��"��v.�SeU��2��o�PK��p��:���Ob�iL�_��5�4��������ߌ+�n��h.��y)޺|-޽y7�ߙ�k�&����q���C?��~��P9�q�2�M�mMUwM'�^b�����Aއ�C_����I�o N{��4	���K~ JI܇�[Y���;��7/ ,߉^���IT��X^�î�Pb�)��R�Իb��!g�MM��Y=;��S۩�U��t!|��ny��< 0�����TQkv�����en~:VV���i�q������Iz���x뭋���~?�	@���9)�ƻWb���h����,t����$G5"��W5:��rE4�^����`~"v�g���f9��L�J9�Dz����N?�Q�Yw�+�-�K�[�;AD���,:Nm�T1;�O확��Q:����%:	��H�$�D����UU���ڻq�=�~���/�ېv�Y�M��Q��_}5���{��׹�o]z;����2�7=���2w����K�㏿���h��t�
D("o@P�,��Y�"+Y���vOw�U�����^�'�$�W�X�q��C�ֹ�.�~�ߌo�����+������b|���?x��x`y���W߈�1�. ,/��z����A|��_�4Z8���V��cq��AL���pViJ9�R��u���uJ{�'G��"0�rNG�:�#5j#n�<3;�Z���G�đ}1>�Yۍ�tMH��	и}�j�����6~��#ͮ8st,>��9@�������4�J~J�=�����RyTH�\��4���֍f���A��z��S�y"�{��Ջq�15u3��o��^��|� Ƿ�⥷r6��^�	�/���_��~�= c0Ν=Ǐ��G?�l|���:�>�"�}�{�܏��W�6g�p/8��Q)�{=���2�cS�N����=��\i�%��O�q�ǭ����i�J�����~TZd��p�@��������9[��Y�k���}�������+�����w]� ������wq/k�Kɥ	c��-@�J�� �{[�7��_����l4c)V��������o�T�������b���H����5����q�ut��Z9�Z�3=0�2�e*nܼ�\������˿��?��觡���o����ø>�[�#�J� 2V��V6����:ꢫ[-�㹕G)�I^�FIc����d��/�T��������fL޼���o��7��"�q4�f���A�/��+�����m���3I��3s�^^��qwV�k�W�>CuU�F|��ߍ����qs�~�~��$�{���$�Kb���z;��/�_����F���ML�۱�<�l ��l{۹Fw���ۘ=� Q"��ܳ�\`/�c���Lo=q*zF���0����'�����&��_޴]�\i�u��R����N�J�Ȥ����(�t#O����ę����r�bO�-! ���w��O�/,R��ӣ�[v��s�nC�u�׸�{� �%In.��0�7k�cW40E��^����w޽���_�;7&c-2��0���4#��:�źrZ�Z���Z����ouh�4�n���R�p�9����u��׹񒥵ݲ�T�L����S�8i@�J2 O9�ώ�N�����-7j~����k�:>���1}�8�Q^�,4�I@L�8x	O:sӳ�*v{����������gc���Tp�s}C��>�7?��-����+�8tI�G�DG�t������g����cȫ�����V��Ϣ270S���`k[0�*iP1f���`��L�������V�m�<9��c�Ň>��8|d4�[0��w���	@Fs$V6��dި�N�s�
"�0Jx>'�|�j"D��u�4��
�_�������
��}���q~k׸�V�:��iչd�)��-�U�l5�/�՝8Ľ驩ZuI��'��
����;���������n��-�(�xH�
@[@��8V��%��/���ü��󟋿�7�r��c����GD��ssS�����jc���\�g�h��k�M�)�XJ7qv�hku+�w�]L8�5�����^����Qt��-0��p�>&=9��6J��8���I�v�m�XDKz����_���N<��Y�k��v��ɍ�攪�SVvݓ�#.�>��A���v��#9���Ȳz���}\z�_����?�څ�������y�=V1Ź�i'����>n�ljGw���\%O��5�H�,Bf��0q�6@}5�#�4��z���+u^Z���p�UD��aZyUe`�"��mB�h���9�����>r.&��G��������Xq��U{LF���^��+�l_\����_�A\�>۵~4�@�V�PJ��<f��h������Q������Ï,��������+>��'�;�ksf�n�W�#.L�3c�-�ț�R�T��!z�ǝ���Ý�rf,�63=��ݴy ���	߈����������bz����b��Re��H�0cJ�MʅL�A\�-�R6�D"W�
�n%���?�S���?��1��޷9�-ln"nB���v�Cy2X���sں�`0?�U��� �}ڀx];Sw.M����V�5�|W������I|���Tk������W]��-V�33l��o�Y�~�����P�OQ�ԍyr�&��Խs{�HՆ��\MZ�Om��ʷ����i"�]�\Mle�6��Gӹ���.�Esh^J����I2�khqm8���*�F0�ј�0;~�>>�d�	#C0 y�s�����O��䨟C�gQ;��⛴�uҬ$��PL�wSHaв�[�tZB�ܑ?���W��u@�����R!��D�#q~�\�T�٩M;��b q��m=A9p��h�kT�+�y��mz�2p:������"��jk�'-'j�����r,���=�ch���_�����Ͽ/�����к���|��DdA�d��,/��k��BE����R�����x��)�0�[#���L���q���:	�<�I�p�*C�T?�(������|R�/�'?�hhNwa�3���e~
a��N\io�u����ˀ�Ά�����}V�����%�����������4먷��C��+{�SA��d�	Kf�@�<�/�<�����B��t���ѯ�s�>�__3on�����Zm�Aݵ�%������V���6jjD���fڊ�ex��aR@�"<7��#̳�/�M����hVI�z\���� ��>��`篓��#�ı#��`dx0��#�%�m��յP�U�˩�����%T#�b�釯����?�f��wF�}_3s3��q�bJ�qT��$|Aļ:�YS�o�~5�$�$=�0ۇ�Ψ]x�ǎ���TaTG �cD�rv��Y��>g��&mY��.��5�߸=��d0.]���t�͹;��j���qs;�eJ�����[�f}��3������%͡�t�N�?�ˊ��5��'��ſ�3��/|���Z�O����46�2A�hLB��#�_�5 �����O~�K���[�30�{+��K� aW��N�=�I,�������ktOK{���*>q�L|���C�@�z<���C��A���8b�b�����Ry���8����!$����+�D���΁�����w��Q��026;V~�)s���Rz�1�r%�[�/"�2K���d0?��׷���>}"��~r�9¸ʵ�,[b��ȏ��$�Es݋��6��)�͌�s'xG@���H��܍����q�N\�q7��>�m/����1��c�u�+���&u����I'�����������i��^OG�6�)	��8ɂ��W ��#�8�ZfB[�n�8�ڊe�������}�B�����X��F��JgY}$Y~�ɻt�����*t�%%;��4�n4]A�3QA��d~��g��/�+ �Ѧ-n�{-'K�#M������X/s,ʂE�$'Z*"	4�'Hŀf,u7���[�i�ޟ'��N�J��qs�SG��o��O�O�tԶ]�N���>��h�$!�^���K����F���G���oF�;?��b"-����������
������x�qTO�82�
�M4I�����TrJwc��{��V�
ƨ	��o��.;|�6�P]����t��Ъ����aY2�s602���d �+Y� H��o�2�$�XG6RV���/�eݙ;T?��}jy�O�m�S��'Bs{�f� vm+�rO\��P)�GJ˾���@�޾�K���p�Ju��7\V���8	��n�-��%#�������5��Kʭ+
䞪<ȶK���
&�y����`%a7��	�9/�lI?��y�� ��>��K ԕ��jל	ʵ�L�ytـ�ݙ��}�\���%� �1khi� @�fҀ<q�v���N�e4��Fo�$�4b	zXGve���j�9z�D5��]�_�}g�z4^��Ԯ�2Z�.h8o*���'~��I�0����߼���/Ad�^q�ډ�c���!>���hh&����tH	������F���YOV�Ae�b���+�;Nb��#�K`_�
�sr���?i�����w fh`���J���R�+�1=���K���ۗ���XG#Y���߷{�Y׻bjv�t�D��Bؿ}�]��jCQG��!u!I$��̯u��a�u6�'�ت�PBJ6˥�ZTUK�|
p֣{���N��FG����cpp�rאxĶ��E�Ⱦ�#lws8�}�#o$B}h�T�O���HLL���C18@Y�^�1���cxx��f��e���TC�y�W�Q��Dj�F�emq�I�ՂP��i�e�)u��i��˶h5a0gI��$�!�h�jV���j2~�E�C���=��N�$^�=i�44,�#$�0�C�2C7fT7͢��'�r.�c�n�vʵ-0��u4�^!�`�5ap�f�A�]���ȹ#~J^�hΑ�Yq^K�ugǖy(�g�ýj��@�ٝB�G8�1>�[�����u�&���i�����+��i�fk���/a
�pU�]g�q B;�T��i������g6Bz���W�[�0mu���< B�q��5}H�\�J�Èj���0�v����$���2��s���	>�%1B�J8u}��P3�4���rj�����E��HfmD�@)M� ֋����sV�����@ـ��Vmz;��K>�z��]�e��Ǻe��{-�N9�S��)�ki��6pnH��Jݮcq�xW;��ƃ�sA60E}�ڪ!=f����:&C�������Y�h��,��������M���H!����CR���X�SU��]���VK����r�ƺ�`������~����1j�S�1?7�u��6��׹]�G :��wL�Q-2�q#ڮ�Fs��6[�9�C�)�罛k����l��l�'!�_���^͖�X��#��V;�Ej>�h,�5a�6w�F`U�H�{�+�v/�Z��>�����*�(J�~5�\��ʝsSf����H�ɼ�Kޡ ,����s�C)WaNF�g��Ky�w2Rb�s����~�n�ˑ����izNWc!-��"V�
���\���l ��M`r��6�� �;9W+��^{�FC�t���6|k�|;Ř�H@)ő�;�x�}���c%�.5ٹ�I���h1���Ĕ;������H7���]�pn�M4ġ�O}s�E8O	�tpH� tĢ��Cn�����<���K�� �m�y���u5���׸�Q�Nlk�,*5���pd��y�@s�ۿ��ۇ���<���=E�K�p�%���GZ�uV�%�xr8�m�w����t�����s�h���_�-Ǻ4A3��y�\(4�܏����F����c��<�h�������<�K�#��.έrt��H�Ƒ��˧^��gg��L[򟶫��c��:�'����;�w�KZ#L���ᯄ��N����*I����t��|�$M���l�1����&�sV� ��u3f� ��Y'�Y\� ���q�ZV��N��i;��P����@�z+�o� ���<��Q��\�w����eĩ�)(���9�LP�I��ƻ�����+x�[X�=m|��Sk�rz�A5>;RuHWj�����Uy5�4�.$fA$��ɛ���kN�L�/��[NS��|;�[���wy���M�U�,���hi&�*h���w�����kM�2EE�u�#�q�⨖;�
�Wy�w_�����E��M�e�a��ۇ��׌-�c��4� ��@xo��ͺ��#S�B�W3�@�֢	�Ƿ�W(Xf���O_ �/ 
�<`�X�ɩ�6���*��}z ���֨�-�X����m��>(���D7Ν$h���r"�-��.�gO �Mm��5h.W��N�d�d��6H��t�N`Hb,.��y�,�-|�q�;���?ܹj_�����(Q�Q�kjV9�*I��0�@���P%d`�(Sl�P4��Tg��.{�����+e0v�3ŵ�������WJ4J� ��^C_))`���Ӆ��$��C��ڎ޲�R��ε(�SF�F.C��|qy�Y26G�d 6=�`5��/�D�T��5S��B�eR���pJ=�m���<�m�^JG�j	�,ѓ�U�N�ޗ�}��������6H{��0�`�}Qz�Q&$��`'��P�^8�/��_aj�NA�DHM���o�cn#�7֝,��~��z)��K=:T��Zʎ�M̃-��CjJĝ���Xy��i[A�2��^/ �P>}���=y�I���_<�$H��N~t��4�/u�i�g�T����7��B$=ȴ~,��._yG� <�ʛ�"���f~��t��Z�y�s�G��{�O�J�tH;*X���s���.5�̟�S�{P�zJ�\��4��T^5M]VN�=�%�@肆�J��6�$��:��+���$(�4\�9�O�a,
+����NP��d��v@��<<zm��#�X&��8
ce$%a��ҟ2��J12l2���샨���\�d��y"��	p�V��9��`,G��BB�ap򨹯���2�f�S$��y�D,�%`T&���s~��h�)��!nK\z��"Lat}���;����^�2��"�����JgCiM2���FQ��-`���5m[hG�O�y�Wv�;�6���t���1U1�g�O�l_'��-t�t�j �����G�2���z4�p�z�^,h;����py��4B�����<�s��ʹ������+��2j�RfẠ�B�0�~]���+O�8@���eӾ��N.9{֝�d�L�����{+/+������l8��LT�Jz�F����`�r%b	�"���
��	8�NR
���s�'MTs���g�)= �t�HIo�@Dͭ I���S���=��� �H���|_-�㜀�����7Y`�e%��G� ^��6i9Iю'?y$�j��ם�uI�����������<yqd�5P9s�Eo=t���CUs�]?X��u� ��#��1?���{mlչE}n�E_�@��]�vmPG�F���"�'4���}�ڝTv��^i2�O5���� �s��]P�^x�9.n����k�6}�>������w��&f�zg���/��ͨ�ҡ���)q�(�=<���K�JM/�ś��<@��" #ʮ��;���9ۋ,:wx��%8��|����)ے��0�C��@�~oC)��%��p瞙"�
�^���<�Y��SmU2*9��8�*����c�k�$�2���ݠ�M��,y����;a2W�Av�f��j�D�!�� k0���v�J���ؗJy�$�~ `�y$�mY�]��@Q��H�5���^��ZPiÀ0*�W-������7<��K��y��JsK�����9����s�%�s��Rv@B;�-Y����
D��9y7��!l�9�Rv�ժRG�n���	"{=ռ$���w<�W���	v`�8�C� ��:ڨH��~�s�>,)�0>�K�!�h�X���`S���%���Tw 4�6�T��Ro��p�B��v,�x��ɓ��35��/�2�f0�X�Z��l��a�`�t��A�"�G*PLnla����Dum��_�ڋ�׮��2��v&?�c��_��R�ś��zm�y�+U|N��^��觡��
�wn���*R
�]=Muhl���$js�=��˰�� �d�ћ+����,�TI1�h�n�����F�>�ecs/UGN���ZzA���;�p]
��6�)<	���ǆ���%�$~����l  ֑�F���q�5dǁ�.HkQ�͜��'���q�5]o���HL6jE�J�4���P%K��Tw�L��r^��A.Kc�����}Y^�~��<��
��{�T����;��NX%Y	F�i��n�g[�������8y^�Z%��j�
��=J�.��
R86�!���=�D�y.ۇ*�����i���^Y �[��Z�QZ�=���d�$��9Z�Ћ���l�N��0jYū�䴅u@�+Ȼ_�Y���x�)ڿf�n�(� Ů�P�:�� -I��O�Gx�6Jo��o��ͦԔ��ͭk�~�P݌S���?�럍�?w,�j0e��vs����H&�A����dv���2ܛ�ޝ�����������t�0H��d��J!xs����r,]676y*�B6��z-��ގ�奜�����������J�\|'##��H�!����< 2���	K°�ə�<��r+]���G����<*���֑,Ys�3��u>@��:��G��@��Օ�]j��}4�ǽ>�0��f�&!�Κ��`����IM���B�o�i�%3@�lM��O|&H�ˬ{��uQ@$�\�&d��
q	P�ԕ���1㧽2.�2��P�O��_��.W��Ir���:t��6��g<�C�������U�w9�}���7O�:8�QF��*���I�;mέ���@ͩ�ul���8����"S�5�L�r�9;�����k�
=ڼ�rbX���CWZ��Ѕ 5H�����I�Q4V��:
U���Dȯ�R)�q�)Ϩs�fڶh��
D�g��|m�NjXû ��$�8}|_������S�c�o�L�Ib�����K�$R}����+tU��%R��vsQ܎'tً��X��s+�23�(*Iu�q&|��Z��v�_@���SW̚�KE��5���1���9�wN�< %^�!�NqJMW�*�þ[�&���8�у~�fR�r�V��u�R�km	-���D�@� l7b"�DZ,����X���z��u�M�٠N��> �mm;&zע����=��oo��S�� 9 ��z3��j�����/kW�?�I�471?7�IBC�c��4�ը�o�m`]��V�5L������\�{�G�����I8��O6��f�{�GO�:�yiwC���.�9�ކ+�{x�;��6��K\z�7��s��� O������F��'>�&޸Lc+�r���<A�~�}m�j���l�i��\C��X�vu�@;����^*} |7�c{!Z�S��:�A���]�~@|�:!ή��/�㻷�?]��Z�2���I�К�$p�4�QMH	еS�Ѓ�N]h&
I�3�4/0�P��� X'�K��=ΗKx���Yj����S���	��z��|��*)r�9�{0���Py����t����������p����s�.oV��W;��AgUݓO=�DQ*��Px^��Ap�{%�ϭ�l�ĳL��'墄��`>�Ew��s�iF�9�JZ�����$)�ű�OA�&7���}E��	����P�F�����N������������B`DU��˯���K�xH��� ƗC����q�Z/}%��!k}5`���	����}�����F��u�Jtw(�o&�qR��Nc��@��ʔ�s,���S���+D�;�$E�Z�q
m��VctƬ����+RI*�#|��@e�t��2��ک�u��P�NL*Y�s.�+��ۑ ��in�D��ܹ2h�Q:,\��@G�x��C�/gwm��/��+f`��D��g�%��]�+^�,LV��y��
LJb����x�׹��\Ta+W�F9x���8�V�����O�y/��zpJX��S��sq޷��� ⨖���Nxo��
l!���4�iɛ���뱰Ҏ���u2)���]8�,�{{<ɑ4\���@�6���Y8-MXD�ߠ�kaP���{�x<z�ɗ�N��1�2�.���권դ��82LE���,�4O� ���?C ��^�r�?�:��`r�����C���3�s W�S�n����Q��
,��#�mi�
��呔�U��)��R� �<Hr$�rS���췩h��̓�/��L��_�������Ny�8͛��W%��1��eAw]ň3Z����,��g�����j�䞨v�~O@�y]���2���]�u��x�+9�)~��y�!��)���r��w� ֕��v�J��؏!Q(�b�M�Z반ahv0��;�Ҋ����[n%��fAfT(r>�{z������#6��#��BGԊw.�{��bˉ�' �W�\�j\�7�SSډ��"�S��|��>w��w��yOS|VD�a5�$h[*�[�D ��53�٩� �;�ae�����^����� ��vpH�N9���H���R�
6E��Q�p�}i	K��HRt�羂O�Xw'�VjyE�\D*8�ق*��
Zҟu���.P�.�7.׃eĔC�:�zͺ�X����@b>~�+|N�䍳�\§�s^@����R�����mU�[�F�1�P��Y�{3���4��7��z��q;u���y���>7v�.5��˻q�U�˨�W�����)3�N���)�����*ոH;��u�94[�^i$)�n�����5��3n}'!i�d����>���'qe��7/����*�o�JD%���ar^I��c�Oǧ:��N����^�QB�9/�{�Y��R��Г���+�lC��eH���'�O>��Ƴ3�D��[%e��!��k��Ip~�é��C
Q5��Y�?�Nq �gGe�ޣ�5���S"*����{ �*�p��'�閜�SZ�²����Ⲙ<�0^X������ȏq����+8-����_�����"��@�Xm{7��uɠI0y	Q�0z��o��I���F�罊qK{�w��\s�\�|�����I�9��}O�3���;ci�j�U	_�3��\��r�2;���e���^N�"R7h��t����ʽFG�����C18�/���w�";��&.�,8b���zW��Z2C���u��a�i�당 C���y��xj���Dn���7���}-����qm���H�x�gʪ��N���ԍN8�;�]�9���[��\>��e<e�~�3�����?��.�2���&ǯ,-�:Z����X�v�R�k��\#`T��򞾀��ib����2GTn���C��Q���3ٮ�������{��r�qT����+A/�U�д��۹��v�s]��������D��2���[[q\I'��TO�R%fz�<O�u����t��{]�{���g��Q *2+�;y���Nd��{�uy_�)�:�K�; �SE:���}@�^>�3�Y��}$��(Gڱ�s������T.{wS�>�l,`�k��c#�0G�W�Ʊ��IO\2�OF.�\G�9OBf&M��g=0@��W��]M��Q��=z���&���k��L^3�)�Z�9�q�~�4<��97�V��� �݄!TN�#�)�s]��\�R����}x�\�0��������<v��r�!m7��F@������dh���z1y@*�t�v�s�џ��h0=qg1�jz���Q�\�M���f5�79�		r���
4ww�>rF���! �Mz���岜��;�qT�������+��ϒy�'���-�pH�W�^Z\���x+[[1�����|5�{�zl�6�n4�n]#�;;Y�W�'�9��X'��6�p3뵸u�rt��U4�M2M����?<����:��x]��2�L�DqG���b���j^�J�^{}��M��|=���b-��>�x���l��c;��NnJ��`��qF�j�$~�?���OP�W>5g�	 ]���F�k�>��H&�i��s��������,I~'����p�;�����!��\��{���ک�*���y��f޹��`r2���[�;�vs���Y��k��a��6mzB��<T������r韣,d���5�����^[]u�a�6�s�&�Վ��� ��Ņ��[��V���r$�]������y"���3G�*W�#Ғf���D�kR�,YO
��@��|ƌt�A�v�=y ��_z!~��� ���B|_r�ũ�AE��ƕ��L��ŷ.Fk�'��7�7����7nq'l�X���O"i����f#'�ݹ�.��A�5"�Vu; ���э?͸:��s�; ��/���u}�d����������ά�v��F�%Ztι�
�> ~�LN[�iF���Z�C�U�]g�~9���I^� Rq�wۦ:��N
IT�e���8�v�������f��e�;���$kjh��*=O;��<J���|x+A�<�}��h���\�]"5G�u��&pZ���&�Dzw�_�,X1��SP��-�I�vc` � ���#U���񓝰"	Vf�y�<D\��6�ZZ�������q治껙t}h~�G�<8d�(W��( ɚ)N�v-�ODvR�2��:5���;�� ����E �ԟ�U�Y%Z�u�Tƃ\���)�zZ@���qt�,�������~��B�I�f�{�̣�ڭ4�C�66uiޝ�W�?��p7���������ܤ3WA��.�F�DC屜�;���F��ثm�Z\��oG����������T� ���R���<���~������&��ă�&�n<��G�'��a8V&�ǾN^�sM��rܹ��5�;�r��@�nQ[v�RRVՖ2��յ��4�ܙ�.@���eL�f? 2��;��I�6R ��$�K펕�_�v ѻ1f>$$�g�d��Ã�n~��c�{�O�=�[SųP�L�,�̭�s�,�Y����Z]����A��;�z�/�Q��������ϒ���8ْ�q�̆��=a�0���Y�䏰*$�H�%a��cuiM�!B7,���^��EC�O���9t�9OO��d��5C;����0��[u��Q,��;U?�s���3�C�n�{5�\-��QŨOG[̆ݎ��@'�S�����o둒ɴv����E֑�Ov�CH�/���?� =FE ��}���<M���ќ0���sR�}!�` ��-�]4eA�O������"f�jj����ܛ��v�����lYtr��fҞ��\���~�.iJw?�������:.�K]�����@�+@��E<�������s��P$���Bs�~jK%|�i�B��$��W�g>3?�l��W��Qe~�լB4~�E�h�4m�=J�d�����+;�Y��\y�^�CX;�=�g=g�m�sߎ�ܕ�r�x����{�v���-σ}��W���8e�w9��<wL��I-9����=x�W��v��3-��:p�F��9/�u^�Vn��0��^�z^E��G9r'�z� 	�]$Ѧ)C�*�u���HD\:uW�"�J1橔������<���t'�t�-O�?|�Y��}�O��2vDq�sh1��磒A�*]2��gu%���$ �ۛ~2�L�K��ݸ�������1!6�W. 9�ŵ��E�{�B����B��,�
-�$c�a��A�`����^&< �<��pm<���'�-77»^#wJïSU�sN��x5�ߍF �so��A���T�{��5I)�Z�ˢ��{��O=��^����c�A��Q�Th���Q����Pd���<�|~��{�{�V{�����,_�I	9���A!K��t�-�2!�$~�qS3��n�O`��7*�=�c��&�K��I�E�w���tY�mZc:Nm��Wz�3���������B�?�"FN��2L��l <C��[]0K�y�>���j�_�v����v����v>��i�x��;a���`ִ%|�XWj:�� �Ԡܔ#O�	�4!4����ݼ|s��M;l:���rU�%��4[�[���E�[�;B�y����#�eb<y�s�����-���^��c�!e�r��y�����]��~d�������g�e�c�h^:GU�^����}�6=׫{=�݂f�#�a~F\tp�ŽV�1@��In��z��^�m�B�%H�{�28�A4�ޏ�K�)H8Q��݋���Yh�uf�re��F���NȄ�-�A�ù��N�u��ȹ���q��sH*u�C�B�^:��� ]u���y&w�!X��B'?��*>����;�<7�z{3^{��XZێ��k��_��3YV�v�`��JC���N�N�2Y��
s����ܹ��]F��+�3���P��2Γ�&����خ���,s����T�������h����K6i�1� �`WrY\�٪�<�����&��;;Ϊ��zQa�!o���d�gk��}+�8�ù	�ZS;\W��j���-Gvj����1��8���&�v�Db�����p����2������:id�$:��y̱�Yu��+$�+�t>+��y���{�*�}�����*���if=״��Bƍ�椵�������͗.����y̓<��U����+��>/v�����$��q�)/:�������ccy9i�`���j������Ʌ��	-�E��=�3�N[誼�v�p\�B�uL��a^S�Ż[�m��j��o�ǫܫ��=8�>?��3�4,�KR�|'�� ��g����b���[4P_\�\�����kW�����wQ_�mQ��?5��l�/{Y���"�f�RAd�Yzd�^D�b�aTI��F��ܤ�m�o������e���@�"�:Ao�8$�TU�"hD? R6j��-;�mf�;[ӑ�w-/����`�z�)�d:��R�w+��RM'N�q�ͅ� l�&�m��ͬ�rx����A�2漋,+a2���QW��k�yw'·��[�t�lO��Ѯ�����_��+q�I�"O�`���d<F��s���d:HVy��:�'�'�y��en���W�|�?"�z�z��\Y���э��}��,��J�~^�}F�&q횻��sx�d#�Y���{��s87�I����=@A����ȑ������?�h���3~�Y2����ϲ�qٙ�ɠ�m&��e@�a�����}�Y���F�e���SqJ�R��>��8��V��C\�+����'N%ȏ�ҏtvRc6��F <W�VD����_���OY��ɰ��ޏ���sD $@R��Cr(q�m�Y�=�D���[<s��m|��w���}JT��w�}e?���@w<���$�e��������s�^��[�5�_�p�kh��\�u��Ƨ+ =��]3t�߀���e9��kws/���o���sW�LM�r�9��rF�C�
T�Z�CANS5�%H_�k���!HܓWڒ�͑�I0�K�i�J��� +�t�9�%���A^'My.��n�?JS�N�v�d���l�KMs$�)���o�ެ:�������
�Y�Q�&Y(�����;��T��n'�N��g?�= ��ʪ��O�J�wΩG�W걀H�Ѥ�P��8��L���L�����NY�a	��4��F#��U6��xg��Phv��u��<�����5~�OQ�$����{η7wÿ��l�������C�a<��9����NQog/�`2�� _��{�$�u�a�z�X۹�E�v�5|��<zE��>ڸ �uȱ�PQ��(�K�'gh�]����-[��h�:������
y�\~3>;��dv�j�n���%�E^��b��
YG���ǽWѨ���h �ʀ���e�u�<|�Km;��̺ /���Q��.�S���o'���
h�9���N��{x��r��p�};�H4)<�|e.�/����={W��1ê�0ʷw �z#jNfQ^YǼ��\�׃�v�P�����9w��sGT��� �L���D0Ԯw�K�չ��VP�W~�{{��g�y���ǽ�����2o���'�*���v���Ս���y�s�G�j�yy�i������k&��q��lO�P-D�	tN��c]3��	�͡vª��췓UѾ�@�K��Ds��ɸ�H:���ޡ��u��/彼�Əp����ԩE�Z�j��tFj>}�f,j!�b�#5;@=C31Ov��Y\��T�{��a��{+F��ū��וg����*����iF;��.��w�Od7n;�<�3�N�2-nxЎ�S���j�C���Hd�9���8"�R}��m�z0�>w.�x	__�Pb�?^s�8�4.��d��k�W��SS���y�z�����IU��%��qT��ܩ�l��v�^�Q��R������i��~N>��܍ε���I����ғ��B� w<|��H&�W��4u����u d��ʙ�9C�#���D��� @88YM�47y�j���Rh�߆��:iM�2���X�C]&g�P&Ԋ��۷o������Cf����g���{8�]���qd#��G�R�t�~��~���CV����.o�N/!'#z�S���,�����uU�g����=��?su�摕�+�r�%�Ļ�]y�z��߼�9�@��L[u
H;�u��[�_³cՎf�hS,�xj���K�q<����#� ���xޓ�r�9�\=�<����N�����Kϯ���_w/ Ts��kp�xHSAW��(�˵�ZM+�r˹��V_W/� �����x��t���X����C�}V�9"�T�k�W����B�ML� DpX̗�=[�k��5�CC�@8���o�	�Kk�0i��BFp>(>i����7��<��U�K�B�y׮�������*A'HDtf���/sE�BMF���5	$���XtJ��VVix���7�*>�;8�����" ѕ{�Iś���J����;�:ad�JjU�2n��;U�:O�q�����v��;E�A���ʮ���]���0T����qg�[�)�Z3��6}1.��;7Iu�7�9�*H�$(R:�[!��-�=�5�������`������U���W���*L'����8�]��ͻ�@�}�#j��~��솉��]����4���!JO�X?x��}��<wu�dp����}�rt���8�w��1���YW����o�n�8��Q�OR�=i��M4Z�4(&~s���s�����t���Ғ��FA�I��3@�`��|H^���&:/5���J���vh�
W��I��U4� �y�M×_M�$W��ߚ�s���c��С��֕'���.#&���J�������q2gUP_��P~o{NK�ݴ�������w�|O���[O%����A:�8�\�$�u~y�#\�����lf�3�0�w�.�FQ�!����7�aw�7�*?�`� q(sZ�b�7 ��F-�����i�������w|�<��!���c��5��o�9w
����G�=D��	�`O�-�[��K<����͒rs#�#=��9Z�e��]����)��]��[�����y�!H�{��s�ۉC�<�%�cav&V��`4�n?J���7F�pB���AM�f����<ރJ���	�W*3�CM�*>��v�U�b��3�9��R'ݩ@H�>�C�~�v����q�/���(�I�K+�ƅ7����]X����/�K��`�A�=���;)�����a�Dd�����j�<�M�y"Υ�F�A7@~'ጡ39O�������s�H�Pt��{�?%�9����$���y"�+��27Gc��V@O���.��[VHq�gU�ge��'�v����Y����Rl�'Fǐb���!�?��;�7�l -�a�i�����%w��7|a}O�?� ��r��Hv�I|9��:P�k~������	�htBn�HX5��$SH�[:��"Ko[��L� `y����zʰ�w��c�U���N»7'��~�*����@�I:��۝���%�|w\u_3* ���{�g:c����8K��*�i�+at�Iz��i?�ۘ[>��� Z��]��0{ch8�gO�PR�g�:�p��R��<x�ɋ���m8)���o5O�D����s+��2�k�N6�������y*�g'c~n&N�=�d��� B�Y��m��.����_�����Z\�����/�u�K�燦r�Y�y�(}+���SW/j��t�Z���j�+S'@�ՙ@��H�J~GE�v����}�X= 6�U@d�� ��i��W�[�ry�g��w���p^����s������T:Nݾk��E����6���N��Tp�\'��G�H�0W�BfC"�D qMF�F+6�+i�j[2a�s��v�͵��fS�τ����q�,�ɋr�/�1-}�<��A�'��{C;�*���^1oE�+ڟO�kjl<SC�����Xʓ�!�;˘����)q��W�����
�\`�C�3d�ꧨ��h �	����҄�_֚�Th��щ�����\����	���6��u כ��BiD�d�Z_#�'���ey�;����_�X��g�����X���G�?��;�tO-��^�G�7��b�**g��䃋���5�+��J�f�p>+1e�9ͭ�(���K�������.�~��������:���s�N��bǽ7佮"ƪ�Ɲ��i�t��_�>ʑ�p�=�^��1�Ƚ�5n3�=�uQ���FK�c��ڈǞ����X�>���I�CM����w�ף��x�W�|B��k4a��~��ו��������?�#	9>����>��*��]O~�s�3g-wg�]�2jr��Ǿ�hy;G�s,�������(<O~��٬��q�'w����K�~>��=�2��8�L�*j����:����v ���=�`����_t;tͯ����eX��S ��1�#3>�����U~���]2�I���U�Z ��<�U@ �lX���+�{O\��N�w��uy�ײ��=��ӧ�c\��-��Wy^���c'~�{��q�pje9�N��2�H:@b
Y���(�O�%h(}��J�Q���|��mHG\"��8�+w�"��}�� ���7io���_��W�8n�)�v�_���/����S��N�Xͭț�
Sy�-�ü�״�s��L��a^�O��E��\�(���u����ۥ���o<����僽��~/���W��GaL/A��몭m�Cܾ����=���0�fj���e8�j�Pǳ�$�4T�~���|±���o.��ʪ(a
�J�Z��u���s�D|���He][g�� D)$���'���gH�W�zN�6����f���I!��x܍�3¨��InE�����f�e�G<;+��f���Ɵ���S��ᘒ���`����g�:�2u��|�W����;K���޲�)�x�8���,+_��R�4ǥ���A�@d��_�:��2�%�W�@�����Fä��4�;Y��h�?�*�e���Q�N}�|���v Ʊ��c�y���r����X�V;@I&H�_>{���^`�~���>�d���)
��:3���R�W�+Gw�7oN����\9����T���S	xI�h���B�[Hhk ��%��>Lg�o��e?&����Z�v2�Л�4�M�+�� ����Z��3��Uq C%���XB�$� G�R�I�M�ɲdy��Fm�]������L�иc����1�x6�<5C=�B��۵��e�P�jm�g��Yi��f���mT�\HG<~�߉:��6iY	9����ؼ(�:�{
��c���I�����RY��i�s�`��J�dx�m ��2*T$�%W��В
��X����-jc���K���4!�[P�,a��ǜuf�RIQ�&D�& ���׺���g�m�oR�����z�p7����h����-w;���zl��	�zk�)@o��,���Td6c��ȩe�T~˗�N�._�'m��E�kځ�� G�����U'��m,���J�i��ԗ_��$��bZ�h �H���靈�Z������[&�+���\���5���"�6q�����|��y���M~[�,�g��!�$-Ң,�K���ıޢ<�U���G��=`��j������s��ܜ�Ay@����b�Tw�=Wi!|�4�"<��:ys��[A��&��/��%J���j�xߵoQ�tɄ��M�#M�C�[=�ǔ���L~�~{y�N�B��b��������9|��WuF����f�nA�-��
,����0l~��P�a�*Tz�-L	��J%��V��\8��ɀXʹ�s�#yHwǓfAY�e�6��gG*}l�J�	E�Z���a�Պ܊���_�N��v)�� V�f@f�F�Re$�X�+{mv)j��O�#���j�׃��G@��z�0i���H��H� fko���`-qq�圈�U�Z&�KhYK��^��6�m��@�j���s��Kѳ1#M��(u�t� )@ֿ�ՙeH�C����ߏFws�~�=�is@Y�fm3��wu����x���un[�2�*�訃�I�΁X��W4H�a��<��ĽD�s���礗��37.���({�`���8���=S�=㖺rR��)��l�����ı� lS���"�:�ZTs��m�F��x�G}d8��a�*�δy�=gK	��-W��"�S8�����j�»���}��1S�/Z��.wQ8��ժK
�S�u���`qi�/�<�<���]���D,��2޼p!�����ٹ�W�b�|q66zi��hԕ
�:Z�	q�
���Ց�RII�=ѕ�o�31��m�=J��cqr*��9�R%��j�	�l�"��"����)b�����}k����󰺮4�q��\FLD��<;`��}k�k��XE��G�ͷ���ڬ�5�P!�'(uwob'���zc �v1�FlR~�Ш�F_�� �s˩X�Q�i��R�X�.9�Qf�:���G�R������o��m�FHwq6��ގ�e�`�l�-B�};�r����#9c�C����V�:6�A�;�_����ζɅ��\C�p�H~&AO�S_�o�
�R��Q.M���2�$0��`�{,v��ו0�)MF��;7�w�ѫ�Xc�,C��~/ߩ���	�;��\�����U]��4	h�@k.{z��R���;��#g��x�����#q-7�r&lNP�o}jg��*YJ�j��2�b�����F���=�ޯ|�g+�h�~`Lk�Q����!����1��w� ��w_��]��5	�;��vBAe�� c+Xj�U�E�H>3��&,� ���c�[��gf�4Oz* Rh�R�E 0A��ş<[YC E_{!��x[N� �`Ӊ>0}�Jn�g�u�P0���#)@���S0;���e$�.������1��5�>4�>L��fo<��q�ȱX�[����n;VPW�����ā���o����j�5�������/��DWq��nL��6�@�O?v.���� �b�zr�]>:z�P�<q8��{)~�_��w0�6��J$������o�l������f�L�F�Z�.��-��&�ۈ��������k�1�ba��p�������-�6/Ry����}%-i��dV��cy���ZS��<��9鐚Q�$�6�X��"�wʒ^��9w{�F�K�����{�o��B�j�]A��-�x�2����N�*��i�)���nxz>p*�eN�ư��� ��) R��� B� ��4�׿���_���1XC[E	X���Y���3�T_f%=��Z{=�ܾ�	����ɸr{ICs݃��6�O-�zj����/=�,��&�Z0Y;q2%�vJ������͒4QxװnRk���h	v��kv�u�s�d�̥��$v�yC���ޞ���> X�B�OQCM�M$�&連phj��$t�sF'@��~��?r�P��/~>>��g���p鏓��c����;�������ތ7�xM`�x,��Q��4��8T�*!���f�b;~�/�g>���7X�>̰S�'���`�8<|�|<����?֌+߈�w5AkY����0�Te�?q9�-��8�S����P�p_@����5��3�� �L�@;�9k���C���w�H:�	�6��hǡĠ6r�w	��\h����� ��ٝ9ܣa;>����2O{Bo2SjiޓΌs��s�ɘz�SP�!����N})�k|/u������~	�u�4df[a�W����΃�Ti�`ˏ�e�T�v��F�cߞ�f���d���}D��E���>���B�m�h�5�}�w�aS7�D�ͮX]Y�I�b���8�z�N\�9����^@��ܴCNd0���2��w�X�H5�//�_N}��7�=�ވ��j��	"�
��f���hf�3��[�S�qzu��� T}���9lG���{/��l�;u2Ξ8�����>�Ϟ��y29{�~�s�˔��F��A*r���H1-�>����t���~.��m�A���4������3O������W~�Z��bgB�e���tŜ�ѹ����'�����_�g?�ߍ���8q�p��fιӧ(�`���7o܌�/֚݉Įvc���4�A���mJ}/���#�����Ǉ��T�:q0�:g���#g�ر�O��>����W�Q� >fں �����ܮ7
�e������ȋL��˰9BB��wX4o�ce�^��C� ��o�'���9f''72�n�i�z�_��̮4-�i��Hx��	D�f<�G;
�����i٢�tʟ�a��{E;���g���N<����ȓ�[�.�`� @ɯ��.����]�������{��q��0ڻ�y���=R�|2(�-���
����F0!ϊ}U�k	��v��J3�f�J�_'n�D:啈�Ϊ�[�ҖQ6P�Wcya>�+|Eʫ�is�ؤ�D��[��n��-�e��͵d���������_����?���G�cz>>����'?�x������~"~���B<�ģ�@�T��3y9���2Z镳t����	�n�Oz�Oj6�eʂF1�f��7��14�cc�0�fXU�Y-�������(�8P�}c�9�ў�C�����l,���`�7�;����h�bv��Rg�`�C�m�Zo��*��ӘB|��q���8z�`<�/�>�V2Ø)� ܟ��O�/������;���κt�W�#�J/�m��:��<W#��a<���/�c���9V~����]�9��x�	���z@�Һ��!-r��jtٿ���y�>'X�ֶ3O[@545&�$$�h
R���t��^C@�@�^���
���{�e	���d��{e�4
(��7������~FӶ+���GQ��W刚ID�i���?=3����/��A��)j�ɣM'Ci*T�rq���R�@d��bv%3����^���q�.�cc��Dɫ��v�U{Z� :����qj���C^M3�#-;\��ʰ������ѯ˹�rbd�#�y�J ;u�X|��4��z3� ���2�r4�NG�ln[iLݢ�тa�W5�_ZJ)[�o�(LO�v6��_Br����0��'�e��Ȝ���7�$R����3�<z.���G��P�wr����$fm��)�[�je�*e�@̾Ͳ����8��M����O��}�b�ā8y�$Z��1؏q�{vO��cmA>0�Z�}(�JD]�}%J:�/�'U�&I��ɼ��(��o��\�^�D�ޓ�?h�����pŗ�?̻�üHI��ޡn�#n����"]�a�����w�A�j���
u�yk��|}�i����>6�#�ˋ`B��i�x�~���t�}�{m��ᩀX�ڪ�̾��#8��2���2��zmc��b�;��M��ѳ٦�@O�B�G�_K#&Gb�L�8��íA�$�^�z%�Т�"��hn C�*Wu��	P�{����1Ϲ%�K����T��!���&�wV����ť\GRf�Q0hk&"}	��e����E�_��H�d��RZ�T�l�Z�)8��k���(���hR&H���J�p���q�����4�VT^�7�r%�SM����k��2�n�5N�  ��0*�`Y`U��~�{�YE��ڮZ$�]�0 y��!\�(:S��=��H��Y>�N�l7���,[��]�=[���8�P0t���Q� �a4${�)ڴ!b�[k �i��RC5���HPc��m���v��D��<f�;������^�y���)�C�Z�|5�Ji[����ﻤK1�)_��@�]�}bh.�I�rH��l���`ߊAMۭvԢ�ǞM7�1�]�܊�u����hn/Ecs!�V����Cݭ<��g��=�����O��X��޵����hm=�j ��|�kn-E�xj\��wm�8f��y��ͭ��Y���Bv��Xc3�k[�ϭ5��i7����F�{.m
X�ր+x��6V����� ����9��̙�O��G��7���g�#��d��/%�d*�=XiN�s▀�;�;-�4�qCXI$�o�i�P�w$�L��gڞ��N	�36DV%/̲�FZ0�fZ���h"������}_�� U�����Rq���h'�G��y�> ���bG"��C༇-��5�.�������B���5����E����A�Ppz��:��A}!�l��P3� +D���WzA\I��������P����[o]�4J;<0(��:\��ʲhGS]�hE?��#�����l��,%��n\+"�)^�1=�eQ�d�!Ҙ�
{��4��	y�'�C���R�Ud���z�wi�Qt���o�؂IS�u5��[C��#ه�k/���t4�^ν�������=�9o�@o��D�R�p�߷G�1O�<�����k��ǻ��H����j����x�P3�L��#���cC����x��p9?5Os�̉�x����F�==Pv��{m1������t�<�u�}��Fw�/���%'T*H@޳	u�љ�A\��U�ET{�!�+;Vo�ǺH�:�B�i�K�l��̏�d��> �����l�6 �	���V�Qe�Ϋ|�X$8�w�kPh)u{�h�� y );�����.}��"z �UM#��~�p�D�@�<{�x�?�h޿u�N,.�,�с��(��à���w�7/���W ����|�_�#yHf��N`��}����P���1==�L|�����kf�ϝ�w�����G�Xj&9�L��,��(t�J��i<^������C9$w��X^^!�v���đC���f��+_�r\�r��WjF����n�cѾg$�պ������O������s����Sgu3����nފ�^y#Z�ud � ����ж
���,��K꠽Ӵ�\F����'�^W�s�@WJ�@���k2K�����y�<Zo��h�i
�Q46��ؾ��@�pb^? �o�����@o폱�Lv@���7Ԉ�>Lݾ�x��x<u�T<v�h<��x��3y������gO�S��������O��?�l<���x���������}������=�x<�����������г���~����>����a^��������<>�?zh?m�����,���'�ʚ��s��)����&��ǏF�ɭS���x���"Yӝ���!:�r���6��n��s0S�:�ڑ��t  �͈PH �Wk>JG^;�T� ��mF�Gu>g�Jp�ڄӈ�4a����v`j+��B����``��[�aG'yܰ$������0Ł'L)��O��щq��Z����7ަ.��d\��N:�W���^�C��ݎ���3O=��C�cee-�#��jȸ����3���br�~7���h�+ڈ�ǔ�wǁ��q�ıx���q�|�ps3�1����� @G�������t=��U��EZۆ��pF�p)��c߁�x��'���# �F,�/�N	L� ���A�m	��ƥ�=�v���`'#��\��L���uT�7��)�^W4���\��~<��:q���t�<�_�{'SJ�lG����(C���X��_�t��g_������:c?�=�H2�'>�|2���٣�����L|�#���^x`8O�����GN�'=�O���'�������GN��C�qx�h=�q�p�7�q$Np�}���\�F����P���6x>0���Ʃ�vG�F�P ._��4����v 'O!ج�g���O |���0gЦF�Qv�p�i���( 188�)���������k�z�lˏ� 8ϡ0=ו7����40_�6^��#Ů�̕��G4�]���.������:�<���,i��Ug����wQ�t����d'�#"�+K�0�YYu4��V���v0on9:��������J��E��H_UݎY�ng��0?�g����@�A�W��x�U��lhb��TǍ��2Z֩�`�G-���a����h�h.�5�F�"��\�QW0ʢ���Y��-�����8M���_�[��斖brv���9���'��7���}�:�,띔Z�J� a1�$D	0grz$]颌d��7�f�g֩Ǫ/�A?j����y��Շxu���muG���}��$0�m���~��4�ch���>���?�{���?��/�'?�>��O|�����g�;����O�?>����F����񑏿g2F����h�u4j
3����?����iB�jw}�U3���57�i>;�;V`�UH��Q��c'���V,���V4|�Fp�"�"5�}�C1>:M�~!�;�FX�ў��:ꦀ�	��>Gj��� �9O,͌�
��aH�P4%�I���qVvzI����y��$��
kn�C��P� �|���HGIs������l��s�7��Hr���O�6isߣ)�����`��8����q��C	,�>%����39�3�1<�� s��{3����17?�y�7�&��##��d��։������j�L�ު�@j�H�L�@�j>s��jl��jA)k!51�R�����&��r�Z\�q+V�����fll�4{�|8;Őz�ܔ���|1�6�)�1H�tՒ@�nnn!��{�08<�f�ZmJ'Ub]z�* ��svz��<�=��/J-}�9/�D��v<Ւϒ��w<�r���z�&� ��[���?��t���czR�;�QkX>4��QX�䉃�7��ϡa.���,��dj�}��������B;Թ70�?j����~ڪan�b~���D����>ۍ�X��h�"̍�~46jñ�;Ľ �xt7'��X�?�\�O 4���}Q#L�����sop��8�CS����Qw��^��G��B��Ԧ���F��!��zu���cxh8G���.�%�LQ�D��x�Wa����~��b\�=�}"����ia�\Kc@f��=��Vv9���SM1��0P,��Z�y��Z#G8z�dP)��j��(��Tr���:8K�r'���<4���"CZ�j����ߌ���x���b��.��X-���s�&ǹ����XV��k���ߎ�7�r���2�7=�����|PovSm�y�ES��A�ܺq'nܸ�C���_���_�x'޽~'�4e`f;y�N�9�a�:�rU%4�Y�?'�#���;W��-����b��-�����7�:f���
6�JjUܭ���	MP��v�jE�K���Qw����\x���W���Kq���h �+�]�� �E*� Ί�I�KU�M�yhx�
۾�8�0	�0jH�J�� �]�4Uݻ��|��$�%�|�sc�i''^��=h�|B/��
	HJ@�Kr����?����g��������[_����V\���__��S�qg~#.^�������z\�j�;7��ǻ3mxi>����x��l�y�NܜY�3�x��$agcri3�Pׯ^�7&Wbfn+._��˷g��\;�ޙ��W�cv�7�o�{;�ïw����;7�򭹘Y؊����[�cn���\�?;7��ηc�?!t�^�SE�@�Po5�^�>u2=u(�J?�#*��;�	%�eJ+3��)� �;����[wA����o�_����Ve�ٻ�H��\	����m�U��-��Mת��$Q�%v�mdG%���X1j��q��R-?I2j����33�|�:Ahx��1"��[e��m �;F��-�k�=�����dn�;��2;7w�މ��j|��ħ>���}���/}=.�v)��¼' �Y�F2�j��}�Aln���ja3Μ<��9��X��|��K��|'��:?�󿐚�����ͷ/Ǖ+7�xH��9�5;�M|]y�&�=[N��H���c��SO<�]{2f�緿�ML�I��OŇ^�p�n.�/�|!n\�S�s1�Q���u�䥾�|A��jԗ#=�q��ɧ��c���ݶ��7�]�!�Χ>����'>EZ��o�ko]�)̍���v���P�N0��l�<VmX��|���&P��~i��� g�kK��{~�����ݸ�~C�p�C�}��K@�%BŇF7hb.]���/}*������@��ֆ�/�q-~돾�߼S ��cM��M�	p�b�?�L��t.L������9�1jW+U��7���+h7r�F?Z�p}8���s�"ql��c�1�&좣r.@��2�0w��d�W��><?�i��>G��k���������-�eja[hJ]~��I�C�W?�D��g��������`J~V)�h"�6��q9=b��WVSٹt�n\�>E�iX�v��zD��'�  ���L�n�bo6�d�lV�q�L?�S���*(��(�K��p;���xK�Co����y�u��j���U��k�G��h��}#��ӏ�؂�^�vi=�tq��%L��XY^���ƻ�^%L+W����׫�>7���-A�PW%���D���^Լ���vs9�����K/��n�BR ff�������71g��]��F#p,�쩕Qn7󱎜n�J�^l�qm3��D7?�� ���hn0ᕫ��@8���VƳU�)�j�!�܋$�9Q	�d`�1������]��ܾq��aҹo���\��@���f�m�M�-���͘����`�˻���/w\�y����|�\z4�}�^01	GfZJ���*���	��m;��v��C񼷆��ę����r��� ���/��f|��D�G�<����4��V���p������E{YX]���fp�E�g��-���R;� �e� ��N��*��
�y��-cg�=��B3^�4_�LA��#�q�veݑ��3���]_��s��ĳO����4��x���u��nf�J�� �G]�!�Y?g�����ΌtS��A���i×Jue�)��K�8��8���Q0�uٓM2@nHCR�V�ij	��)u �_x�=�;�σ󪣴��<��S��A�aﵣ��sX�5y�
e���bLN�<a�1y�FLa|�k���7����	�L���*�:�G|��X.L��pR9�v{5�]���q);W�wծ3CW����q��71s�S�MP�'��A�ͨ�̂�R�Q�-�;5G�ch�?ryiP�SSwx�7�24،�qᵸ��+q�껱�^��~�s�Q@��s��Y��s�.J�a�;jt����~�]���A�=4�`Ϸ����o�+/� ��*��Jr����2��ci��ޕ+mW��'��"��MW Q���9
^�J��*Wy�s,?�9g֢�;W�A{�{d�n�{%��%���EV������1����v2\7��f��}h�_:u��g��vh����^u��(Ĵ]�a̐Qlܡޭ�ٌ�{�����T�m.E}�fs5��mt�#n���u��
~�hcA22<�Ν�>]dE��H��Y;º�Z脓v�W�v�!�S�FƟC�:�kY�8�����@�4R5�=3Hbz�%c&.m�E1		 q��z��o���@�	�4Mȴ��
/�yz�U�Za0�6�[���e��H�����ۨ�10�G����c?`�|�t�s�~!���YnM �8��LаS)M(]����@�H��s�VJ�����ȇ_�l�ϝ��Ǐ��Chw�1�wģ^Ǥ � ��<���bm&��1��fÎO$��<���e�8766Ǐ�zcyq����Z�}5.����DF���ƚ��J?��j;y������:y�Pn�ș�U@���sm\g3=y;�9�a��7���V�������8�q�Y�����lW~��Q2�I��'Iz���r�e�D`D-����lU����m�i�NGn� �3}��J 3
]�I P�}q�׉��X�h@O~k��V��t�j�F��	A���5�4�og��c466�˕��^���ŻK��;�>3�8:���4�������U�D��l��D�Z�b����hn4dݕ�vyߑֆ�N}W�Щ���+W8_��eD>�;��]!B;Z�p�A��0N�J�/��w��JN$0^>��S�i(M���L�+	�u���3GnL��$�z�49�_�W=���d�:6��۷c��ȱ#�8���q���8u���m98���LN�r�Z�iVXf�8� pn�����HP�܎:�9s:N�8��1�yJ�}�U㩥��^�NCB�and� N4g^{�jͲ8$���!x��P-1Ф�0����Pj��_'^���5/Էd_Z^�z�y �H�
�Y ���� �Q���$�i>|�u6Μ:-���U@b�72#hR]��6�rS���$�f���wu�G�١�ԬqPl�RQ/�[���t�刢�>�&��_2>e�ׂ�ixO�ִ���'�#O4��ߌ�`����8�sӱ27����9�[��uG[I�B���5)�=�Z .�Xo�bia1;����ς H�9Xn�д,N�\'�X:�-�ea);�ڑR��[��k�,iV�Q �"�ﲑ�5:A�2��{!����#r_Cg�X"�u &d8��u��x+��Ɉûep�5�TF��NTAġ]��������"@�T�ǲH@!11��}�ǎGM�����3��a��_������'���;ws$d`�&*��0Z�����=�}S����&[ݘ�h ���G6�,&�;��:p����W򏏏�8]h4����1::��������Rܾu#G_��?ʔc�ԓd+�7U3�C	��.�j>{�T:x ߕ΍��矉�{&5yh3(i�F�P�������+U{��A��<|�(&�@�I?Ǔ�ǓO>��3������TKB���a�٩�L*��U�t?]�y�B��$�Z��B�H�'�P_��'������<�o���c�M��}�u�>h��1�ɩ.�tA�u3�K[�n�5[���ѽَm��:�^oA��(���ZA�5�EP�9
����0�}ϝꫯ�mAw��=5[�@m��n�떔+ГFHj�_��E�@����&�������� .AF�ŵf
E��ԫ�����l�6�Ív��}L\�RKЋ�Ο�l#�?$p+Q��r��$&U�B��}	���5���HK��d�~T�p���C�yE��},MTA��#�)G�]��J;{uU���3q���hw�¬ ���.�;v�x<��#I<�1�I<Jm�ى���4n`��NCכw�ؤ��2h�>u*g��<y"���|���N�S�Yo����+({,svT+K��e�Q�G�Ch;��������iv8BV��UI�ږ̕�Ľ��kXT�b���\[���o����(O�v{)&���o}56�X�Z:����{f�G8鯢����po;���_�wy�4XF#�o��j{��n"�Y�Yb��BH��
�: �\�^��W�5�V[��nʜ��@�)H!�:��~6�sQߦ����ke*&�1���]+��\�8���碹���2����Y��A��� ���wc���=��<���� ���N1�o)��E_���80��m���\�,�QL�SyX�6��5*�c�54����t[�Р��$v�U*Le"�G:#ыs�|.���@�4�ԣ���k` Ɓ�]��I�tW�T%	[�������a5ێ�E4	G�(V���spz
��^��s�!1�Z@`iR�u�ao������+��	�����À�A����R
�KKK!����ڑkHl�<���Ea)W,/-Ü������M��Gϧ?�t�;d��F�е��a=��l�QpG����^�������(��/�)��8�1�FD�� �]��GUP���^�CQ}^k����$MGM$UZ��90C���g�ĳ��!���h����6m��hB����u~��8���n*��p�
Q��s�'O�Ȕrר�+iri�6)�3�Q"R8i2��L����F(�6����0
CN�+�@-B��k3F���z�ꋃ���Gㅧ�cc�g{&j D����n&���ǎ�O��D|����O}�����=����/~�������0@�9��٘h��h��|��`�c'&��Ϝ��?q&�i�E4�e�T��[��m��m=�Yt	Z*�+	v�ɶ#<h���{�d�3�<��+ �;������\�I`֔�Jo�رj����z�P%֒!}^TB�y�zZ�y��Ҽ�bj4`/��v��^�U��B;��x7a�M�~�P�m:�<�ރ�Q=���n~�-�M�NMƝ�wr�ՉrKKؕ�p/� �CϪ����B����PR�,�LT�B%j�PY��>(�`�GtE��(�	����E@�E\�%�ZϦ�sxnMZ_Mg�ZG�I}9����T�搡ZG5C�g�=������z%.�eQ��>%� ��3^?Ҝ�E?�>;����,@� �`?���s4�l/s�gA���kr�%,U4!���V
	�'�:)u���cz���貃4��FHոֻ@@/�X������ �[��	��z���!��}�B�*&	4���x������g�~��O�?��_������������؈��������<��_����~�3�����?����?�����  ��K�|6~���#4�P�Jhř����������Ŀ��_��G��.�j�~L�!j��5h�ү��B ����W������3�wx�Z�iiRL:��=�:m,}ut����<������L���"@ձTE.���|΅G'��3=���
��U�\�����0�@t�,�+�	n�\#�:��Ƀ�CB��˱H��{�G?��M��$Z]F;�a`����~��f���ɻȓ�i�mW����無���/+�[�,�� .VZG�smP&t���4�/ĭ[����/�o�W�]/�Ax�%�Wъ�vN�*�$ ��i�9��sM	������m	�!�w�^�WH��][߈�wn'8��~<)W�D<�g�v+�x�=AC�5ɜ��ƅq�ƍ�|�r\����^Ko��p0�5L�$H�3i���D>%�P�@~"�dR�ŷG�|��wCA��Ͻ xMs]�MWM����m�)���>9g��	^F#��N�+�$NQ���8vp_|����ܙ�qp�H�7cd���l|�g>��韎G{,�?�D����L|ⓟ��ёXD(�h�6q��6��6u��ss�S��t<���8x�@<��9��X|�/�M�����C�7G��Kv��&��!�
��C����Hm���
o+¸�ԩ�i�����OяrU.A$���e$;Y8W��	.~�!����J��p��a�K� ���n�=�ʫ��{�3��
�;�쨃#mT�̎��}JQ^S�F�Ӑ�C!��9��V��-� %
;WcC��X��~�"����L�˯�/�����אĘM�k^�ȓ�Z�R��Nw֪���N~��v,���[���� ��$��j|��ߎ�ɢ�|�J�����*��Z� .hw�_4:>ãc��/h2qO q����|��K_�J���W�z��y7��|�A�m��%�#��S/jV�0��S��7���Ks2��㺐� ʅ7�H@\�բ�p���i	$
�'i��/}�<�I9�JMW��^M��Я-��pVl�[��6�߄�68���bE`�{�Hg�KCηМ�+���8J�Ny�,��4c��P��.�9�����9����g���W�����K�C���|l�֣�/a�,��f�%hm��h=�̳���L�¯�e���x�C��������;<<BE(4�}�z�b���W�{�ptr��^����K ��~~ҹ��h��Q0*�P�v@D�/�Ŝ$qS+�!�ʆDEIB$�bd�����D�>��@bo�{L���~��z��!1Aq������L~�d�ǐ=��;G��9�|9�ޣ��Jae����[k��7�ߊi��49=���������H$BM�7ގ��R�s�2LY��}f\�j���f,;�ƹ{k޽;��%{]�58oܺo��6Z���P�P��~�x��+��8;R-"	�c�F�y�Cy�D�ޝ;wcjz&5�F����s��4��`5ߟ����V�og�C�����%��\)�R���g���v����9�"�(��y�djf�z�ŗ}RK�Gv���?	g�R�����,�]�}ܩ���P)x�$��5���~���G�B�u�)�f����&(H�{�Ȩ��9��*��3;l�wJ͝�?5
w���g���������_m�[���ٻ��ca�Nܽy%�n_C^�:�74g�֚#�?4�C=i�Jҷ󅜅l���F��Y��Y~e�2�#����Y��Yg�o�X芹?shp0�����
@��70���q��$��bז���3���/��<���tJͅ��HFP��9�e?��99���06ہJ�z��ș���$,'��{/����Z�A���v���Qَɩ���-+�7�'!���	HW��g`�M6{�y����h-jS�d�5�+���bzf*�`xO�N��RSQ3�ռ2�����iɴ���j�֟^�EuW�]�w�\�4UV7�Z��&��Ὃ�\�k7��̌�$瑬:5�����mmq����{�Vܹu3g����PC�֎P,�����Q��ԻC�ꑲ��A�ie�
H:׻~��mx��]o�>�~z$��K_.��|�Q���E]נ�>��[��ݦ��S�I/RGj��Ѻ�<?�E��E;�����i8\��k� 359I{��)x��U�C�ѳٙI���6��.�;y�:���+ηA�f�s(��øK��4��jk�v[�\��۷'s}�;�ۯa>Ϳ�/�U��
���B�<�ޮ8���Ǐg��������$�֥N^�0�[;�}�rrZ��Pp�꽽�˘w@�\��]�!P�Ml�kT��i�8?�*?�L�F�	�v��B�=h@�[��}<��Q�0f���p���еf�_�*�
�*�f��F�"	eV]*�+�� �ȋ`��.!C�ۈ%wu~d"j�b�������<��f\�r!�foCh4�7���L���m�$�����2*xK�㚛�XZD+�p-L7R������x��+���Wbj�&ug��z�Ï�$�x�ݘ���S�
���~K�����ڻ��׳�B�p~K`�w�\�;H�y��a�����{m5vf~1~���
&J���k��g�1�b~�.�# J�����(��7�`��O��ۤs�\���G�ȑ}166��r�}�6<q")�V���Q�Z	�uq�u%@��'A�R	X��V��w�%Λ�� n�c~h�ǚG�GF�8y�y�z��uѢ}m�Gڟ�ȶ_DS�f��7@��8v����>Ll;����� �]�0mgs��� �
.#V�bM`�9��MrM�<�[�ڞ��_���F�)D�k ���3���ȵ4K��?0F�8��F�P�x�;��Q곟2���na^�I `~�}e�	g�ɦk]�2�i/��Vo���b�Y�/��r��-��P��S��u�i�z%hv!��s��-��S�Ms�dR�ϣ����!9���@sD�u�97��2�as�
��~'!�#*�c&�;=� 4�*_��C�.���_��x��Ƀ�n_�r���3�ȑB��d�i<GZ����x�����X����4��p�C}���G�Ʊ�Gblx�"t�-��0m��h�3��9�gz�<� Z�����As#�����h\#�1��!ږ��b;��<$(���䄣��r�jH���ȟsN�9�����q�Ё�@�;01gO���gO���9��[�$M�͎SG����)]Qk-��R�9ǎ���>b���������Qѩ�s~vTS7�ԭ��՞V�������PW�N���|ʛ����9������j��~��s����>�SS��j�z�i�y��q�Y	�i��%�A#�����B_B+��a��r"��+tّ�o��˱AzCC1N[fg	��l�Is0���L���_$��]��?|�嘚��0��zr�m�΅�}h��E=գY�`OW-�Gƣ�Ց�����c'�A��sU�#bv
��pm��#�mS�h�Y��yq
�_sP�U��w
�ȫ{�H⓳�zpʂ���,��u� @���DOfF��"�h��}#�km�<f����N~��a��a���Px_�v!T5�d����=����a��)�e��5�U��	�������\ܺy�
�GE��۽q∌�H�;}.�|��x�g��'��g�|f<~]?�� ϭ5�d��_J��.�m2ڪbl�B��Sg�� #����q���d�SǏDS�ZYH;�al����C]����#�:kU���o��|���8z�h�O���8�"�nc�����hQyt_�-4�M���qi܍E� T���혛��_����8}�X>�/��C ʑ��  ��
����mƝw�ʥ�ܫSp�v�/���<h#�# 
���i�@�>.�d.�gWj�EXU=����u>�~�+GG��Hm9w�Yʚv��bY/�e���p��[��fA���70�nN�����I/UD�n���9L���L�j6f�!駙�O@`/^��#_��|b�3�GGcx��F�:�Ғ���>��bߡ;�ױj �u#�����12:F\h����f�Z@`N�N;��Dv��YMVT��.��A����b���X�=V���T#>�x�6��y�����Ϫ��P�xrؗ�� 	<�(xߌ@;@�	��|��f�$l!�|��S{8����t2y��dH��p<��4`���tf#'�5�!ܾ};G���F\$���O>\���Ȑ��@�E�4�y�v���� ���^�v�^�C��}%쒓�c���m��,��� ���"��a�	�f���Q	�4L�͘Q������Ӡ]���	�;V�D��r�UT���%,{��}H&7YvN�r���Wݮ� �6��[�46�~���|;�I����Nn����q$���C�z���A@�$����X]����iʡ�S���_Ǭ"�!�m(z�OxtujUSS�Z��j�Z��4��Б}.V�z���0�õu�����l���6����g~M�n��^86�aڨլG�w���u�Ⱥ�f�f�EJh� ��oO���e�ց�м}Z�N��e��Ѳ�?�\5;Hzu����Q^�E���b���I��Z�dܸu5.�{1nq\\���|^F�9T��y��a����o��*S��Y��%��\���o��|!�)�+��ɯ����]��r>���)��+q$�՝ޓG9$�Si� >���
͝*l޺�D��{��t�u>+>��S�u|R�Geғ�r��麖����f�`ʭ,��ޔ��	�:�=
���~�wh�n8{ߗ��˨�����Ht�O�������l�����Dr=j�4�b�����=�v|mcl�9D#�F��w�P�RD�"�����nT/�܇og�%��9$��64؇�K<���L4��U�I)J~k�   �"�߿8�� 0�y֏w1�P�#��z0�I4W��7�yg;���A2��}`2.#��~i>��y�=�������3���p[s�W��~�lua!V8�8��Q��ZX��{�K���\��i/��i|܃;����y
+�Ά�H]�n_���W9W�tg�l����9P!�pR��uR�h�׎v���-?����Eރz`^��Z�a4౱C�eo\�>?|����_�7.����q)�����W����o}9���?�����y�f��x��q�H�~lb<��&�N�!������= t����}j8Ո�>'κ'��N���x��sM:Z Ƒ��,��V����0��T�s������쉋����	��v��eA���H��{�d�vƜ�Qe!p�Ȁ��N>�<3��	��l�df9�2g,.�_�����k�>�ˡ�+p,�5��������c�<q��F%E��˚�!������pܸ}3��͜�N��:�1?AA��pBRn�Hi%?1���MfL��q+I%�А�1�H/��o@�c��� ���E�����R�H-ȅv�<r&�{晜(��ulpgMڟ���q	�k����K�&�T��Q3��]���ǎ��C~.�������c�ũ�p��~���# ���H��O�>�L�#�N�� juL��Α!�& l�짠�74��P�͖��5z����PWՌd�k�V��9G) p߷?ǎN��~��g�w�� �.�C�֑Z��� ���L�$�j)H8�����f�Z��w�M�y��@���	���7߉�^���+��0�uL���=���Оn12:��3 ���ګ���cG
�q�W5�%H��{�� ��6d�0�#������ѱA���"�.��N\�O���1��=h(A����g�y,N ,��� �����Ӌ�����R�6���b0A����;O�ۏ`����uP7��)SA4f�#$(\�~d������{��a|�ۯ��o�2#�H �ǆwBO�q�T�i� ��#
=���T���nC���m��#ak4���;H_*T !Dv�r�*�}#��(����L�ʍw�i�I<z�t���5Q��ۭ8r�;{&	n��1~W�
H����(��/���A�!R�_���#��;�\��6 �C��;����)OS�k�����{�R�fs8�\����_��1)  7j����;m���A1�G����G������' 6�w���|��� �����br�nLa�/���~N�3��C��P�&���_���0���I�扒������Lhn������җ���_)�_���>��r7�.4%��$m'��)w�~�-�Pu��<%�X�Y��Y�ַN�����fwT��֑�4�D���;C�>�m���3n�e��m�}��Ҥ#n�i���m�w�;9y3������������Ň?�8�h3��_��ߏ��ǿ�}��ԛq-�km1��_��8q�`(�0���J|�+_��h#�Y�e?M�<��Cڱ��o;k��{wr:._�05?��O!�Q�
B��܊���g�?~5V6Fc�E�iw�!;�'�����+�?u�ϑቸ5�������f���)��hJ~r���& ��??���a��� ����e�D+�F�(�ɸ}�� Ʒ{���;q	��ME��%jS8�{�@n�u/G�*XoC�P�0����6�������)���{W��`��h^@jEw�0O�= R\�r����j��{����_�K�瞎s���r7"Vլכi�P�eX�=��I�o^|'�;������TG�$vhML�C��ºC�9v�x��;��D��s���Nw�(�C12��s<.�y1&�f���؉��?̳�8tԴ�̃H���c?�ú�\�A�<�3��$��9�I���eh��=7������y����L�a�49�?ss���f�>����ܱ� qN� ̷��A�B�[����!�X�[���_�~�f�ɱ]�ɥa�O��f���Җ��R���y�#�Z���Kx��	T@�҂�O3�Q7 �;�e�s�M�'�MGޠ�\O�;�Ve�-�k](ҫ�%��N��?�4�<y�>��ŋ�<~=�V0ss#"���Y[�O}�q�v<��a�}�����=$=�&�c���	Znq�:M�@���0���ô�a�i�:�oƛo_�-�� ��{�(������� �.�v��?����ߚ&̓O���g��������V|��1@��j�9���:��6Ts���'≳r4�2�"���S�_'�R�yJ�z%�m�Q4����
kW��s�%C ��C\2���mU&��R�N?�_H@�Q�����4;7���z�KB}�\��m����Ki���$~̀�&�6x������Ɣh#�t#	bfn)�ܙ�;w�cva)�����܉+7nŭ�阞_����q��d\B�x���<���71��@ awiw_?Z�D̠|�/ū� �.�z������F��3N?;;S�h�[7o��K�`;���9xGo�ޝ6�0������|7�菾�����ޟ��[���&[���]}��Mǻ�^��|���߈�r!.]��3���P�UM��H�;�`���,Bc�o�Q4�L�@qs����R(6����ٔN����dx�֠�]��Ҿ�m
ۘ��k�^{�0�By�sCl���q,��DKsHf�_������Q�'����bOgKCkjhn砹���.�P깬��jvHf��Z֑8��W��g��м�_�f��/�7�������@��Gh��F5L�5��K�\�����}p��5p5�o��O=�d��|�p/��h��	Y謁6��3j����:$?��u�9�Q��˓�c�I^K��;���й�}e՚-�����h"6�3&s�)�H���)�OB<���S�lDN�~�?��"��
�A���D� �H�k9rR��e�s�)�6xJ%�H�%�!�8	�8
��ix�)!�$$A!�(jD��6��v��e�N;3��a%�-key@i UU�ݪ  �y#����_��/�x���Ugl
"�q{�ݫ7`����vf�r�F���ո	�\\���2��:8<� ��*t�nhd4U�/|�w������T\�F׮�5��7o��wP�'s6�]�M�p��}�H�{�8m���jTN{�җ�_��W�u~��s��u���t9�%�+W��/�Ocjݾu3�^}7纸����Z��>��[m[��t6���;�/�忉o\�>���:u����/�a����>6�9/�A�wnˡp��k�3;�l#�W�x4_�$���v�_h�y������~��ϲCt�y�y�ם04m�@�S4�Z?�4Ҵ��0����U` փp�<���5gNKO��I_�+�8����s��&b�+����~�t�ȳx���g;>��&b��~���Ko���P�?�?�@���s���)��2����T�\˵�H�5�e)�|�K7��FCт���^'?��[�$۩I�JjQ�zw<���q���jj�
�/���'��m��òh�%��Ǐ��g�`���\K�C;zv;V�X��~��[�O!m���ѕ�Lx��$�d1`�,R�olq�Y�/��E4<`��`�ش���
aI�We%�7�[E���?���{B�(<
�hH^�|�9Y*��nԢ*��[oī?|9.�~!�|��x���r/�>'�����əx뭷a�/�7��M��s����\2���7s�N5��!<��s�=����>���޽|�g�q���x�����0�k\�s��߇Y]q5o��$p��U2=;�Ms�u�]��b?A�
@��W_�o}�ۤu3���<�j^5)$z�i�������<O]�V����,`�N�ŷ.�@z��{#���o����/��R|��_�o�[q����g�2[��QO���d�\��i1�	�&?�¥�`�P�W���^�8�ao��o��Q�]�A��gR��X����?��:6җ�ݾ�oB�9Py7㆓�6��Z@��h	
Nێ��|�J��M_�p1�x�2����Z1� ��ħ>��\��w�/��%h�;&@;F��5��r,��@��ۡS( �9����&�L{�����_X����\i^�?~���?p���B���{h�����q��O�E�%��Xd~���қ���򾺺��ӄ%@P��i�Zҋ�=ii�AzՃ���̬��H�	$1 � �nt�m5��7�ߛ�����&S�_���孮*� g���6�cGĎ��^�sW�1��%�ڷ~d�[�,dv������*�	��;e����x5'��*9Q�C��"0$�r"�j�OH����]]R.!��Kjx�@JeI�P�$ `x����|-D��"��A}�^c�����(ueq(<��c++�0<-���(�ʐȡ�|�a��M[]^��{���b@���U�Y���7ߴw�}O=��v���� �`���w�+�7R�m�� "��y��������V����^Q/�r$D�^��BbAsca��lr�<��� �~R��� ������,�dI��
�հ��7�)�8D)6���\�khX��1 ��*SBd�*>軱��_�o�S�+��Zݶ��
��R_�=�©�T��JͅH5X��F�a�X�.z��UXNL�<��3w����:��~���4)�8�v�=9���1�*?R���g�Z���Q�	g:���.g�������F��U��P�2`��j��Ⱦ�g��j;�B����gM|�"ȼ�Y(6?=e�e����+�.W��NXU��1�kR�*�q$:�M��ȴ�����[�)/F"�]�����!���=	4(�}�����{�{E�ŷ���`
�9=����-��|�ѱo|�e	�z�_�pL �!�i՚��G����ٲMO�Y¬�Ea���E:��]���
���bR�3�y[�h"���ԔTGItң�0؊}Lc�Kp`,�SH0>R&A�A(1�� �s����9Fs|�ZKD/X�LY�� D$ő�W5�zp�wt�q�Ӥ��~r�Ky��o��}/�E��r}�I�,Ģ?=��L���	ËG$@�nd����)�bQ�XY���j��F�gL�r��}�.q���J�v�X���
�z!��v�� �|��p��@Pb|�Z�̛��P���YG2�2u5���s&"<�F�# Q���+���7{"\z��ȊM�$�0��L,���0��6(������F�U�9�s&���|P\>̎y1�^B ���ƅAa�'�=�G<��GB�FP���,��¢,L�8�JtG}�Hp*�3tݺvB]8J0B�Vc0���U�|��K/>#����Mig�D0�Y��5U]u6=��ް��86���w�kh�;凙�Y�����k�h��GD{�]m4$d���R�3�+��c�i���L�o�oI�ݐ&�%M�oΈ�Fb��~�A��%"E	��kv�?z��d��`�"D��K��}��=��Γ�
�!Z�#1c�Cw �X�Af`|0Baa��D0j'|½9�+�">�!�M@�k�xL����(_��y��`Ud$A��"7y��jy � ���m������#��_��x���q�Ԅ80����)�h�w���B%@�<�ՂUPO�Ks|?K����}9�p6��"2	�q�N�te&���-a{�0O�vq�O�滕3W6z1 � �$ឞ����A�XH]�đ��*{����ۙA=ɨ)'�0�ω((|F��+Ix�@������A�?ؓ@]U��:�@e�66log]QS�s���ʳ�Nv� ��랴�> &�.�s����� �s�g$NOi���/��Ge�����Ϩ����w���ӳ���ց����h�\��Q��*�M��X�>P<��\����l��ؘ����n��i����j+7���� ��A�&��=AH�y��&�Д��7�vw8}N�c����?�ᱫ�ϱa!��G��u��S��Xy͞3va���;L 0kt��5㳭|�5`����\7%1k���ኀe�"�E��x���<E���4�W~���%@PQ�B�p���%�`Ȟ�8�h�s�"h�m��h Q��~��z+d22�?3}��.yY5��H=��|��A�eZ�+�{L��zHzU�$8�1��Ą�%Y⽺*�Z��"flK"��`�TjD������^���ڕ:��م�TC��P��z�7���؀#9���ms���>��A�3��1!J��-��|��Qv�6�;�� ��I��e�����?PQo>6V��@4�o5�Tc��ܖ���+�L���[�ݰ݅c>�AOX(@�};��ےZ:߷���RU���Zy{^�M^�þ��ɞn������EuPo劊� >{*F����+Te�>�Q!D!�T�T�S����		Ssg�w�eVM�-���,������<CݨU��JG�� ���,���/��^�2`�hL�^���d�e�������юh5�;�̔�@t�k��"<
.���@m֓Y.�f;���&��fG�lG��u(=�QI�������3�!��y�Ke�oU�[
�usN���I�f��6w}�R��⻮��5	"i��=��MS+�x�ccy���g�=	yu~�~SxQ�������s�ތ��l�Z��Q�Y]��ėb�Q��g\��Y�8�BW�wSFi1��蚷*qt'�:4 fM�G�s|�Y�V"m���:��D����t��B�K
��vɗj�Qe��Xv��\x@/>:LMT	�yf
K�9�MߕI/(�9খ�Q�\ ���,����P�S(�WxI`�(�R�-!�Z���(%�e5(���s�7���"8�5ϿxF�(��1 l��lZ���"���R���UQ4:�$K�Y<ƕu|��Q���<���Z��3��f]Elx���@̹\�B@�蝈�,�j�����S��N}��('b*��T�/ƫ����a=� 1��IURZ�9``v����O[���N���vĽ4���b/>�>�h��W<﹔���=ǒ	L	V���L?h�)}�������>
_�!+��� �nӹ1�--�͒}	�}�Yi#����Z<7o޴�UΉa"Ae! �B�#�	T�$絠u��E�J`ϋ&��U���P���RǸp=�+�X;+`nf�gB�f��Ϝ:igO��S��6S�#f��Ƕ�Ԯ|�s��� ��z�m�X�'S�;{�&V�@|������R�W��O��#R^J�;�.D��!��'	�J��(�H� ��o� R��B��#�X�1 d�=��ȇ���� q��'�Oq}
Q�3���aP����,���Z15>6��F>N�ʛ社!TX�CX��,���aJ-�<�J�����'-��A�0�O� Kx�DX�'��t�?�1m�`���,]�GٮI�|�&V������t8�a���t�W�V$��D�hL%	𢈸(S�7�!Х�I�
W��{�O�㜎���/��Oj�L�[3g��z���2]��-��]U@�MG�w
�I��4��%��S�P��%��#�m�=�Yֵ���rv��.v%���te�&���;Rz�b���«����;w�]�x�?c��#��#?�+9w�=p挝=��Kz��]�p�Ο�`�Ξ� Y�]�v�ge&'d������}�3íi#t�X	h�ca����3k���b��p�x�W%�0��]&� "��y�.ₛ��@���E2�C8��ѱ��o���]!Xe@�8�$�{*�G/��� %���ۺox�s	�3� IW=�08�L���������%s!��^�]X&&�v)��u�7��Ȁ���^F*+=����ϼ����7�=*$����	y-yy݄S�C����[���p$F.�B�䜙8�T$�HE�K�ׅ����*�f2ر�?�H�"���}���0:LA0���$x�������d��ޞ�ՀQ1YNT�I��g5&�M�_[�P��6فXDL�f��HJ�g4��~B�������Xw#�s����q��y������X����1X'�VM��r[a��X\&X���$։,.���g�ʬ�M`ڠ	9wO���L�J����r�8��8��a���@�%���N�B8��'�c���!�"��X�a��o� J���A����p����P0��p�]I�Bķʂ�U��@�A�<�����[����c�(4� ���wq�Ɗ���@�ċ<��@B����<.�g�9d|�(7���;�Gx�pÆ�'	�xi�,_ǁq���'8�nr�{8�`���9�˔2�L��&�����ց�ML��E���R��eJu�e2�գ��u_W�S�y�|�DO��s��@�E���C�h&e�����8C)iH��RAFd���@�T�f��݁���#��	D���|��q�(�%�XS=9/���[u@}�\�T:L,�Ue�
GE0+F�(㡋��+�:�)��l� ����z]�3+#�c����Z�ݖF!���
f���%�XO~|��]H�fG+�XQ�7�@�X��
�ra��\#D$|�����9�H��L���rN]N�AKq�]��G�+!�@��kD�7s�(i�8 s��^ �N;qt����O3��⡲����d�I�'�qxЪ����ơ�����n0��I���3,���y�4��#]\ӳ_�����;|�����\`��#e���P��G��!lb�+z|�?�	������p�[�Fp-W�_qJ"Ȓ�����1�0&X�ԶeDxYq˼�Y��S&ͧ���ء�Ut%��{�wL5"ϼ�>'MiT��`�}^W`"NA��Իw���@Lʁ�9		�#�$��Y�ز&��,��D���ufM�u��t+aL�0a4p�i>Cz��9����ë8hjjƵ�C��2�Iw�q7y���3>U�3�VS\̛����f��Y"�V}+�p�H[���n2%-?&\��l@�P!�p�Бw����DX	�6q�w(D���|-��q��x�k=E&3�-�ŅE?��AD�	��1���{�;�������yj<Lq�;:ㅄd_��G0?�	�i� �I�I��DA8���ɐ�4��:��/1%�~�����8N�G]�+��������u��|/#K˻� b��x�}�f0a�ȟ�禸!4*0X��\�-���U>91�z�}����m�nmZ{}M~�;�����w�/3���Ʀ�76>�X�(�w��u����_��C�FZ�q��ֆ��Ζ��_J��Ukn�Yg{��=iNu�L��q� �p0g�#AP�����yP����k2��2�-���c����t<�ݬh��Knn��C���z�Ӭ/@�f�#,0�b3�.d��!܁���Mi9x\>��贋)t�6�G@n��2�zG���:�)���h���}�b��ɷ�^�����ΰZ��"�9�@$� 0�W٘<�ل��ɥ��	S��
J=Ô��0(�@S�d sA�^��  pHy>I�a��R�Y�|��4�A�#z#r����T&�A#����0Q��3�`��e��1��AC=������cp4�Qv��=y�<�'�7�MD�(�k��\!cD���k�o2m�I娐��E]#Oo����]����ڀ��ѶO�(g��\;<��bh���|��U��v���Wؠ]�5{ϴ��Jc
�u��&�b���	��zgM�'�Q߶�����]��e���ZL�gt��E����{rƔ?��-��*M�!�C{�lR?򕒍�sb�����D{��Ǿh�+sk����dr�󃎵�#�WdunC���Т�Ĝ���u+����D�zf�Z3��,��q��%@����ǧc�3K���e��f��}A<�w�i?��#�!:EՏ��k�[Z�7��ӳ���-��%�Ƴ���Lþ�&_ū��^���ǚv�C8��*�-�	 �j��C�Y\w �g�"O=�#o����Q�W�m��m_@Á�l�B�C�[�++\�g�;5�ٝLY)��~6�{�A���2=(\Vi�`����w\�A�����h�>�0G��������x���Y���K�F�q\=���S�I��a�p�҅�8Q�T7���"�h����S2\�wG�a��Ug榜z`�wA�c)���rF��2Ō #����<��� P�.S(�IZ�����p�������=��$d��:8��qּ�_?ו)Ut����N�	���جn��D?o5'f�Y^�@N����l�^T=���2f���K���k�ٕ�K����BD��W��ȍ�>|M�Q��,̻�4b-�"i"�6e/�Q�:	���Lt�)U��c�NMMJÙuM�B��1ɬS�8:�]�Z̚�B�~���������?���O�����'�I<U�% /9?�.����}���B���S'�3��%���^+�}�C�tB&%�3��FB�Z��b�m0f�8򀉒��� Yi�`*�B�č��	w�!Cz�6�1@p�m1����N����ic�d�C4�'��w��&4��\zNe�.4�^�y�B0L�QFԏ2�

y򜦘��H���r�L�2~D�!|�S��<��x����U���1v$M��J�������vŴ����#��U�AWz��#�gh�b�~)�}Z�S�7�0����'q�K���H�G�Gl�m�N[���mT=�4K�^��3��t�����]�|PO�ݐfqP�Aa��qk�~��yr�H�,@"i�u@c9��?�S���G�����nߓ��6g�aW��N�g�;���6�Vh��
��o�mC1����׽��k�pb?�3b�cn�m�r��_7%>�TLR`A@o�U�ˌZ��YS����M��c{��l}���#��4�:f�!��UP��>����\Pj� BBM�K��(h�1�qHdCG�{'��ݑ()o�0����
�"���3`��gS�g|�`ZII�GxQL��������G9�-K�<��T4�Gha�>՛�#&�¼/�]���{�"�)�8I��p1s�e���|����Gu�Akǻa��yP�
_.4h��z�����M���^�7Vo�jPd¨|^�,<�ϊpM>=��'f�n ��R��X�:PK�`�=%Y��{�x��s��'�l�y�.���¯��6^����S�S��%�C)ٸ��Jy\=|U��Đbi	�\��]�vӮ\�%	P��ڴ���U�'�Q7�v�ž�f�af� � ���h�iK��y�(�T�� ���@�C��4"������l�
ㄾ��|Zh�,�0��	o�RY&Uq��HF����Ĺ�>��|��p�u'
s��]��~��*��#�@h�0�.#ى�����!��3�\������n���_)��=���BAa�� 8|�%�� i%	��\����
�=�QT��/���B�E��{=ӃӨ4nZPH3�"T�W,�"�p��f��hJ�p8e|#�L�H��s8�)z|m@�Exj��k���:'w�������� �����-?��s�{���!��J�R��j��ҴTO�юʀ�j;[dב�j�| �` ma Ma_�=�w�V�������>{�{F�8y��nY�Ք�����Ā|��0����uO<�̍�ߒ�˴�a�`����_�K����o�1]�{T¤������6��Y�槽)��d�2y�����+� ���v���YA0L�ޞL%i��;�!�iC:"	@��g����-	,�p�~	74چ�Z6N���)k�BE�D���5� ��G�O^�����@gG��CZ
'��A�a*�\�DT'"�R���&ΜǑ睿�J|�!��]��Eb7�6��K������Z*RG~�#���-$"VRo��y������(,�s�� =DY�Y]��H��r�0��!= ���dFQ6.�Ap�@�q���!���>�w�!�G�T勉�(܅V�	�8�p w0A�J�g���|3��s��cWe���+�þ��%�繣4m��R9m��+������T���bB|�o�|�&���#��)��-a�����FV�5�\hY�ж�R�j՞MV�09b�5��JϦ�M�*4l�(����U6�<ض�`���]+�7�`���mbH��:}	7Υ�� ҲY/a�ɍ�[��F�=	0�łBߝ+�GH`�`. (�i�\���&Hݽw�n/��sq9^�7���,nݺ�ep$'�9��$ Y/�W3:�DۊVT�tl%\�bƢ�F��m�G�.�/W5�����L�1�![N�����Y�W?Z����+��ݱ��Լ�
ߗ�w fPA5Ie���W�)��w������A�.T|N����j���jٶ�W�K�N�"�P��Ίyٝ��#ֱ�EeI��vyU��#�ÊCI�n�8)�"�+��`�h�X��(0/���,0*��ǉ�!T\�H�(�'.u!8��B|�&� 
�CP@4�Ͻ7����{]y�s&,x�]l�Ј���+y�R�TǣW�t��Q�t�4�����D��%��"
�|l�%��gg��Z����G:��gz��*Th�pM��>ơ6T)��&���2�Ke%��e�Z��q�t����.�����4�*"�"���P�YH��1V�w愶���ږ]���{eJ�D̚҂|��q�U ��	ߣҗ�ز��]89oO=r�ʢ[�`���¢�qHt�h!�C��O�|�fc}C�k�9���A�kj����əE������}��ڲ֠(u���b()m�W&mU<"�Fx�լ��UONEC�a��Ĥڮ`��:8ś������C��?��]8=�z3��`�h����>�5|�����8P�s���k��������U[ٕ$�W�����b�UE(�9LaX�ŀ����+%kK��%i��ʒ�񝮌���n�"�7V�m��۩E1�χ�W�Ir�G��e�pʗTDT�%��%�lez'���֮KS�"��T�)���t�X��`�h@�	� 1K���T�Xa�hq��`:\���\08*%ZH�G�Ch(���#�3�~�ǹn�J� _��U�CA!��=�4�I���,�)?��)0�[E.�o��d@�,-b�&q ?�c�����E0�A'8Oyxi*���t� �7�V�R��?v���/�`ϝ�^����FS;��R�1oYs��acb�,��|�h���T'�2;����8�e[��l��_����������z��T�b�	�K��$ý�0t�6���=|zA���D��LPK>`��́:�Oo�� d��.��n�Kp)p��e��1A�;q�v���W�u�T�����E?��g����9��GFn�2��i	�3�����¬�����~�	{��x*ub�_��S�I8�+C�(|b��X�����bB�8�����`6$�SK�09�BN0��1�0��D��ќp@����K[�1)S�Ko��Y�,��ciM����� �!,��|�L%_�8d���Qfi��G�?1���
~O�x��I/�)��\qE�JH��J�x�q=,�È�{���1�p�XP����q���'啹#�Qߏ�	�ȏ97o(�[��f�}�Z�"�\H+�3�ȑ		`�^�sA9��!�-���@�9��J#PO���H�Kʰ,�Ƣ.QÁҌ�|ʏy<S�Ssv���6w츯b� ,�N�D�8gd|jފc�6>s�O������'l�آ͞8i�s�V�P���H�Ҳ&�l��i�����4�A��&̬�@uF[�J��
n�E��8�^QY��t��j�{6�_��Ѯ���+vw�a��%�\�bk�>��[�m��5�]�i��U���Ti�&�6Y��򫍶ݏ�d��itm�8b��Ԇ����[r£'~B󃢨Bx�z4����nE�^/��/x�Y7Q�qP��
��,�SH�Ew�D�E�Y��+B�	��ڌ��'�����%ؖ|Eb�A�T(z��3�W��Ĕ|�\�AM ���1vbz�H��'t�xʦJp�4��fx��="�"�T���L����"���h�9G�S%_�Ө�LZ�p�����G���ϼ�l��i���2��  ��IDAT��{���'��.��ϴq�)>�(H>whn>MadN�==0b>˔�}ԍ6W���UqÃ����-y𧫛�L�r=F���>y�$O�F������Z�����lck��b��zݮ.�ث�^���������={������޷�u��oܰ?�����7n�w߻k_�}������?���֫����/���;���U[��l�3j�Ę­����P���~:�N��ԍ��/Ə�TDN«���J�����8k_8�c�H��<�$)���Ydچ���O�6>6�k7ph��o���6�����t"�G�0\��7�ц�O�}�#sn�D��j�G������c����;��Fz��;���#��)SB=EuLX�Ѯ��V�%�;;�_6�7�fRq��1"s�)�hJ"RHA[� � u߳����抛2}!�S��>�<��ʛ�E�2����(�E�(ņ9�eI� @�d����1��b��q��c�8�$qM��S��IW�°cA#�wد�Oq|L��$���@	A ;1�`D���[�00�h�=���%�4"�2^�� �
�?���u�'i��Q�`(�[��}8`F��/��3�uf��&�w�]��1�签/��2�7�τ'N-�0��+�B�DC����apP�r���<�E�q�r��`f����������/���h����}�IC��w^�����٪h�-f��"M���gbƶE����Q�ִ�h����J�ϙ6�O�2f�h�u�ƞ� a���@ļʷ�ڳ��Us]�[�/<i��5km�s�����c��f�k^0�Ԧ�\4���k�9'�?���yO0�'�cSv��m�޳����핫�̹֭�7"}�'S��o�%V���S���`�>�Rզ,✘����=5��ˎ���<k����)[`Ju�r�&�ڡ�4\:�Qf��$G�q�To��w� 3��Y�
&p�']����_b�}!y ���-=��eL&'���y1T^���
�=)��ľ�����0 B #� 	D�0�#N���C����5�V.���gg��Ṓ��C&����a�dj�"^��`C`,��{#���ҳ��+^D�)R�;�O���0��Tf\��+�t�@�wV�y)����G7����5�s�'�"Fz�z��=}��Ջ��3x����9c<��^�����}���?��?�o|�M�m�AK5�3?���[�P{��V�o���5FƭU�ԳI���[S�;M����d&qDcmF�F\.K������FCf�UT��-d<PGђ��ow�M0�/�Y5���.���S��!��Jܴ�g���q��\T��+>C�^��p�@e��vbЖp��&�`q@�<�|r����Q���D���V�E�����w��/ �![$�KB!U��kN�"@!:2s�q0��=c�0)P��FO�ȵ_ȉ%; ��ČM^�JQ��s��)�i����ȟ��I��59*�0<1Hr�CS�(��/�0����7[��B�0�ϳàx܇��)$��VI`�.҅V��z]q�냚Y�D8��3�癅�V�{\p�w��G���i#�xtA,���#M��CH��'�Q���H0�Ee׬ .�Oߓ���U?��Ǖ�|�(<�C���ҫ�����w�Ͼ�����z3C���fX�^��qL7C�BSQu���iy�Wf�����L�>�8ߧa�!@��ъyPCw;�Ӭ�/rc2@�ԅ����&"�w���(/��.��Wh6h�=��v0��`�J�,2Ὅ���� �ޓ��;�/sY:w
D�=�.Y�q�f��]�>��%!��D X��TK���,^�!�@N��%5��B�
��"���_	Q
�~j�����#0�	�R_*�z-�/���,�U�R�|�{Vq���Q	�q�2O���*��#G�����D�M>I��ޏt\�&iHO �$Ř
�"�޸�}B)�E�'`�S�)����``�z$���<��^��֣��DzҒ'u	�]����޼���L_����߸���������h�Pg�wv��}|Eii�x'�a����B��7�O����o��}�������,W��{f$(�17i=i6��f{s����AaT���Y@At���q����Y��y��,3��u�u_�V�C�,�dHO��3m���#����ޢM%T��fѾ��Q��}���ù�n\H�)�s�w��%<��"O��"��������I���g���^�9}9�$&&S�6V��Z����D$���}�L�#��>�sE��1!��~��j��A۪M��w䷭�۴���U�[�o�YYa#�u	�=�w��t?�XW���v��۶�Ѷ��z�Q	�����aT��D��&b�q!�j�&iC�K8	MO����'6�sD���	����С ;�'΅@���)�Ԏ8�'�S�玄�|��z��n��t�Lϩ>	�.����Y	�!N�}���<o�:��N9.�uO}R=�2=���I�����z{�,͖��_���?��ٛ��O�*��g�6��2� �KjrN�
�pQ�!0�^��3���s��Ln��S��RR�)�%@�j_B	>��g��Te�L�;�U6{Xk�.#�N#!-�~Է��]S�\�O�����іL�F��B��q4�E��~���WX�	op@�ǋv ���Ĥ��~��ی����8�)�
w�W��@���4X���iJE��
)L�	A܂X-���n�ڶ��͕�P���6Ҵ��=xrڞ�t�N/��L-��©Y�xf��̏۱ɂM�;���(��R�� "1.u����և�&G��B�'׸�Jx�B��}r!,�!q0.�%a��:*l!$�0�z#RPW�)|�+�@���'q7���e����p�<~�y4��Ô��{Da��$}����)��P��<��8~�p�~��4���A��#7��cֈ�}{���
��H��햭n����h��*����
<�:�`d�R,��#9������ЩS��3pl��Y䳟g�$�ʣ�UL$Љ�)@�VIxA$�;~��4�o|0��w�|-�	J7��`�{�\�&\����6 �h?%�%O�)����~N�������h���I�gg���a�����o������k�F����ٙ��;��̖0+S�ST�����m�vG���﫪��J��kL�س�<j�_:g�^4z�!�&'��{�cղvsc�+�=�)`/���~����ǯ�n�M�YƂ85�"�t*A�h�mc��*Fgw��0���+E�_��A4FMy -�eW�i!9�Ǖ�@0.���.̣xN��2p�`~�sf�7ze80��#>�D��9��|r�uX3Xp���Qw4-����[,gO���M��;� q�������$Hꭞ*�)���>��(_E�}�2�Ge.0�� #2[Y�-]5,�;��8.�{xE�P^����p�r�~�m=�q	=�쫜���C�2�V���t�61f{�m	��^��ڲ�=��b�
�
&9f
(;�쪑:Ҳ����$EA��5����JM;wb�~�ŧm<߷�囂5��q�89�C�P_b��p̂��"�����i���y;}梯���7}vf/7a�m�^S�H, e� ��E���I�����yF��OL��Eku�[�11^������W��`O��� �:���p�y�z ��+�i�,q�����d�0�U�&��H	ĨA|ui��;6=Q��}���/����/����O����ů�3Ͼ`��hթ9�;}�x�q[<���>p��^���gmb���f�[y|ZP��}�)�JL�`�j����m����}ܓ.��OLe���"<�c|�q��8=r��La��Q� \�S�ۿ��q�G����ꑜ��Ļ�'�&�#�<���Ǻ��Ќk*�;A𑭗�)��'�q��e��ӧ9� @lz4��X]���-7�+��m+4����d.|"Sr�:�s&����ͽi,M;j��s�JF;V���x�&�$P1ݕGI��@�с�0"�J��I(/ڹ�L�.|o��Bi���x��df��+.p��=�t��+�)�D�`Ը�����L�e�	甁9����3�o�H|�I�#�#/IŢ����yg�޾�a���?�kw�$�V�楹H�K�Ā�嫶'm��mK�yE�9>��ԈO>�����5{��i,��;W��?�����HJmzv�66�����h��	�Qk��R�z�z3�5�~���p�V5'Ev�i��-�!��#Ū���V�Z"6d�pN���@d�����4��HB�b�
� !�I�"c-��ʌ�k���)"=���4�_�(3�1���>�����9�<�G�����h%�4E�����i�8f��cV?��c�'X}�R��2�r?I9諬Q�����N��P���k|JuęaqV��O�	{�G}��׿�=��w^�M�=�֒f�~ه5�4�Ξ��,�?�������5;�8i?��w��bKҼ9��U��hq/fn�eӃ��Eu0#�6i)�Ѿ=�0a_|�!�����J��>s�-��	�NKY�-)p#�*y/���
9$h�N�<'1X���|�~��k�g�'m"��,����LS+,��a��=l�C �Q��z_�6;�U�8��W����|�..V}-�/���f�-^rS���!	�>~�s��5:]�qg�������QIc��CR��7E��5{�)�h|��Zs�n޽k[4�ڌ��B�y�G�����������U?�emm��-�J�ܵ����`m	-��f-���/d��L9�r��E�� g6r��	2�*�`ɕ|#fj���g�KLM��\�Z�QX##	�x����Q&J�K�e�n�޵�����I�%<~U��"��s�������fԋ���m�hM�þ��HG\�/��y�M���YSG'�LU�? �r�&�ӕ)��~�NM�g?����_��}�s����'��S6�p�~����#�g9>͠�TTEVIcB�L~oo�~�W�j��?�;6[+��Sǥ�Ĺ�-�;m2	�4��v��T0s/���UFQ<2Q-�ɹ)�(l��P�b��t�V�I<�n^~��xOYL+���[q�D�6�B��҆]�[���%�=&�k�2�b������p�+�)��Љ�R*�����瞸h�Ѽ��;�����xp��by���h$H=0=qQk���Q!�Kv�r�`����:�����w��������u�mk��V��/�\���i�R���_+���S��T��vTĠF�,a/��m�"QF�Q���>N���D
rCX�L���+(#N��I��jʶo�f�x�M|�	�p�駴�,/Gy���r)?<�R��������8|	L��u,�F'\���<�z�+\�p�C�!��2X�s{��sB��@�҂�(S/?������͌�?�����͟��:c�b۶�����]{��[� �&�T�ZU���ھAt�4.��q#vwe������^���}�������}�����㘄G]�c<ϧ\�Ρ��u������-�ۈ��8�:g�H�g	V44qY���Y�=���H�8�������=� ��q�r;���Oqȗ��hk�c� ���P� �\@���2&&'mjz�UW?�'+D���W� 82��D�h,B��4M�L�����-�ޟ���]�lE�F�&=�R�2�ݵ�ޚ�[j�ۻj�����5|�>XO���dT��-5��PA�qR�XmH���O�F>1eB6��w'й�F�w���òH�#<~⽧!�xfJ��&�$Ϡ��m�'=H<����/�N0�R��y�] F��ë����	���uԳ�J����u��dT:��Y�@7����0>ab���U�L75鄄��i!�49>2�/�E� '���<_J ��롲����CvJ�y�&��d:O���˿����Ͻ`��S���������_ް����O���ץ�֕][t�#��';i�t�N�m����5�g��{�ږmw������=��%�xl�F�6ڒ�0 +h��
�?-�gK��<8�$�,�Y���Y,S��>�&�'k3������UB�Do��{�ǲ�W'|p�U]�J"�;s�K��<���M8W�%��j���b��^�7x�?S�~:���] N�����!Tx�@m~5w�F�J#�eqz!���\�(oOW2M���rV�1�\�9�g��Q[�����=tb�;}�<�h�]:k/<rξ��E����\8e/>�=}�M�L�Mټ2Q$���D`Q���t;PO~R���%S�����Pg`|�5]��F�#5*�6��Ϡ)�����G8��,�a�b��O_x��IC���i�=����Ǉ�C@I@
�w��{��U�~�5�x��F&�XyNx��}A�C,�\�B�=L�+�A��Cxa*����"�'�1�~�X	<��)�nl;���g��0
B�&y��r�\�	S^�0g+�����K_x�jE�W�k��?�ُ���؟��#[��Z�:��e掶�Ft�z
��u��Z�J���ڷo�����?�����ukts~jؔT�/>�������I Qu�1��M47	P�KE2!�U[���_Z ~�g�E��}?����A�2G�"���~Bف�=k?"��X,�H!��#�������s�-��a���8*�U�y	z���y�Έ�ᘈ7h��Sb54�޽U�m6my�a�_�c�����=/���%�u�Ry��YC�H&KcUI;1����`�W�~�����8oO=��=���◞�g^x�~��=��c��W�`Ͼ��=���67?㒰��'�	q*�1q�S3*�/�V8ҚՄ쒜���A.�e�6�L�聁�@H��AC`�oҸE��\�S� \����la� !�H���+���p���W�A�'!�GX�?ʊ:uD!nrIhN�T��7�!`xG��#��!��rb�o�b�!�8<8/��dT��R�	 �+���=�"�op�~E�<��Ia�2 ��c��g�o�l���w~���[���m5��#e����#��N�rFG9�lE�ǫ�:�I��D�6�	��lo{��걱��K9;��i[�\��7o
�w#C�F������9
w�r�Pg�>�?c�����Sۥ�H�\rN����)����@41a��Ą����Zݱ{[Mi�D9��X��>4����-چ<SӒ#V-��_<֏:��'<eO?zΪ�X�fh�d��r�9���=-y�`���L��*`�O��;2��Y1���iv԰]���O_���=d�ϝ�cg���cV;6o	����k��p5��씽����^|�&�<��*�SBTr	�N�z�
6�E�A>1�s�"8��ϯ~O�Ta >�kʛ;���2����g���,=����p�]���S[k�K��;�	L�B�c� zF �SG��3�ǃ������"?_\�v�#	+ 
,��q�y��G�r!K=�e[&��W�~O��]d�9B��g9����%��@�;PbP�(���۷��V���k~���x!��8����빧-UG�X�nWј9��ތ�J�~��}�;ߵ�zݪ�q��=wZy7e!E�Ԣ��JM�z�@{��]�b �("	�#��I�x������+�!]��x�K���½��e� ֽ �|�V3�w��x($��JY��WZHpY�������\��9�fw�g� #�
��3��sU3s���Vļ�÷5*����}��i��?����|�^��j?x��}덛��Wo��޺g�}�e�Vo�����J�����g��<d#�=�&�S��N�,���B��A���ddݧ�?��#�[�a~ �6������t����#0iԗ�x����G��:�A���1��(��D(����8�!|r��w�����!$o��fyd�Å�ųÖ	l���=A�N\2�.Ng�2�E�*�0�s�h����)V��B`�=�a�I3KCx�f�N�ը;���2.��������	��V�=`��0=9nR:�]�\]�1*�v���!�M.�O�1ć�+{.y�
瑯�åiF�a��}%��#�!���8Oƽ¸�D�6�̀h%mC@�O���?���^��K\�*X�Н��/��.f+��+{�h���ö������B�A.5��`���X~���&k*�LL����k�ۿ��g�����O�k�ۿ���ۿ�M�������?��~׾����7�Wߵ�n�ffge�|�.\:��&Ĺj��;�i�(Z��3�C�qC�G�`�&�7��.��CX��H�P=b�Bx�@x�0@�@��\�3&B>a^�Q���(r�9 �M����=I�8q)/�=����R�#<9�Ϟ�.у��l�!dʉ{wJLG��E�A�R
�<�{��V糕𘐾�D8M�:m)^-I�g!~�I�a�F�`L(�� �Ѣge���^&k2_z��z��U�k,Z���ک,�)�a����ej��+��tU����^�I�:?������T�n�g+��V�N*�4��c�^��:�Ä	�!��7�����3����z���<�N�!D�]��ar���"�;�#�p��?�-�{� �q�i#�X��h�S��GN��sr�}��R2�%��������G��n��|&�'��0o�N�26��zoe�./mٝ��ml��Ɔ���ݾ�f7�N����G��5��׾m�k[V�Jy��);q��#x(��R2X��{����%�H&1N�A�8>C����@^b�`�h�!���抏��rh$x��*��1o��}�9K���p)$��_g.� EK���G뗄����~Nh�C����E$a�����Ꮥ�	�1z�?�z�$������	��Ιȅ���!x9P������������W�����Ǭ��l�\ˊ�m+���4`��c�����ۖ�o�����t�0ړ�ұ��5�l,��e�{?�e������ժ~N�k��io���5��]a�5�g����FB�k9����WBcVKu�^�QƘ܋�mD3�!��t��\����Y+o�G<��NAn^fϴcDփ�|��<m��A]�]�"�+�����&#��>Y�R�����/�`�ωE*6�O�a0'��+���Ow��(�~ۯ������xE���w�|9�|����m�|�n3#��Xڱ�3];1Ѳ���v˪��J4\�v:���R�>��2h(��`O�Ax>�!�A"uI��ʝ.	����AĘ<��P7p04�B%��4n�3���yޑV\�s(X�a�f�s�Q�	v�r#�¥|��%/½�rX�pXw�\/�~�#����{���ا!�:��dr�4�G��B�D*��`��{�������+7nٵ{6R���O=���ݿ�+��#gm�:��}�+�lbt��l�����g#u����H�NO��|;��%���W��~�o��dMmq`w׶���K���]��|�s��pY�:�ր���\����f�?�k�W���m����I3&��(O��1"τ|�n�ȇt\=Op&�q���ئ�T�����뱀X�i��S�Q/`�JHxt'�6�;0�����#���ʽ������]��a��ZS�rbN{WnS�1�ݮ�)�	R��o��j�U>&��a��/إS�\��C��b2lΒz�����т_�nX�7�3����� ����׿�#۬�
	���L?���ґ��qF��R_�RSل$UHf�Ϡ�u���� �0@{���Fť�q4)(T��0�k0T��)�Ǌ�Ty�'<�".�Rø)�Cb�#O␞������]��w�"=Z'|��p~
��TQt��#�fff\Hb����FS�\��ؼu���r��h�Gk�C�>~��.��oBF�0V�*[��CF�<n]q	�^W�/��������`�S%7e
#[��lKח$�djɄn�[�ҕ΅7������&&�҅�V�)T��<=1�x�ַ���������5ۨKk�T~-)0{~l ��GY~�щy�:���������h�^�ƺ�G-
�TGݼ3���Q�i���2���x�u�͔�Q}�*��♳V���?�����/ۀ#*{�V���Xj����a����`�[�w !!�K�-r��%kD˃Q[���_��G�׿��]8�w�S��T8�t(D�� �q�p��Ǝ���e?��å]	���M�KP�bE����&�e�P��n��]�\:�]	������x�~������=g����K�h{��gǏO�Ԕ����u:#�h��
2ET��_{�~���a7n��~Iv0��	BD��I���Y�_��r��b;�4q�.U?*D��������H������ ȇ0�3	�az�Ia����w�^S�G��>	�#^hz����B�"�ϑ'u%�TN�9��:��n�n�
�yi�����e5d�1�Ֆy�G�GJ3"���F%Dİ]a�o��5�.ą��أ/�=�(�������E�0CB��{�yTʣ����_�	rjq�͕i�]U�Z���~�m�{*����;�N�n�"���gi1lȣ�L�����W�٫��m/���ݸ}Ϗ`��Y�VL�*3��|��
���*�ϧO�]��Y���,Z}���TW:� oD���)j:�M�asus2���r�8-R�:�\IpN�t�f�1jS��׮ڷ_�b�✵
(D���8��q��J7�����m�Z��$į��V���^G�8�ۉ�i��/^�����s��^�v�؉��FA����T����2>���a�!u�!1 �ב�*�Fz������'Nرc���������Yyr�J�36:6m�¸T�q�O,Znl��A��������[]߶<�,�>���(�6u6۹�u�ȉA§��&����',����w)_�Jq� y�xtLh/3%̤0�\/��KeR�����x]�U��!�G��>�'��I�d9r�]�+���K)�cUkQ=9��(�˂	T�3J�D@�2�9����>��§�b����k����եM1��wtt~�r�
RŅM��]�S�eieu0l$U��LV�Yq|�6=��������k�i w��$8�bX��g6�ݎ�;�m�������5��]@Oj��*G��v��v�3�+آ�^?ц���Y}�����(>8�+��~h,8��0��Eՙ�=��ؠ!�B���(�@���Ь�8P�z0e��	��$w��Lq�4��z��O�Z�޲���S�����M��0��P������Yd��FSƕ�L�j��G��ٶ5I���k��lٷ�ܴ7>�e�\�c7V��x�۫l��Ɔ���W�xϾ�ҏ����*��F�k^��p �4�P�,`h5���N]��
)����>k�a ���h�I�(�
�s(,>�Gs}�c,%�|�OG�$!cFY�A�F�pC���Bs�a��?�����]�ɜ^{q&P�m^�-�{�z�2>8ͷa:R�Y��weh/�A݇�`���?y���]����u��X�6�}�aH�]�~�n޺c뛻v��=����	�����{7��-+f��|YQ���մ�K��������n��f�o�ҝ51dٗ '�$�F%��ML��y��_��f�]N������i�j���M��ĸ�eF8b��(x�Y������C�h^�hԣ�5*���L��Uj�e[�jۭ�mk�ON�x���&:dO�O>d?�����g}�xk��kh8�\��sR?*9���ɓ�{�Ξ���J�:���+3VpxPΉ�QRV������u{��-W������|�v�OF�����/� �Bt�� $�@c�"�(|ImӏߗY#�Be쩷R��rV� AD-��m�0U��JA�U��h}��z�`��5���.e9+�^!RR��R�Zj����3#�!��#�%�<,�%D������!�`,�ӈA30;�C��=�C`SS��G �y�t	.`r!��4 G~�EO.�	>��S�"r�Dt�Ɖz�;�Eo����aL�x��B����#O����v�V���%���	ɳj���@A"V�O��U1! *���eWj�s��tԜ��cLm�-�S����3�;5^�Ņ){��'����m~f�Cq�Ƥ�.,Vm��n�����G?z��.��^�.h��zcE�:��@�@6����;������=��%���g��Z��k�,��[��;سse{��3v�Ԃ56WE߻�T|�<S_d~1��
,��kn�^o����s&7"<
YUu��b�4�7�oٟ��#[f�K�&(��\<�G������������O����^z����GvoG|R����<�Q��vSB�\��}�~��S�����cU�tU��5Dh" K]���"�D�z�Vפ�䋶�ݲ��,�^Kbb�D͋ȕ��8�6�t���Ⴡl���q����ב�!Bd�	��N[5n�i���֔�`f�����ɔ,�Bg�Z�Y �a�DM$����ΝH�g��|��Ј�`p�#���<$�y��I�˂�=�yG^�/��j�xZ����q�S�:&��+)^!�(K�,���XDh+h-�a��?�#�D�������}�I���g��+�*#<��=�ظ��!Xٟ�"��������c�7�+k��g����D��T��G1	�^f'��Q	��̔j�e��)�ӫ�^����ڶ]_ٰW޿b/�}�~��G���~`]�g�}�}�;?�o|��:�E|�	�,1���	�P�$��4w�#�p��/��o؉�9+������5�h�>ЪJ��m�V�Ei"�洵}NC;`@��S����r/O���!��lhc�������/��Tj��L����ݸ�e{b����H�?C��U�+/>oO?x��+��&e������;�|�OZ��	m�U1^���Y;�8&?e��"C,���:m��D@~��_ћ�S�a"�����C=�<,Бu<s?���)M�'���>+}N>g�f�}k6�*+~"�����`-i���A�Ttx�z�0�<o�$z@`A��|0RA4tb>�L~��sϘ�%L�Ua8��I��.���8�f�w<�M8��i�1�v��Ub�a�!� 8�	^|�'��F=#`�^U���n�W�9��b^6U*[���ë<%J�-����VHYF]P;����F"C�|���<_s!��'�e+|x�;�5:����M5ICx�7Z������҂���dr���Zݖ�l؝۫�twծ�Z���y�>������$����`-���ћ F�i�5;�[)U������MNO�#�=l3��m�m�/��K��4*S�½4�������:D:E�i�':�q���Q:���+���:⏮<�[����{�0\�#O�m&|�XD&�P��]��n�x
L�'3���d��er1�����%�P���oW8��qp�G�9�@�����lh�`��֔WB1�9Q�0>RN}�7*'Y3}��{N��"!5��X�Ov�P�V*��[^ ��#��PU��,�.� � �"��>��Qk�]r�`�=_�#�9CQ����)[��?	KWny�T# �(�Ï{��2�M�|R:��A���$�������	����q0'B�J�ဋ�N��s�f�������s� qMF�ք� *�E!<���)�m8YLؓ6��s��@3��a��"��P� {V�~u���ք8])>~ �tT&�|���SjV�2&�vS�)ǥeT0�E[��iU�'�^1�/F�n��`]����!���]��F_`�Ǧ:
@c��g^�\�C��֐�Ǿ*��s�JS+VjV,�[yl�&f���)[8~�N�y�N�=k'N���c�|̣T�YI�
�8�2:╖Ϟ귋0�����P<	4�>��h�(��pTf��������H�{�z �Ú����v���T�H���5xj0�sF�BMX� H5� qU�{Z�a�`�=�0?���8����3��Xc����+"]�R8q�i�����Q�x���N��{�ͰT- ����C�\xs��n:� B����=�PF�heL)i�~�!	�(+4�pѶ�q��Kur畋[�����0��)�OHWY1���Y�p�����#�����������:O�r䔞HJ���e1�ٗ��*mR�0B,���=*?[Ƭ������.O��`��>j'�/>��=�ܗ���}�{�K���_��u}���#�ڥ�>g�<��=�}��E���=��/�S��~�i;~��;y�f$��$3jcU	�7�"P�M�]�	���h�8�u�O��G\�c�s{{����3�*9����B$�nc�*v:_���R
�=W��h���a��7��P>���:�0�?y2���#���k��U��Y�2���2�Ki)���L���g�a *�!B(�0[`6pLY�G�H�8�A�H�2z�������"�=�q��D)	�h7�J8Z:��9�t��Ӄ?�5|�A}xGZfB3
ܤ��zH9�wI.���F.�Ou������R]���^h���sQ������R9���!�"Z���y\mWm�la�=����_q�p�̃6{��,�����6>s�Ʀ�[ebAҧ&-aܧ���Vu��K�L��O����v���v�����g?o?��_���Sv��%;q���ƫ��D�҄dr��r�{,bS�&��!
"͂?��������ݳ��o��S;gw?!D�#
t�г�NQ@���z��"�Lբ����.#��cy8�;��ݙ.���@ިk07��`�`
��dO>��"1$�g��!��MZF�	�{����<�'�9�>R$�ɵ�e�1f������4~h\���0y^t��+��!����g���
�a�I�ҳ�"O�x�(��"u����6����O��;z�#6L#�0$�1FV�GuPZ�Dh��s\�:3;m�������bb��S�Rv�aLZmb�N�:g�=���=��զ�8>c�ʤ��j��N�y�׶l�ud����N��Aa�Z2I��L�)^�h���vٗ�q��Y{�g졇���).S*g㕒���%ؒ6�F�[+T'�1:�Wֹ82�����q�!4�@�ы�[$���� Z��#���2�E��8��t)�8ʋ2?��'����3�����+=G5�V�g�D�I`B�i��q��$_��@6�����!�g�8�8��!X�0��e�O$���m�NB�įwo
y)�G����h���=�����:��K�-ס	��6l�t����]�����a�%�S]�ϊ�?$�C\}�,�	�>�K�Sc�1�H�X�o�f�q �H��NډSg�!�݆5���~1�Նf`�ʘ�k�lt=�L��Ꝿ��$b��~^�M��+PY~�Q��2Y���9Ru�CS���v9o?�^� ?�$#�blQ�P8�w����0-5���(n]���@R�����q��:���pÌ�S��@J�_��X�#)u4/��Gb,�@�����&D!p�#h/�h�GkIB�<���H�I&�>&1�C���!�C0)χ9+�&-
3G�q��D�\	K0!��x2��<q���� ,�ɋz�x��[W\���'���z�6!X�c��*�eO�K�
8:E�x̞�5�ӶY��i��l5lks�vvwԛI>�BDBC��T%\jJg���#�P�����d�Z��ԭ��5T�N�'�X��u��9˂�\�7��Ϫ��zK��39��քU�|�%@5�6"����0�,�-Fg��D��|�z�
>��[�9�A��_��s�I	���Y�*��wJxMwQpjX����X�)�~��>Ɛ^��Qb��9D�%��]����q�'_��u�+�c�p�aL��8�\�dp�\�:�$M��}��PSO�!�3a�\*+	Za�K��i`b5p�B���6�G�j-�]��I���0�?t�pz(ݑW�c8HLzz.�BW�B	G����a��v��&H%�ϟ����Q�[����	^�a��ӹʎ�H�G�9��w AW��^pSM�sS�^���}%~f*�Q�Hnp�^�W�"h(�-h,|d�����\�[�YT��bMx�Bsi �{����'��/Y�+U��وʔh�b�Mw�  �$8�H��Ԏ8p',9"�E+�����w�I�I�{�c�2|��Y���Ӵ&5 .�%���L!�[�P�Tp���:� �KD�yL�r�9c��<��r�މ\ϩ���ȇ{zu���} Yp�ž.����x�!�FCو��y�CXh%�S����-c|1�_����1.�k�<BK��81��Iz� Cxx��oݥ��e*7�*��L�|��pq��F�tƀ���u�M��	�q�y~�*w�y��;��6=���;�K��y�C�:���^��@�G��GRp-T���d�����<~����|P� ��h�m�7���4�mi/-��X8���@��rx�8���� @�j>�
���N���K�0ݨ�Y��A�4���aΰ�Șf��A��R�������X�T|�6�ߠ���Qw�ONy�Q;cu���wA�����1��;W1�)1�ե�D�OF�0�<���q ���>�&�7�X��y!%"�Ȏ!ɧ^��A8�����1�D�W0I��y:O����`�0A�z�r���L�o�Ð1.�L�$T�^��	@�y����|V���<�W���K�	>�g�-�Ï��+9����i�Sf��귟�p�J,�SV������;G�B~Kۊ)u��G/KV� �Wf��V����Ib����s��n}�V7V�.��^��TzfU�8��o���r�(FK�mI���A_0��/Zӵ�2�E�ME�R��ࡍ�2�TX�Y�b4̜�=��c�&¯*��A]��MC��6�δ�p���z=���t��s!�0_;#���U(�b�dEAdDa�LbF���tM���/#��i.�I����t�U<�qDI�����0���#�xH���c�����"B�.9�AHN��p�6�F����4�$D"o�^����a%ar���_r��GVY	/x޻p�<��}b��u��rRY�U���?ɑ���G*7?R��;�!?��!��{{g_�Օ���I*�J�"��U+��\���Bd�����pfo5��>Ą]���I�ٱ�^K�m��nX����m�C�o������DB�L�����J3a)}h�-�����L
�5�S��c!�h���H?�#����L��9��g�(o��AO��+�p�&����N>l]�;ATz��_��x�G�d���'8��Tm�3p%���v�����f
��Đ%����ȉ�I��OZ�w��g�@<e%M$*ϕ��*I;�S�6����ܻ��Ӓ�0����$K�{����E�=1|��;�}����6	��g*�=��/{��\=�Ow�����>;�_��ua��	8~�%���Ѭ�~Ą�MG;55e��S>cCۨ5��r,ǔi����4�]�	"��Ɔ$�� ����m���;z�xz�h�>%��`R�d��zaZ�[M[�w��V�e�@/08JZx2�Eg*�Ed�V�雄>�#���sL1��a�$�	e�H�%0���P�tI&�A �?�"�?�9�p� I����Ow���_���E��pQސ�AF\#$z�Jp�)�	��5K���(�?�g&���rN�rC��-��Z�D!8�=�G]���~�yN��q��Y�D0�|��w��Qx�n��a�H��aTbh�y�+�J�hܸD,�?������%7��3��?�y�q{x���P	��S��GY�������8��bf���_NzgO��檭m�����!d�k·mƫ�ǾƦ:���ó���d��8�#N��LY��{��]�zծ^�����+��|OBCy����bF�5Pa�I�^��W��!�:�O#O��J��Dע/\���kty�)m�����B(��rC�!ǣ����� 4+/+��(�)|ދ2U0u�������T��3��e��"!<�q�φo8f0t��h㥼#,�S<�+�/�C%���|���'�ƥ��~�č���Q�p�6�nfg8���%�iNo���g�G�g8��`��E�"��#��q�!e��ue뉦�g|�Sӳ�#��^*�U�{��mfnZBa��7����]��ް���5�u����5v�!M�#D7��e��ٮ��͝�ݞү�\!>G=ʼ�ys��=[YYq�ON�lLBb@�&��J��$~��	�<�ZB{�'<z}���Ak�)i\8���vNb�=Y#���)��c��MJid�+��)�nO��x�z
Ob�*����0*�z7��9�'F���T!=���)�R�� �Eֲ�XBN���o�"v>/x�L�g.��3�@	��3����H��w�j ��:����� .X��@ <���0	���,�����3�W�x�G�b�x��%z)�*3z6���B�"���xNl�r�0�9|�U^��S_epH/_tC�0��uUZ�����%'z��lJ�i��*s�,��G9��.aC�n� ��w�z��h ����R0�p4�@�pjPE�rN���������i�78ԟ\ �p�ﲀ`	z�C|*�8VVդ���J[���rmDV([���W����}�s��sO>c�>�������mە��w��L�[����M��NӶ$l6�W�^&�̙]i(;���o蛝��csv�؜�?w�}�a{��g���_�ǟx�W���=��`�����8�&_��K"�n1]-A��J��
Kj]Y��y���(!0��7�S�b��0���a��l1�˄a�G�y�w%�X�1�OE/!�P�x`BL0� )����b���Q�)�*�4T�![��@�)Z\y΋0FU��@� at;w te���J*�o��u/&)s�{TL�Ì����RX�qT�<\nP/�!QG��(�_ 5"LW=�a<���v*�˔��-���veĜk�z�i:9�&��wVaj�J+��������j���H�\{p� �la��6�9(�	�Aኋ��=��;*�sz]V&�2�ΡD�o�)r�ʴѾWa��M*2xWC����ؗaGo���*u6F��;�	! �9p�UZ1
g�C_�ˌC�ӑ ��&S��ٱ-���`\��`SHz�=�q�UɁ��6>�}���Fx��M& �Ct�f��Hߪ2Gf&'majV�f	�l�T�������������=b_|�8�`�O��z�f'ln�f�1uҪ�X�`|�rzb��%pN;f��>`Ξ�sg�ԱI;渝�=��9�җ>o�}�I����)iG�Ν�y4��4#�|0'��ӛPե�/��>.7�{ږ�X�C��Y�ɯz��J	'�Im66^��#�	n@��kz�Rud�:+bR\Te$;�hHso�H�)�'�f��)�<��Gͧ��W�����b�s��Ud�+>ΤP:�u�sM���T�r����T7	���j_���J�S�ʁ4����+- CT��%��#��C�x�]��X�7����'OW�0�$��;� T��-Փu b��k���վ�ė�	�:�t��z�.�Av�T� ��IH��e	���cԻѩ@�Gp�0*@�����|�F!�2 ��b�g�	�G���=��C��RE�Kep���^WJ���)��|W��	W1�>�p�\R١}Gū��G��ȡ����� �!hńu��֒�AϏ�B�w����	kI�j�i�[8c��Y˗$<&�m��i����	�8~�<e��lvq�ffmzn�&�615oc����jmʏ_hwebЌtJ��<y�Qv8�Qu Vp� s=4,<uԳ�9
��~YPW�En$TG���/2q	�|:��F
'�X�, �(r�@�b�D��{c���ǟ;�
�͑x ���$U��zH�ͅ��縂��<'�0�ה��?=���$D$k��_p�9ԥgF�'���ŉj<����i�U?�����+�"�`T ICpd^�OϪ
���R_\�+=����7��l�	���ؓ���K��m ��4�?��Q|L8it��HW�w�N�dT=���F��ȏ"2��4���Ę���FO����EC;�y�{N#��aB�A�.���x�J�A�@W�H/�p����9cp��A�ӵ?�(8�>��whx��8��6�qe� �a�a���3�Vo�Ec��I?Izkw�^��Ĵ�e�MNYilL4,���wRԳBY��$����0,"�|���M�;?��2G�Q�{�p�S�ز���K�B$���O��L_�_�� ���漲���.d���6���,��EJ\<Ī[�	���^\�dy�^`8��v��}��4�"����̡6���H��^% }010$�@���#C���H������f��xp3���9KB�����J���ί��Uk���
������Y�{ɅJ���v����JD�`���Ui���+L�)T�J���]���� `́�죥�~_�.�ف�����������|&AŃY��g��uI��j�x�0�p�Yؑ���U^6�����;2����z�p%��RG;1]D�x�C�\#<9fG0�Y�833k�O��i�̠��T^���m�w�k+|����%{�w�νU�3i�6�xBBeL��(�Q:L�l�/V��åw�:���c+k[���m�{�'�$Q��ls�訕�1� B)U��3yڒ�I���5��3�8B�$素|�"r @D�#1��	g�<`'O�t-��%�|��]�1<��0E�'�����፼7�!2��W�44�_�@qKP���9�*)u���k�D ��0��\�@��A8ʢ�8� �g�U�]�F���J����j1`�5J�<L�z�Y�>�:�����<+�� ��V��F@>���AW�D�Ս�MiUWaY�Q����	�N�*�}� XB�D�C��7��1�Fshr�B���Z��t�js3�1:nEqnIp��p���*L͵��:���s^R��������0�W2_&L��K�޿����y_<�N-��Ɯ�)�u9��D>i����i�Gx�5��x0C�=i�R��Q��شkׯ�m	���5]o��o�n_����[���ݕ�)3�Y(���{.++�V��D���$UN��z�ի7�7޲��~ϖ�ܵ�][Ww�޳�K+voE�	��+��s�J��� ̖�{�+<t6��!pr��5Q��h#���9�����5�H�B��_dt��?��1���N�w!�$�b�oHs�_ċ'DВ�TL��W�`� t����{�9QP_�Eo���d+��[��������LB�#0pfW�&�$�-a,�K˖'��Y!�c>|M��o��zc����iUJ��E���y�tm�n���=3(����N�3BI�D(��	]���K���}�@�����ݴA��eq>�5}���w$��q߁�{uB���ے@��a9�z��i�nǯ|�_#\�Yvm�A�e�bV�%�/x���:�w���%�]�Y���c��];�#i2�ynnl؞�����@�Ѹg�y#<yK�xOӼ㵚
�x���4���Ҥ�/~&�p���VKB����]i+Sv��V��lue��|��я~`����}����$!�|o�"�5�y,�Z��^��]��延����|�i�RQm|`w����Ғ5�T�nϯ��t�,��!4/у���t1K]�(�ipŁ��s�cg����NM.�߹��#�YQ�n/ݶݝ@8�����!��P)}�^����qG8q",L�h�`yL���Uyy�v)(8�=a#3-�WN�O���G�~|`܇$�(�b��H�}κbP6G��08N)��TB�|W��y�1;?T-���39���3�UL
Ç0Qo��p=��C��	gj�5����hU,g���q�]Q�JO��sbP<8������*�)$4�-�)�qA,�@�M����u�Ixt�b��:�8�~`;ۻ�����-y�S���:=�0���m{�k�~O�/:j����q������z&�E��������>{n��s��̞um�|�ޯz�Qy��=k+��;V��}��욂y���x-$�iS>'��)�5�	���L��]�H��Mg�Ν=cO?�}�K/�>����I[[�ݸnk+�ޠe���9Y��g+
��b&�3����M����ر����ab�W�b�R�V�a�D�NNY�x�(���#Lx�&:3@���92�&xD�P��|���lnnzF�,��P ��
��#��������DD�S�q�쒤�t5ɉ^1\��)�i�T��J�E��ǯ���Q)%y�]�hUN�A
3�KcO=���)Q��]-�g�I���X��x%��VLN���|����9iE�W��p�.�\`�1?�k�6f��cʻ�Sx5��S�����rt,��#�\�H8�H�3�(�1B\qmל�Ŝ-�ge2,L�����TJVF0�~!t��g��I"0"!P �?6M~l�Ƨ˲ו���͎��L�晊,]�@�M���|�c�������!+��B���O�v���5�<�^�:�����]^�x�SǑS|
Ki���L�2�<ȋO����fEy�=�¹�j��L��i�ޔMk0?g�F/L{� 64:���0h�(u���3{g������'�4�B1S�FBH��U��T|>bvz�{�!{�����������S6�v<6?�kAFE�{�Ģ��y~V�h����8�0��fy�О�F.��LǊ[�wQ����P���tIc��-<Ó�J�>��QX%.C�Յx(Dx��)�P��3;�#�J�=�"/��0Ff��O
;�O䗼�CĈ�cùY��KQSY�'*�H����p���e &���<yG���9�O�a�gQ^8wF��)]O���C�4NIH"����U�����u��#L�� T׼T\>��G�ϞS~=l^�h�?��=�أ������Ѓ�'7L��VUQ�$�荙&U._b&I�D~vv�.^<o�=���CN��ΟU/u�*P������<�Z		C����g"6Q��+���%�T�C�>h_����/�`/~�{�s����ϟ=�=ZM�T,9� 4��c��T�W�&����2����q]Ο�\Us�=~�Žǉwq��3OZ�	��U���?������{��4�rv��p��0ۓ�t��k�l�;�y�]>�WD�h��#Eј:��)	�Ӣ�G��'���!	�i��S�=·�lzz�N_�wS(��:��L=���īh?�m��fJ��pƸ�l�,{_X��2$�p�SM�9��3W����֪a@�[+�?^ō?������/���{+>e��p>�y�V7��p�d�tN����8� IL (�����(A��@����@h���Yb�^H l�Q�� x��[�������@]����Ր �+�]C>�����_~Q���=�{������:om�
VƁ8MJD��Hi��g��rO�xƌ@�ɓ���g��\���K�=y��/,�IX�˫�@!�̼��Qyy4Q��Fk�ކc�1��N�<i�W~Y����#|��.9�3"�e�[���
p/Z�3���Uڄ�� ��O�J;{�����g�U��ړ�=aO<��=��Ӯ�ܸ�du�T��lW��Gx"�).�x�&m�W}�	�}���R���#�����ͽ�i��MC`�)�������z�W\��J�\���Ž@t�Щ��M{���ts�$m�,az��m{���t*2G��q�.�szD���ڀ�B�Ѝ؜��y��>�l��Y�W����B~"��e��[/U>t�}�{�0�9ۦ)����.[��6W{����`(_�|��'��¤4�=啷��=��K��NK���'\�6��4�¿��G/��c3c���)-�����e<����fD���x�i1xM���.��UA�Q��';��x":WH$2u�L�T^���z/�k��/X�(��\����̡��+U'�����/��/������/}�+���^���~�>������W�������UY`3�4[UH᳁��h>@D��w�9��	�`6��O�s�����/����)�����^��O����_�Ͻ�%��[���b�Ѣ�CY���Ĵ�Ʀ�AG�SQ4�ru�&�fllbRZ£���Kv����S�p�-�z�癧��'��3҂H�J���;Rk��c1+BU7o�VQ�T/7='��E{��611+�(lz=��g�'��q�G�?K��zʓ�)qnhZ��V�\��=��q�6�����Ј�'<��A���!&�A����I�O�<����č睴g�:�:e��e �y�s���:惯��}�D�cF�4?V�r����iEO\�5�I�ϋ{*W&D�S�#g�.�ĶO�U&�`<�x�AS��f@:�ģ8&N����n��ם��k�(�ʈ	�����_�G�5Bz�Vv(�|�К��x��S|^r� ���<ez@��Ct�.��U��"r�a� ���b1i����D��dg��9�]��1�ku�[�Z�G�$��g���m��1o���ŦL��Z�#�W1'���0L���&#v\L�ēO��6K�*ԠQe�8���������K.�`>z����P��fG�J=��h*���p�L��i�4�u���eb~�~�);~����W�q4�31��G{1�8���|	�A���<(Ux�Z���پ���m�6m]�ٙs����!������%���D���#��~!�{`�aB��a���=q<ޑ�#q�B��t��'��,�"s�J�C���W� .�Y<�zϚ�꯬�J@���%����(�=�������j#�4�
�{F����ח��m�˃�/Z?��-I�����\U�ZS��ˏ)o	�%%�E��)�U�yCxq s�D1��$�$l|�%㷨�nx��m�II��K.���b����Qd5�@�Pk(��K+-�3w�����YNEx9.x�z�'҇�	�H�K�ǯx��=�c��t�7�2b���Թ��X��|��<B�_�͞���M������m�w��uL0�|S�� U����
c㓓�ȣ�٩S�mk�s ������]���S~{�pXƼ(x.|J��;�f����	�����5�9fA6�G�"�X�hk�i|�e�M^¾A��ގ�����m��8���B�F�B�T��Q�?x�{��E+��E�R��c�����<�T��279��&����CD��"v��m��2L�>�����4<�p������q��Il��1��^?�>��S�����L���t-��~ܡ�p&U<	3s������ި���+�@y�����eJۭMMۄ��5	���, �$���G�����.H�W^369��Z
2�߫Ҁ��1>5e����Y2~��Hi����g�z]p��d|�:y���&Y��&\���V�<-NA<�w�R(����[��p��`��SH9).��Fe��)ì���j�ԣ���^�<|�[e�W( �D6$�}	/bE��fB"����..S~у��_�jǠ���/��Tﺾ���g�ug�ٕ7==���nK����-�6-��*b����73)���GnZ�3*{i�5�;�˶��ek[�v��U��gV���������2V�*<��]�2�\u8�0o��mGp�[}�ڬ���z�M����س�w�lG)�����T�Y!|�s��,PN	�[\���e�{oY�X�c�n߱�w����[îݺi�{;�5������0�,z!S��t	�'��mM�A��@�~�=^/��zߏg4,<q#�Ӌ�%��?@�R��F��S����X�G��G4�q�f��a|ׅ��ڤ?uF�(��I��ޜ:����Տ�?z�޹�l�X�����ז���+���u���eK���C��Y��FNZ^q���yk�&m{P�ww�[���k����c�������{��+�ڻW�w.��x�^~�-m�X#��P��yp�miN{Ң�v-�R����C���1Zl�q���AC��1��WX�a������F�/t�^-�Fox�V���m��Sk2@D��$p��/Z��x�d�[ ��3�̦b�$b����/� hD�+� �Lh�z�ԓy[
�5K�����;8@�@B��l�w�iXY����#ˣ�3��y��F�d�!h�*s3hO*����c�����t�:����r{��Ψy�
;��:V�'���̴�JHш#�i-A&�R�ʼ!Au�֒��b�[���w�CV}�Q��"��`8&u��)�&�E]���Ɩ���[G�OQ����{���-!�@��b@uT*5�'Oz&����>�.[���(A2!A���.3F���4���t�T}'�7�zK�To(�^vWBFDP�a�Yy��������T�<i���\����d�w��8��ޟ�`S�M �\�)������\y��rmZާ�L�W��o�?g�(g:K�B�}FL�Ytɸ�sO=b_�����|49u-��{W�w���M�N�4�fg�Z��]��i��s������-{烛�[z�e��e{��=[���퍺�������+v�����;>wԦ��˯�f�~p�>�0���M���e�V�9-��������n��lIH8�<�ժe{��'�G�[�4bՉ	����xU<�*N�gL��4�O�����Ǧ�������ޙz7	�ަ���X8聳"}LD��̀��C2��Dx\0��@��PU�;ݺ�r�/ٗ��V�Q����*^�ǈ{]<�x��M�9L�
!Ei��4���s��ں�p�R"uI;ٰ+W>�9�e�b�'Nؙ3�mnnV��@�L��aV�j3���"ȕ��}��5ŀUdt#|��IKs��<8V�)_F�9�.'".�l��E�|O��Qx�^_[��n�ZU�7%�6^�/ۃ���>��S���� ��Eh�ׅ�Q�F��ݽc׮^U��V�/�q����6cu$0 '¾\��Ls�[��1�r���^e���&O+�W`_{\��%��Eo�M�;���_�
���\�C�<E�V��a����6�_�@�X�3E�+�R���sQ��Pg��-qҷ��� <�m[kw�vXt�|�6�7l{��Z"3\��7����޴?��K���߰����[���^�����w���?�u���ް�L뾴�A��K�+�ö�`Aߖ课�a�_Q���v)	��Ҩͪ��T�����6e�7G8F�-�l�Mt��w�eē��wi/���L@�Q�4S�	��M�帖����#̽�G�d� P'�`�*
�pݓ����ى��ҋ�X� �(3��`�<yʅ(����3L�qN�jz/|��U]ה�@�i�f0�dg2c�TW����-��(6����n��Q\��X�HS3"L�ۧ�n�h7'�/..Ⱦ�P�4��P�d�Q5*�'�fOVF@$�Үj�������N �R`�%"L0�|
Q��	�I�p!"ᰥ�WD�;��"�?*��lZS��ށX��D�fǎ-��$���cV �ޛ	_q-��g��}�Hc=��ɮ)-擼�f#ҀG��=�����J��W^�=��h�c��ii[�)1�zc�2���G�@.*�:�	�I၆��V�޵�Aǯ�с޳�G��}�Cǅ���mB�|������&#@����4B��D�|झ���qE�T�\GE��ܳB�m�Wk��H{�Ƭg5i��~�z�]�eJ�yCg��#l��t�C��]���Wh��Y��!�K)9���������E��\����G2I��w~���)HBI����\I>�K>.@R:]XU0��D��[���Ny|��z]j�.'c�D��:��co���4���R�;bj� a1!f��<T�\Tz>|N@8L���#���Y�e���Q�������ޝ;P����oK�ɄX8��er�� P�}�u-%ic�nК$���v��]�L�3��*��و�l6lYD=--gvfFu��r�pԎb��q���`�������o߰%�{���a�V�í	7K��>K[�!Y�P��3.M�&a2*��c{t4�����*�&�S�cje�yi��n}�W�(+|�
!��w��{/�Ds�h1�k,N�A�UqC�i%2k(�m0Ë�ǉ�){�Ĵ4��uGBD�`WL�c��-;�J;hoX��f�-����u��g'F;6�ݱ��]���\gǎ�v�W�E�c������vjaz�=-�dq�b����TG��L����:[��=�߰�ʁ��-��$q�i���z)�tD��8��)xʜ0�ad�N+"�h��'z��N>�'!1���-���m�[����޺n�}���<��%�X��$j1��� ʔ�벤tY �EĒ�Np2ی��|XR�L�7�mz��S^��	$�TZ�K��x�f�Yȡ<�+�@��t%u���=��ò	�v��w}��҅K�:���@�P#��a�b��>�bKw�$$��Ǟv��^h}cۮ]�!!�R#d�HC���v��04����aI����|0���� [��j����۷��g�ٮp���/��ƦUTG
47�fǬ�ڴ͕�Re��3����.
�Ud2�4hK���ꖽ�ƻ���m'8�S�Ҿ"�����Ҙ����yvfR�DEx�٦g_=��Ϩ�&���+j/D�!a{My��/?c�'ev�ڭ;�ֻ�[��I�f$\��e�h��ɆW�>kMD���M�#O�ü>���� s%����<�H�V�K��J���Ui)��q>O��B8Z'���������jyu0�-��ч2�77%p��~��1k�T/���O���5�|�	峦��E-�cs�"�����L'���0_񱽹��TwOf+�C�J�d��F��ůԗ�2�g���ƃ~�&d��aU�D�2��3���{����c[ݕΝ绾�Ҡ�D`��ނt��ة����w�eO_�I@�פe���"0=�`V�8���]�@��j+�B��o^�Έ�V�|^�ɱ^B 	m��1C,eƌ��S�0�[�9J!"Vw!"L�.���a�+�ob�}!5���@E���$�B�@p^1!����T�>��C��6d�޳m5����'��V�U�ٽ�+�s[Z���|�3SS�v�?�L��5d�^�~ӷeWT���Y��v;u��Z���w��;u⤏W`�0+���ڕ �f�n�aT%D���c�&�U��7����)D��p�؂���%[^� �۱�'��'�����0Ɏl��]���]xy����¥��X���cϿ���p���0?훸����ݴ����qln�`��z*L�`D���o����m����sv��_�rS6��o�cִdB�KW�Z��}�ŕ�7Ќ�w����㎼��#�����F��7A/����+����Er	^4m!��h���p�s���������_�����ڸ��R�i���(ᘼ1S|����uDk v�T�A	�0�˂U�,BGZ��s8F�:�c20hQ�+�N�<�|�/3mp_1+[}�[�4�4�X{�Q�lr�}p}��O�����vBD�C�U��o+o��=*!�������ii�y�MB���d`��p^3�)Ha�"
0�w�^?�E_��g7?��s4B�����R�����}� x$�nyH^1(ϳ���0�Hc�k���S���FÞ��%���0��O?�`0�ӺY^~��řW���51��T��"����,
*7ċ��g����MOO���#e�J�$��|�L���y���쫌�5y�a��((�0m��?6q=����"ƕF���i�D�<y����#_fc ���|�b��'��ip�_�u';31�&���I���v�2|���		�)���׏/Зc��/VkVf�mm:�N���p�S�5���5	�	�&��k-�����$T%��s������u�Ǖ���}EWһB/L�Rw���{%�p�99�3u����/�2�	���.�np*�H�:���ʫ%�qKB�β��؆��憭�n�^��(�����Hc�j쉙�
۷]u��$	�/��0��Lnz�n��V��p��ZG���Q�m�a]�M�QWYh%�QD�4%���� P�Aq�vd���س���̝�Uoh1���31d 8c�Z�90�|(�l��P�\�ꞁ1_�+$�����gfA�Q��}��8��+n���
*O�;9��Āa��H������`V*BĴY-�lj����.����y�^��(L]s�ҙ3g2�%��\�	{�����?��p3C���i�,W�'��`��\�P`���	1"34�.�y�g:v�������O����l�c�#Ξ(Ks���L3��W�AD�K;=����C9������ĸ�%{�!�/4�RxdZ�ך��|���`����]puXX\p��A ͊�g�g�ر�>S�/,��`[A�I&Sql�r�Iˏ᧬0>�X��������^^��	�p��'ė�<��U%6�ٛ��'a	��|N�F%�FI�I�ʏxeᵬvͫ��yꍦ��-��3̑W� ��T
c�:�����/����ɷ^��A��KS��I�/�l�7j{���sD�zI�ͨnӺ/J��Y@����U��~Y4π�:��c~o#�GN4���I�3%��]W%*���ĨYs�d{=ю���sk�h����ٕ'm�ٳu�O�/H��W������vOa���+w���{��#a�Р�j[h���N8�O�nǫ<��EӼǹ�)��*-C�X�� A���-l�L�f� ���"~!w���OsD'�$P|@���w��'9ϕ���N�8W�i�G��$�<"v�S��m�ԠY�G�Ęl����؃>����Ǥ�K5�0�.�)�Մ�|YL	�48�H�|��=4��.�q	t��`�9o�>���{��۸��8�ѳdkI�A�E�0���*���4uA�MMMډ��������֕�s��I�"h�)	4"�g���7C�¹�%@^��ٌc��h=y�L����քֶ(�R�y&P���{��sP��(��%�d��jZ����o$\�;�>�*���	~Dy�k�T�/��M�h��	W��g�Ɗ�xc���/�g�J^mD]�o,�B�pOX�B�x��67��_��?�?���v{����b������ڞٺ�7$Vw���Z�nޫ�ͻ{v{�e�-�=	�z�j+m���m��۱�R	n6zvW�ݒ��k��]��x�ѵ��1ܑɱ��r�F% r�7��Ҳnl�k�޲w./{9חv���v����]��ݍ��}y�^~�����{�k���ݷ���?���������ɧ&z}�7��91c	?£Á�#*�O}L*c+Syɀ���ݱ{w�mvM����a�����_�$�=��K�Ϻ|Tg���7�Jc$_=EGL�5C�����H
+�̱�SF��ʊ�r �0@T/�zѺÕ�i�D�o}
�js"�ǀL�m�ӵ��;�h3R���m��u㼎�}ܾ�s?Kb	Dֈ�lnq�{��?����?��b(��®���m��n$P^~�UۖfS�NO�����z��5�[��u[s�g��]�h�VJ�YX8fǏ�ta�����؇�����~NҿdK�V��^���?��^S����i;6�`�*���o/��֊}��?e������@t���E19�<?�ޏ���O,/����Kʸ|c�^~�-�(�{`s�6?#bd`m��r���И�7��oI�:f��=�}��s�J���{`wV7����6w̺�/�����u��GXVO�D�y�v�Yb�$+���;���b^�B�h�۵�,����;�H���O�r�@Y�ue���M�50�!�P���H�y1��r��0��4�^t:'�Kk��=[�ñ0m�x�::7Ig� XW9t�~g�0/�`�2z}Q��+EŃ.NI�i�K{�7�V=/M/�ΊC��6������4穎�&�'���!��iib�nS�ҵ�S�+`n5�nF);�~�;L_�#<��$��@�Kz"�x�f��������[�5�)�ˊU��H�ѓ�����[7o9"[��]��j�W����\<�N� r�F|�>�5 D�����d4�{!M@뿈����y�J�����R $h�q��fkC�F"�^�`e���m�^�"!�d���'S��z�ފݼyGڈz��E�T��0`G��m1�Ϟ�C�n�K�R����%x+�z.���&
�@Q���l�KXp���K[��5Zz-5�����A��"��z�q�6�"B�'�ٱfcׅ�Cv�;ێ�~��Z��-	��O�\��&?�����}�����1��G��v�R]z蒛-��w?��r|V�2�>�����O����{������4����}��	�9��.s-�~�S�{=��1�m��.������q/|_Wj�x f"�u-L���\0PR�S��C��&�jｰ"1�V�����߼iW%�o޼m����߳��8ݹ�b++���nK�����][�}ז�/��7����U�ۮۦ��e�}Cy\�mw�O��+�����]�z�>��]V'D�lu`���n�V׶��R @����:�=[�\�c'���rz����[4]�1}�B��Q���,*��\-o�=q��,Ju4�Ɂ�Q4�?�1&>]��%�!��gOMf�(�:��γ�� ��"�������F�4�)&>�A�����L�|��læ'Hc5A0���&)֋�%�����ʚ�u5	���0V$�+�m6;����� fpĆ,�}��c�#مJ�Ƴ�}sS���fk�+ʯ�������N�|ѻ2��I�9ɑths��tE�&-��1��z֥0 
1oom��q�!5�++�u�������Y�N �Qg$%.�gd���Ξ�{{GĹlW�\��E�s�(���N��i����/��/5��Z,fb<��[���z�EX8p�>�s�aѶ��y�M�o�ȏ�?�w>t�M����ս(�
Ҭ'AXC�0�8\ri썺������	��BG#�z'�w���*��S��ꫭ8!_y�l��vC�G{��/Zi��}�O���%/
ǣe��}�:1�Ξ0<�s��x���T�V%ԇ��m�*�0�B���-(5u�U�Uǧ��-�	�j'T��/>��~𡑅��n���A�1��Ƣq;u�� b�u0����3>B��92�Dc|� Q� G���>������B��Q�]C!E`�����7�&��.���,�w0��涄Iݵ�o!>Ʀ$��z���-I��h8v��w�Z���i̤�j�6%��b2~�#�Œ���g7n^U����U\�G��l�����J�e�U':򩓗�!����T�-_���DUf4!�!aŀ��xM�.�����B�����X[�������� �hrj�g`�_I���/�;���{�w�W}|����UR�XC)��6�"L��t�DbL�j|�S9�3��O�F�*K�*ܗĴE~^B2����Ip�M�!x�������!
.��̒��������{�!A�Ե�2:V.
�qX�8Q�$3�ce1��̾�����%fI��y1��@�'!q���G
U�>α�VF%�U�_�g:�(U�C?�bW8R�T&�Qqӄ�¬��ΰ��B �RG�p*.�1Ï�m���d��	����Y��\�3������3��7���Ko�v�kR�7��W!�����	-f����)A�Ll��qE�س��� bޝ0'��J)��͠�
x%�w�����N�" �ħ�`��25;;eU!�G!�}��p�OS�99��__al���Sol7���U�'ᱭx��T|i�� pЗ̘��x��%����rr��ӧ���lrzRB�MD��aF�פ�^�
{G*��Y��@�c��깿�.k��zmfz���0 �ыmi@��E�2V���)�����gyuK�.�����,����M{��8�u��m�=�أv���U�F/[�YƳ��<�zk�V�J7�2��	�MK�_���1�&���wU˛��H��� ����43^�3W�f��z �c��4�Cǖ�'�(+2�Ȓ#!�q�Y*����#�4%�T^ �te
����������n���#6�B�Χd&~��M��Fx+�S2mm�dJ�j�HZ��� ��T��W���	���P*"8�#�!eE�I8)�4��ħL��QO�4'H)$Ĥ�tZ�0Y����3vb���|��jC����N��TP��Y0r@��;���^�V�.��<��R��~EUE�����xt���S��HE�\|T*�� ޏ  ��+.�o�P*�Ծ∤���R���`+�vCL89o�N=`/�������)E�X��X���ǟ|��'�X�f�iWd����YuR�q���19�uD��~�`1�>�Dd��궭7�V���?lΟ� (ٕ˗��wޱ��vg�n[-˱ӗ��KQ�,R�kS�F�v��Y{��'�/Z�s{M����؄]�@�����E�1�@B����ܑ�z�/՚S�9��@�(�S�����鎝?s�.�;o��@��t��1z#��v�䂝?w��Ai_�v��m�'Do�H����8/_yU��z���ZQ퉏C��\��ږÛ��1�k�W�mDy�1�8-JWޗ�'�8|�}���ꩺI3�����,���ssd���Z1�.c>b��̴'�Y���]>k!F�7��� 4W�U'ZDC�F�:,�B����蘍���2��AK��R�,�j*+4�䝺��V��J)�/�� �w�SqSt�C~<�����#D�����w~�I
���H̪�?�FH1�؇��'��s�q8:,	̜=	���P*��[�TDi�`���Br.��|aq��l$*Z��j�~w�#�?��y���x�q9�o2���Fs�.�T3f�Ĉ��5��#�z'��ǅ��l�Gϩ���E��n�^=�
cv��Y;{S�k��K����)���8����{5&�/��a=g�^�g���߷�^{�^y�U	����ٙ)�	K~�:�PF*G��U���'&PS����Ӂ��E{��9;y|�n^��o�L�	Μ9i�>zI&U�>T��oޖ�3�i|�C/ɢ�XZOUj�E	��|Оx�1�۷7�xݾ��o��/��vw�d�J;9.��>�]��qq6.���omZc[�G���ķvw���8�OD���*�)�a{�WW��y�yO\��7�I�5�[M���*JH���8R ��C�T<c9c�I�t%fm�ؚ�����j�aLP��M�̇V>����N�|��/�#�N��bj'�ɋ!��5������E�3����v?�S�!�X���6�FN���@�w%������7	K�ﺙ��^���,���ͅ��{�w
�������H���4��Y��|��G���������Ot�*�q�6�FGx0��	����#Wdv���`Nu �plF����a�{��1���	��-�u+�H�ĎG��39ӕ��
44�����O��?z��7�I#��Ԣ�Ņ�m�C�+ ��Z�	�ݷxP}�[�.ۗ��8~|Zeˤ���*��9�]��/���*o-1�J�����Sц�z,ڑ��0�?_��٧�Dzf�v�؜$����T�dv�wl��m�j��Tc�zV���B��k5�7�������|�j�+����|�J�+���}lm��d�+�#>����)�b��ﲰ��C���v"t�.�u1��7t�ݎ pzh��t�
g�rN
��3,q������i���`����?w�3���D��>L<�RK�w�NВbx�x��+����/��=f�/0�9�������S#�X%oݧ�e�	���z�1)�����˄H x�{�ƢM��0!��`��z��i������w�>��@������?��.�}K��=�=0�:Q��8���U�8�������ޠg�3��ҹ����i+�e� ���Z�yL�VE�.�06�&�S5���\<g�O,�i	���O���	�t�!J=kX ���G�AuV�RoH���>
�W�����E;{���&�,���̏��}&_�2aǎ���IС�"�P��*������������ߊ�U}�xqq^q�z��s�{�{�1_�O�Ƙ˾��q����Y����{/���7fĆ2����Kp��aX.�^�b^�v��\����y��c,|�*D"�$���6BMBGpB�h$�X��z������X�����>�=ee	l��E��Gsؗѓ��l!~��p��nmLw�e�D1���L*�%����Pː�D�j_ᛍ{ժ�J�b���R���8yHԇ<��CC���]X�q��
t�gT~����s!��� ���|h">��=� ������dGގ��+���?��#|�Sc��8.O�\��NY�?��#�N��SV)K���ʦ۷�JMHa��eQ�[�kvBdq��(���.�A�Y�)��~�oL�a����w��Kw'Ĕk���}�q�q!z���l:d�Б~EP��]��;o�IH������.�09P�ZM�ШML�۔�M�AS�]4�MSY,�g� ��@�{>�X���-͠^�nJ~����1_��/P4v�_p��^_��'��+w�p�@;�!}�J�ߑ����2�0�:�6�3qM>{�/����#�ښ���	%�UN'�h_bM4�4:,�6�	���^�iR�G�`�I�D)U'����.{wx{&�#�s�2�4ș�8υs\��������0K��G�tuŗ�ϋ�9B~0;�
��>�5`�U躢� ��8"�LK�б�$1�5�1�L��O�?��De8�Յ�)I�d�Kg-~�#���_Ӄ.*'��0�ɮd�h!1����r��'�:kB�_��u�]�BVE�1.�[��1aK�<���8�����3'y�Q)��F��/��
`j�F`�	�`���!-�)_V�"�{����X[��U!8z@Y�Z�i�hL�H8z�d}cG�0](�v�ږ91Qo��♀WD�i��
�G��!�B�HC�	Fy�u!��5�Rf��`&��FC=�`�����h,�C+�	1��C��B�|�2c0=zP�,��0�\}�����?z�0���D��ݑĽg�ͮ 8FD��A�T�>��;m+)m !�	c��.W�Ǘ�n�%��^�T�
�t� ������
M�Bt8
�{����ƪ�".��`�2��1ܐaAq�l,dŪ�-3��8�%�{�p(M�A5����BǼ`[�M�@����N��1!*�ጐ�sIu��$,�E��Pc�"=��"�>˩|�1��:��Os		��A~��xHjZR����SV��{�ms{�.Ѻ�0�J��2�[��)�|7V*1��H��PZ�jǎ�sS �v��ga�)���/���/�|3�P�×Y�4�z�R�� ��">���}zY���B-�LbH��� "g�
��	[�ڶvo�*�����hG��p�FQ�g
�L#�?��-�K�Y��,|���
�y���ܩۭ�{��Q2HZ�'x�_e1K��V�E�r/˞�]�!FO�SκGgj1�"�%>���������ÄU��Py�L�Ƭ��D�t1t~��G���k ʁq̼6�[U�).���F��P�ϧy�xH�G��G�#ĝi]�N���!����M��Hț�I�Eh*=߷F��#8\�"O�zA�������Iv��L�XhG�Cg$z�r>u.P��	i�8䙺c�f�Vq�ֈ��AA�`qfR�#i�;���OS�H�2��}�W9�P&O{��?��o
�T�����6��+o�9[��/��[��~�z��v{����h�n��hIx��a���EW�� �Dh���)���.�#�ʛ��u�3w�pi�bέz�ׄ�*�6+���T��pH�B�e4C�7"۾_���M	q���m��D�,�m�Ӱ��N�n�{;vos�Б`ey7k0S��D�/�C9�z�0��iؽ�-�uԚ���~��`��\k�ѱ�5	ح=�(ԕ �U{�#R�h�F�Q�?�9�ϐr�F�F�;���:V��X�H��w��O���<����Ny��Y��^Yt�	lP
����'�4�%ŀ3&:�8�е1ᆥ����Me����Y��$`��0�6S�xС�M�c�c(T m��sAu^�B�a��*R�`OK�͘�yG���S�C����D���7c�x8_CC�<��b��c)�g\��N���O�K�Ld:�j5*4��"T� *�L�T����ǠJ� �2>�����?݁�$8��tYޟ�� Xz7���B]���N�9�5�Nĸ��k}z2N�QvD�[͎�Y�n[�{`�K��_^���1C�'Ӏ������r��mY˱��)�=1��m���۫��{W����|sٮ,������5Uߝ�������ĉ�%B���B#����c�V���ڶ-�4me�m�׷�{Oe���vk�gw�$`F�[���89w� 0=Ӝq$ �Y�VV���ߵ��m[Z�@Z���^��E[����o�۰K+�]���6_ �kl��I	��'���'{u).|�g�Jϼ�׽_=u �b�L�L:�ef� ���%1���
D<��hf�����F"��oð`����)(kC���W�qF�?��}�����^y�j\�X>L\�EG�)]��BҠxC�㐳��'50{�-m�3u]���:\*q�������X�!�9�}�3�Ѳ}t��Z޴A��c�a6�Vi!��IPL�
�ыc8!g���<���i4���8�1CLv�'��������wb�W�H�g�X�����Vot�.�|G�N�o�F$4�1�ڨ�GWn���^���]��z3	��ۦz`��cWsx��Xهc������k���m����v{� #��}�^������yӀ��թ/�Q�B�?+����y� �nْ��ֶ�.���|C��;k��ko��Ɩo�cE+����`�<�F��w%u��?'��흕u�-MdSy߹�f7oߓ_��_{��z�C�����Y��x�����Te}�S'ow��|?�8�Y�P�ǯ�"V�aOOXv�{�P�S4Z3`�B�D�'&��t���2ɟ�\Ä~YK�l�|������Y��;����'}r������ �QB���}��Β{uE�����?s�&{v���cUuu�~9O�3�0d�  "L2H��M���+�߮e[�zW�5�[�d��eY�%ے%KԊ9!�0��{��{���cuu��~�V�{3�@��O{�o���|��ٮ9��\A���橀r�����ZGi��}�=H!9'��j�w�%��@[
8�^�$�TuO���`����K��ʳ3��_�a��/|'6{��3G26�Z��Wi��Ulg��$CKu ��*�z��%��s�㩯��.��:���l(���"��[yN��[މ�F��\_ղ[y�,�fk-n���8v�p,���6�IIP=5L�׾vߜ�/�ˡ�͍�� �fk�A�-GM�Rs�����9Щ������V�[n�5�䜓�2��D��\���j\p�'�I�T��\@dIP*B���m]!�c	z͵��$�pc����o�ʜ�@�:C#�ij��\�en��"�@��?����	�����<��z�r}kg3�j���]Iuz;��j/Χp�#�;������w���T�N�V��_/$Sh�D֫�
����P��t��R�P��m���M��h'�]��s���Ⱥ���e}|�׎�qʆ��`��Ʋ��|E+o�xU�y������:�ك�j��k�鿅��vY�(ϓ*�K��q��X�<ѹl����M4��ޝt;OG��I����5�+���]}`8��x
��ӿt�5#�������G��l�4�+`(i�&Ba���i� U;��~��U�����X��~~�H���U*�O;�$��&���܆0�۰�}EI��'\e�����l<�J#�J��ev��k���LbMmz~)��K�)86�,0f�@�fV �v(�=�ڇL�FND��smc�*	��Se�A���A�/,50]Z1͹sX��Q�`Բ	�)��ۚ�8iü�th|��9L�K�+�D>j"+�ۘ_K�͘Y���#�d���"!�4���~�@f���^��M}���u�:#U'kwo�s�qN�}Ѩ���OG- /f��`��F�fz�����_�ib'a+�w��uD���	J��)Q��C򆊽+@��t�)�!�ӤW��F���[�d>�x���r%�j��}���k��������RW��% e��_:�!��S��cr����y箹$G:a)�Anq��� w���MD���v�����鶰'G!�P�<�P��?VMMdϰ�����YA���8L|��h�E�ti8���6��)Q��f�A7d�D%��8�\_��k��R`�>z���۲=�D�d��u���h���g���v4P�W���!��͝�,A8:�\�R?���n�M}@8�w������7b�Qtn��%.�g��ll�>�[ c��˅o)�|��h�'�L�,H浳@�:?р�ќ@����[�Q��vn��q��)C�U%�hS�lu��ap���<��"�."��*�djn$��f��Z�?}���N5{~��X�5ʝ�ak��"��Ba?ӳ���zњ�^,{Ȑ1�j��Nlԣl�o&�����}ǥ�pt��u}u9V�پ�@V�H>�Mt@��XO�Ѯ��X�ΐq�Oư�ߛ�,c9�k/��Ʋ%˧���־$���h�<��}�#����W�=���6�a����e|Ұ�ZGc+4L�%I%�W�\(/�UJS>Hې�����H��]d���N�*U�G;�7ߙD'��y;dΝ뫎�E�������9�V09c���V R �z���H@!�'5�U(~�p�ɦ�r����Ԝ�z����*���֬>��)9 D�T��)Z������p����Jt%�d�]���{�/U�3��nm {a�=�DY[_�|ZɗUEu:;ZmC�_?m����2��J=G��b��P�%J>Jb�,iZfמp�pѢ�U����Ij��Tr�\ʘu��
'|9�"����;�hSдc"�U��W�uT��Qd;���[�"���l��h](s!{TLF@��s,��o0�X�4(�p�m�{bO��)�:W�FF`�C)TY/`*�؎�����	Y�N,�ڡ8;�L��*8f�;�脒�5m3�d{%�λ�c�.���o�ˣ���%����72��"�2X��@ɨs���2�!ﴟ�ܐJ%�?�km
�:�pg.��u�݉l�����{(� ���"m�#��{����M�E�AU���h���$�9`�wf[J
Fw����ه*����s�:�6y�\�.;9w%} �Q�hD$M2�ib#��P� I=%!Ȣ	�ݜ]�"'����,����t��EC��Jz4�.L�,i���r�e+�hvZ*�!c�@��<ht��n�;��Q�]q˕��+��Q}n0V�~#V�R���U��Q��jt񠹶L��ؤ[H�e�#mNh�Lؼݎ���jnWcs3�.H��c��鹉ZO=,o�"o�I]���v5��枚�̕gF�bIMLs�u#)�Fо.��f2k��jsm�"1�����Hs����0Q;T��蠨h����Z�O�ta[&=��UT@����I���9��m���jv� �Xh�9��r����i#1��$��k'|-��<3O���15�?��ѿf�p��*qH��^��Y?�m��Kp���p'��|�c��^Z�2�'9�ȁ��|`����}�+�C�N
mg����Nl���Z1ȡ�J���5U����ܺ�v�؎<�}�Aa<f���~ $Jm����)����@�ps�&�(���['���JW��qo=����w�b���o��T5�,��l��my�ȋ�yn�i��G>�;�3E"	���*�� ��0�-̳y�`rC�X���X���阚����@h:�Ah� f_���\�| ���v��HL2f���{>+���
��w��ۀ�֫�*1��o^gAA>�y��BB�v��r�J�<H�9ʔ�-<$�+;]�F�Q�8罼L�K��rq�\�C�H_A�X�$z`���vaQR����;���ot��t%p���c����~փL��+���|�}� �L�}������m#/;%�|w���A�1��IY� 4H�#��!Ԏ"��F�w��e��h)��B�Hx��m0���.�%��5w �9�c��+�w^3���`��槥=�\�,G�[u���W��4`jhj
����iV�^Yp
��u]5K?M�n�(��^�S��I�t*�P-�u�0��C���!�і�\�_�?˙�%X�R�r�j��c'�~ۉ�����}Ż��We�'f�I��"t�ٖ��'�kv�;k���2w	S��&\����C���4)]HY��M.{7�!a�1�^n�?�Sk�yW�h�~�ژ�[n^{�w��y,i���"�p�k	xk�}?�޴Ǝ�p�j~i�L��[PBf�[+�����U��c� +]�=]J)��d�N2��_���:��4�ڠ �M2�Nc���y����4��;�X`�?1Q���9{�TK�9�n���f�/-��,��� ��x�� ���a�|xg�
��עG�izJO�t�UJt%��PX�#�r�-k9ᅋ����~�wx�8*˽��!!���|�:�OJ�L%S*^vfl-B�h�f�lU#q��~g(��\j�MB�&�67�^]sǑ�<�̲��i���j�w\�[�ܐמ�s?�χ�Y�G�?��v,�y���-�K�N���f���%�Û2�qYh=�ٿ�R��SM�HdI�o�s�w,S"	�K��&�+A�ia"~�Yp���~W�^(�QR�y���f���ţ굱 �IdJ��<�<ʐk�yW�J�XE%����zh��'�("��������Z�������Fz]�6���Dr�̝��y_MO�u�G'f���(���)Ǉ�����el�9��&!�z��ERR��m�i�g�ǣ�Er�O��j��h��`���`��{�,� ~�$a
��=5��`�UL�	�,j)�հ��2�*#O�M��S�gJ����{��2�Nlg��i˖���wuyޔ��������>�2�\��PT���c^2���.��.`isd	�ru�	\;r���B�h���_s�c6�ׯ��Ym�����m�T���Kd�}�i�I���&L8�����8J$���\��>���"�p�=:�z�Z�Ig���WQ'�F#�<��ܮc�ףk@{�;zɯ���,�<�0R��.O�u��0�x<3��{�媘7�!�M�ټ^��y�z�J:�.�Yo�*S	��Y&d�ڵ��-�����Jl�m�駿�h�ԃ�֛�:�#}L��o����*dQ���Z`T`�啐���NY�~���;x���o�Ϲ�Ēf�����J{�<J,�����W����%H9o,�OOM�Y�iu��3!�#)����\��.e+*���&eE:��E�V��Y��F $���k�]��]�s���[�Ae*m&���㘌�]��#��Hh�p�^��r�2�٫����.:�l�8��o��e�P:vI'��v�Ex��|��G�"=���]�»W��e+O��,sa~��C7^����/��|���7_��Q�;~̲"���<7������7涇ecsqe%Ǘ�������ͳ��/Dm�]K~�]��)��		�Y�"a��W��Jl�N���o;�y�C>��ya$�:��n:<^�p�����2~27Ir�+�3:U�u�Q��������8H7��nw<?��ѱ�LB���!p���^"ls�+(��E�!�~��M'5%Ґ�D߷kJ'��V{���=��j
k.�[�*��%��Y��W��VF�G����1Ix�>ij��meΪ�\�GQ�#��*� �4�l3A�~��U�I��q��b�|���z |Ws3`����p��������J2����]��`ON$�Z_u`��Y�ʶ��"��a2c`b��>�z�'ߔAK02��M���K�~F�1���]3�6y�����a�e���$L���2op0˔i 7�)�||�Pz�h��n�
���=Ӥ.�����e���4�L�}��2��d9K�,Ksq,a�� ��W�m��u��?�ShM���g١'��~�}�&��X�u �^��|��2}�[��s5z��p
�{��!��w�4y��N�焜���t�v
�BD�w8�K'��k�7x�u*�������n��:��x��@��$N���	x���=�� T2oq,�y�DP�~���j��i��w:�$�,�o�Ի�[�!� e��a^>WC�-�9΁�K�e$F��Kƹ��LQfl�������}��UNtF�&���������?Ǘm���:q����������=����+"�������Ƒ�����}%z��S����c��&3~y�����v�>���1!�4l5�+<�(�O'7�j�.�vb�t7�%?R�.�V2	V�,�.��kB���IE����
���_�0���%MY^�"��H����<�8����GF+\8]�6�����I�Uz���˿<�x��V�S�!�s̿NW��f;*�������:���/���d<m�|�PʗI� ���.o��t
�������C�o;�l49��˝�����K��m��4����B�vpT������;);0�z[��6��rr"��E����U��+>�R�$��h��G�d��[�m�K	KY;�Hۄ��*��0����%�W�|�`zbr6 �{�X:q�|�F�;cc�����9V���X���~'Ӡt���奌��a)j��3~� �:[�v�|C)_��x�y�镺�C�ݎW��/�ލW`gLm��N'dZ�����r\��S�*ӹ� �$�B>0C�Ki��i�F�K�
d��W;��)��L�*�k�g>����ғ+��NeK�rf�  ���w�ъ._��Ʉ����wkvJ��O��j������k�,*�w�Mi��#�i��}HpJ��TwE>�޳+�ܕ��L�ȩes��~�)({h&����~~ef�;@M��,KW]o.7bͱByj[�4`҆I�D�8L~��nѮ.£�o�hb�S���K$��$�-��{�0�c��������^��+�òg�f~x�[��},��v��I� ���/ڇ�๰�^ql�������%��/����$E�|�¦Ӿ�u��$9��5^ōċN�=Cw����I��r��|�E������L�}�	WҺ�竃����`T�֦ +/tr�y2 C�|l|,	��t��L:*�Grh����5���4�N����2���)1<vb�}4�1��\5/:�`i�'�PMO��P2_~ޓ�x�FV�1�V��Ue�5��r����s�Z�]�sI@��՜��DěP�Q�W�L�-�;[U&�+#!V`
"g�3?��:b�Aݚe��3�[��,@e�\�	&"#	��Ӕ��u�2�D��p���$��փ�.#yE,p�@��t��<�w�n��U�V�h'�z!anl�[����Ic�9����=v��@�y'��gЂ��Z�oS{��/��~�d�R8Q�;�-�n�	2��]	�,��Q��iy�4�i�^޿�/_�|��k����o|��:��4)C�;!)̤�F����g� ���f�q�����`iKa��������ȷ^���L`���>�Yd^��2�+�_��`&��hH�)��D��,bl%pf�7�n97�)e�*�Y�RV�0�"��*[���(Z���w%�v��çw��>*靕�tK�s�R�H/�8K��ua�T�I�]ԏ���ƴ�ZZ��Ս�&5.�$�J�ڦ���-��r��q���ٖ�8K��O�4��l�N}>��&0*c~�~���g~jL¹��k�|�{��^}m�x%O�|���s&�H���&�]r⑸�
�/x�2��8P��%	uǒ���h�d�Ѽ.��u̼,6�y��!o�<�_�ί�5B�[����뤔���7�7oL�w�݈�� $�#�Jc~"�=.FN3�����x�dW'm�ʽVH��_*?����+����h�_��y�	6���&!����uj��f)�;cu�����\�����k���5?M�(��:Mc�Ż�DwG����3Z�K�j�a+b:�17�bj�Q��^;�|���5�9���B�iG��s[͊�K4�{��P��%4�F#'��rO~�ԅ�v�+�f�2#g�����d$���e��u��,�'aY^��oq�M�J���8�-å�噭h�eP�ߕX�V�g'p����:o�~�YI;3 w������,	�[����>|f]Jم��M�<v��xiA��u���{X�,�IԄU���m���'"]��$Ԃ��K�nY�̻����� e�U�c��o��V~������yzf
�bn�_��}[���H�IK�Z��f�;����)���sVh�`Y`�f�=˖�gj%�h�]�9�{�+��n* X���Q�F��س�����鷶��{�r,�9�?ynC ڶT��H�no�wO,���v�b�w�+K�=u)z��8߈�M�
iR��}{c��5#�ӠI �w�^�⁑<��5bFP����V 2���4:NU�2�u`������ێ��U�܌u�P�.W.�1�sf�Y�n�������Z$!�!�H^d� �ֶS��c���s�\���9��>J�T�����we(]�J�i�<��{�6:�yon�m�1��	��l�)�8�Y�����������H���d�բ>�0���ިM����0v`��U�VS�U{H�AҶ�,/s�w�����&��#eJ��ѫ2�Τ�9/{���7jf=���l�ǎ��>���x��mS��Q��I[�оn"�n������vlp��}������lhCQ?��9}2j��F0S�j����&3>2.��W�]��{0�n�l;�32V���%2hRI���N��+��hҾF�
�v.��{]� �)d�OҦ�{�f��G^��:[�0�|��/��Oh_%Gsߔ���cb���ҙF-���s���y�~'�����K����˞P_h�O�����i�~E�=��X��"�;�I}�N?A#Ԝ(��+�l�E��"z!�g� >rmA� <Hb�6(P�,c2�,A��Q��<E:��3BW��c�����,�̉k� �T�17�������@����t��6��dG0 jhB؛]���m�\00cm����>�����j�*�����[U�#��k���20����v�����s�����Ț8�L@�D���ps�)�Ld�N.z�%܇j1<9�c�0��*R.E086c�&c|��K�����{7��f��B�	C>/�SZC��fF����W�3&s�B���D�{�#��9�<̵H�{�V����Hc��5���ԈXw�2�8R�>�,;�	#�)kD5\@X��1w:����O�N���6!Z�D�I*�
����</!i(?4]��#��O���]����,^y��2/_l�7�q�Y�������u�H����>�~�� ��\�����x��r^��;�U��H8���ڄd����d�.R�Q�υ���=}�}�.q129#��vdV/*gШ��V��C��޵�[K�$�g�k�uT�~F>����nм��@r�W�@�Ŗ�{�T�]��"�p{ֆ�^�<��vmQOg�w��.��ˋ�AR�������yfD�n��J��k��YT�C(�Ӫ M{�J`\�2���ڀk^(�l�Y� �q���GWsǶ�Ѐ4]��'w��UbA\}0�o���1�M���� �=|��l��юֶ���ݵ����P��t���:t����H��w�vnA�-�*�S[�䈅	ͅz �.43�T�Ԭ�G=��вj��2��p��6;���k;iϭ(�j1X��)�F��؃�$���ƃ�M�u�f�mj���Cݫg��|iGU<�SB�&b�4�g3��ޕ7�С�-�u���)ƛ2%����0�k�S"5��L���<�r��k?�JZ�d�w^څ�;�fh��M¹���&q�Mx�T�Xޮ	k�s�%Q�&��O��Q�*�s�E�r�@h��R9&��b#��:��4�x�	mN�R]΍���10��K�SAU";��ls1�T��a �#�������0C�\���ns��q��{*ɩ��[a�]�Fߌ�ڕ��u4��j4�ע�`�o�]ǭ&��8�G^G-�땑`v�aj�����7��L\�		L)�\��ou���h=UL�:̆��5�;��2L�w��8�Ac쏁:�
�D%�=t�AqBh��
�7�k�\�!�@�����+��Qm�|\:�ռ�O�[�1�X��;�Ѧz(�
�A� �9n�hj�9�A,�ӥ-�!s��ȧD!&#�ijJ[�L;�v�6��i���/o� ����C���8�"�S�j��8��ò]�fnkBosq��3��<7�]Ү@2�݊X�bV��~y��.�w�\L��D<vy�'e���:5U��J/��D
�mmvǪ�4ϯDc�U�`Мޏ~~  @߿�u[�pa��R����Σ 1�jW�9��њ�?������Z[%ߎw�j�@`]:!@�N����������u��*����v@���nB�h}��0�%��N��|�������������@~ls��.�m���
&]3� hdwƪ��ʞ$��ƨpo@=�4�����zQ咁�[�2����|l�0��ct�-7�(W��יFte��έF����DC�؈�44/Wq����`󖰬WW���̼`͟<P�lG�iR#�R���e�b���V���R��54�>w)�\�0l5D5�m���,[j��2i�4L�tT���A&���y�k���G	eA��HhA�k��Jz�J�}���Ґ8O(L�ԮN�}��L�$,��Zp�N%�9d�2A �Ca yR��@�V5�k���R_�W��Ү���~�&����i�JԶL-���LLW����B�
�*����P��������TYџ��ڛ��\���2HD끉d׷?�O�igW�� cky9G�����T�dx2�ռqW�&�첅;Uls�S���L�����}�2��#�%Q��Q�JV��l�Dl��}�4��Q��ז1��Q�����?ۢ��@��p/'�Q֞*ڒ��ØuhcHQ.�b�n��@�����KZ�V�c�Q���%nb*7a$��V:����Ҏ�^,�$��uP�5�2�2X5[�qe,AF��QZZ.�̅�]�Ū�1ۖ0]�WWc��v+똾�ז���=�&��߮z�x�G�zX\R�[g.�����5o���-I8$��Yjiĳ<捼��K���?���_#�7m	7{hH����+�H���%λy�ׯ�w�wu(I�`��(�3��>���w":��@�B#�CL�/�.��*j;e����ߍZ����Ѩ�E7v��>�º��7����Ş�^�Y<��Gj��3�H��ڙ�y.l�}�J�Y�H�ͥFl��F?Z�>�̈d< Z���dPr���[N��De	>TͽC�!�-��)X���b9:�� �.�5�H6'�;��n���r��nӪ
c��ĬYY���Sc��'];V8����0;���H�p�E46���6��٪ʻ�mo/p��m����n�;[:�h���`��K$�I��4s;H�#S�꘭R�~�k���d,�;��	�С�`��;F�ƭ��ش-5a�1q��a�K<s�M�6P�
��z��EZ|菉]'�p\r�GR�`��эj�m����<�1�.�A�F&��Wrm����k�s�r���
v�6�E�v��3�<�[��Z1{! � �1MX�IO4D�s��~��oĆ���ڔW�L�h���N/P��|gz<�ɂ{�ǵ!����*s�,���<�j��ݳn���O[+kH[I�I#�صH��C��Noe�)�˶ML}[-��-�"�����bR�C�Պ�AӇ1?�z��5g 0��t�L��CsW�L�z�(�����FP��T�> ��D��1<�qX;�TSȘC�A^J&�R��Q���t4L����X��)�ߒ��)�&o� �3Y\^��'��?��zZ,�rC���I,���N���QD�0������lE�F�cw�摆��<�#��^�܈�\W�
x{`T�B03a��.m��=3�\8�,v��S��B��2�U�P7�8+sJ_��6�g���o���}��T��n�50y[1ԿC�<�Y����ѽ6ýѳ>u��p�924#�vu�b�쇁�u�i�u./E_�şik�z?̴����xhd0�^���#gVcj�v�i.�gG��y+{�(y��j����@9�u�tSz(�N��� �
ߓf��sC���gF�U���=���+L$o�2��r�. ��*�ת��ډKϷ_�w����H�V��~������|��_���$��th5�c��������sD�"Ib�"��颲w77�������빔A:�j�B�t j�	�C���c�ѐ��UdR����e�W��'XV� b��l�Z-͛��F�-,�=�c:6�W ΍t����X�>������"�ע���ٶ�w���6��w ��^���l���n�v@ƽ�ڇ�ML�u7n�}ǡ�e�@[R��w�
�Vu>K|�M2GwGԗ3 �9�<�s�߲�a�e�4T>@��D��<��nk�D�V����h|�h���:��w,J��J�� 6cmq�{h�<s�a��Mv'��i���/�+��㕋�3S��@:��)�$��Fc&3碹x1*�%�bt�L�����i�9�o�`�+��U��(W���Yu/������^���g0c/c��D�o&ճs�E�5b��`�Tca�� .`�
�}~` l�+~m���y2�r�4B��^:1�a$�?{u�ω�2�N�->w�����y]>���,��t :E�aw���llb��tv1��������d\XBJ����j���mM`m�-�]-wKnFcWA~�F4AD3ϙ�ؖ"���Z+�gf8r�΁7D�����	0�f��!L���
�fw�4șj���ȿ��0��}���@��X�āH��[h_���P��\��K!Z-�
uq�A4��5�Cj�@r�PCWׄ��*DjRL�^��uX��P��5�`zHg0���!9�&���=�_�G�Z׹�!��ၯĽ�p��(ec"��7�����sNǝH`�@fm�J����
evk������HM�-2�-M�EX�n�-.[���r�
�2K�?8w-�p���|h�dtS���F�t�}�+�0ǓP�L����#������Vanh��h`���4]��Y����7���u4�߄:�R:��="�R@���v�����0��#ո��cd�#��	O������-M��Nq��L�vq��&Ϟ�	ʁ鹲��d֛h3�!tb���#��g^�'�;��_�Q8�Lڃn`�9�:�D��G��h���Pn"O{��%o�n�9����H>���_��D�C{���~�2��N�96�P�sl�C!(vj�C䷺�� È��f��_�l|�����w���C��`"����z&bt*���|<�̅��C/�o��87�T�:�b����RrEl��e"�k~�D`Vb �h�
�,OϨ��h��x�LsG~�
zy~:F!Ƒ�k_��h]�3Y~�W�� ���:Nn`�//��C�����?��n��F��L����$�� '{Q�2�~��if���D�G��]���F/ҡW�O�? �P�~�톱�������z�ѩjK����DߌcPj�\�U�l'�T&���Y�}�[-{�d}T`G�kMs`a	������_�M�cE�75W� b����"#q�}2!;%���\��f#&*;��dbt4FQ��j��D���q�¹8{�ljz?#�GS��_Z����8p`�:l�ԛ1Ly�j������C���,Bm�6x���gN���N�VƁ�����%C���5�-�c۪v\Kok%�����O~$�9��_�����mai���hLv�h&�֭��W%�̵���3��K���Ot[a�����_�������� ��\�_�#���D�E?p]����LD&�=���1
��`X�W1�Nu��v�~�?9��)��`���>y�(���I��!��D�τ.h��D�tqv:{�||&���|*.#lz �MTT���g"�&Rw^��0��Y4��;|��D^����a㴐~
]�nƻ�~O\w� �6�P�����R&��&�K��1������~7塑 ��eL��?z b,����[ll������n�y	F��S/�C�<C݆i0�j�F�@Nf"�
K��AQv�w9��ei<�[^7��������mw�{���/`[�y��ij8�:{-��J��cc(*h ��h굢�,�/���u�OE���v��rD��.�}&���߈9��=l��U�:lB���k:J���m�u�8�`N���>���\�7��q�m���ރ1><��u+��Kӗ��� d�L.��M� m)s��C#���;8O�)rln�0M�t��c@�����?��/����_����
(�
mʿ�N��jؘ�s��-7_��_��q�'b�1���t�I\�4�+�wc��`Ƙ�L�(Ӱы���:�Sߑ0���Jh�jA��Գ�����<����cd��m��'a�~�X����Dh{}:LD�]g�����[j"K��H�}�}r0⟆�ڎ����������՚��/ݙ�����]�H���ə��מ���ʣ��T�U���k3�]����Dr7-IK �D��]�j"�|���D�@��Dz����x����������~��ı��ر�i�kH3�{G�Df13=k ���9*l��p�&*i�V��!�!r��~��h�ull}�U�(֑���7������J�{�_�46�l��.�m$]Y���o9��	w�n6@�[O�����q�7�u3V��}�i��/�>eڮ�V�>:2��Ҩ��L�Y�Lj!5W6어$0J����"D�eW?v�@<����o��?�ǟ9V(�v�.@`�� ;rw�j/�&����p�RWs'�i���F�3��;�]�)���ݎ�EK�L)�i��_��Q�; �F�F3E��C�U��>���8��d-`H�c �fw���D<����W��ߍ���fw3�;�V�5����kQ*1��p�b����/�O}�1}a�v��Sz;�m0��"fT��y&n[��k�ժ�f,I����N��פy}d�H�$��^*?04��O�e����>@;���f������ёX�]l�h��/��-?���.ik"���Dvd?,��0L�/a�|��C�	�3�]���!$��SJ	7j�G��z��vՁ���_��^8K�l!�«m�\TͶkK�#�pa�I�*����U�$0=2,�/����JfE���%[�Bm�7���Ə�����p��)	�I��:��-X�@��}�W�{���v/ZD����p�XB
.o��|�ĳm$��{��������X[�0�̎1�5��&�ȿRG��@'˞�|S*�.B��ۆ!�{�M�ӟ�8߬���tv��c- k������6��&�`ae#��c-��2�����F�a̯m��J+�V�<��V��69?��w#+`��o+N_�;0�u�e'��SCp.͆�^� �����c��UL�w�����{މfT'�m�sm�Ab%��i�뱄���E�6��7�ƴ�)�Xݠ�'��@PL�/S�M����~�{[��e��;����_���b��$vqF��PF�zKj��U�wSL�lG�wO���B�Գ�Z�|�3���	�秢E���g���L#�;u1�|�l�|q>�;=���d<��K��ǟ����7���~<���>=�|���@����t����ȣOB��Y>K��q��+;4��J?A_�do�_��W�)M^*c�^j��+���j�4l�A%�
�Ԣ�R��ߓ��;����;������M(Z��&�`mo*#�?�p��j4�f�2x(�M�W��߈�T�%���Y�&"�[�,H���^�>47Ur/S��J�ݨJ7pu$V�����!,���qv��s��Pj.�EZ��������ßG:6Pw�����l��1��?1>�Z��myc��A�j3�,H	K^���^�#���qme9�V�ht���uGƭם��1T��j|��ߊ��������x�T9 �o�I	2J���������!���sm)>�������R�.,�7�z�L<�ܩ���b�` ��e;�3�1��v	���`-�ܓ��4�can�� @��c4�b��P�v���k��h-f��o��ߎ�=�t��ǳ�V߂ݦ�+@�n?iy\)���0l���&̯�Պ_���Ǐ�筱�r	�b�D=��Kq��b��K757�/_L8Ȭs [�W`h���HZ��.�E��;RS��:�{29��{�[���goԅS�/��/��h"���
���i@��G��/�p<Ϟ�z���>��FX�Ujqyz1~㏾�|�)	���pX�]ƎX݀)S��l���)�Z���T,/-d��h���?j��?�����#�Q����M����?�����FK$�P����̊xF�:BZ*�
��v��(��N���<�:� #����&~7L=�I�}r��i9$NJop�Zu�F���Ł�F����?��;ӱj�d	��
��R�d �H�z��+�sQ:�'���_��[H_TTx	�
YJ���y��)�W��3ij�G�� X'S�A�d"��`�H�V)�#��rO5����)�����}�6��_|�R������;O�'/�G��U%p��uN��Q�J���l���{��W1w�2iP�h�ı����x|��[c�x-��_�����L �H�0H)���ZXi1���D��.�>�+��3��@�W���γi���������?�sH�m$qk��I���X���ZK��ױ�����^�-����zbe}3����>��g?�����X��D~�o���ⷾ�HF#}8_�� �^4�~ګm�*؁H��ȿ	Bm�/|�C�o��X�z�?.έ�?�_+������:Eƒ��h��M�d�0Dh����Cé�oB|}1?���-lpOO�q���ٟ�h|����0������W���+��F۔��wB<{����bo��ʱ07����������d�㞛��J,����~=���|>Nϭ�&�ol��`
��@�8�u
��0Us�QG��O_>�3�q[�V�Gm�~h�M��˟���}}Lb����?�����EN���|�D"��iI_0l8��))��0����#h8��myf.}_2�.%S(w�D����-�HL#j�L�Y2�=0AHllV)�Pk��}�]�ޚ'�ڄa�(�NP]j�UD�M�{p�4Y�(��R�x��1$ёn����k��{Mt̄&��XA^&���Q[q�ܙ���~���=_���r҆�����@�>�'񹧈�d�ш����/3pQ�H���1K��z&��Aq ��(˕h�!�Rn���J��F��$`���58����@��C# 	�Ӌ�:T1����TQ]sB��ǀ�*` j �����/ģ�&�:ve�^���{��abl$w�_��A�҈FWC��,��!�	�C",ҼxG��=Th9���@?M���=�1�=���y�}[��k0g���#1Z�Q�bc��#F�~�4�p�!'�雪�E�8T�DdoA��k��[e���@��������3��� 27���b���u�;*�i��_5��r�o�`�*u����U�� 
1G��J�N8����(R����t���t�@>M��g�-W�s�Ûr	ڑ�u����Ȅ;{��P!�Td�I��WjQ��~����D�M���Oe��u��H�[u�d�9�۾��&0�AL;� �N#w5�#��xe�Ch+� *i5�����Ǝ������q��Q�Cx��Y�v�)��ûe�jQ�f��F����� �|��􃄇M@D���%p5�)[���7�!�����z��=Y[L�����:�|�����\]��:
���Q�ˎm��#e�E�I&�f$j~�ܶw����R��h�:�����7���F��a`<1�&C���+ѳ���\ݫч9׷�=Į���{y��vv�NU`�l��U:C���	�2����9�������A`��y����H�����G��e!��~�[��o/� qp�rs.�{�}[�{}|[D�h{uA�	����ܾT�����a48�25�$�R@��������!�^9�������J���{ޚ�N�7e"J�$��dVRǋZ��Y�va�
|@����ݽ�����1���T��έ�!��o��-���9�Qtm"�X�k1�q��MDA�@\׌��`��p'x^�i�
�Ç�HP9�\� H����ԯ���H����?08��(M������W�-�Œ�.�ԯ�н#���[��8����jLֺbr�{C}1��`�"V��D��L��`��5̀�H�o��1׆��D2�#��8�=����d�0#W�__�^�U}G����F�V�{�k-*�ʺGƺ���j��܉=�����Ğj\�o n=q �M���vBx�};h5h� G�ZB�����CX��
�	k�%�� *|m��=.�Ȗ�]���h��"��t�{�zk��qˡZܰ�'n$�ql �:1w��;�7�~��h�5�2��4
���t�+�;��uh��=��.���D���B��;�L?����e5��:�A��2.!D���2���c� ]wj�/��p!�.�m�E��:@TB^��?�df��}|�7{��F,�'��*m����*=_�����a=��@�qt4��[���쉷^�7�~����D��VbK�y��.�NBպ� �zV�V@�	��Qa$j�s��G����0Qu� � ։���v��þ��E:s�2t�k�p!���N�pp4��p�{ӑx����vK<x׵o���Ȼ�'�����n���H�z��k!��~ F�h���Av����f�ہXd��v��g�/�	n�d�ɸ���D�ZwJf��:�^�0��e��P�������-��`�~|�2��������|���w����񱏾=~�������~���vӎ��*��c���#��91����� B��'YG�Q]҂1�P�o�W�T�	�
�~�̻�)>���ǃ��������?��ƿ��O�_������g?����{cb�M�;���B�j��А�4��������b�`�<俼��됩�~�<v���Q�,�����Ua���)�a�����3z�ӖD(�!�el�d2%
��B���t"��~O#�]����on qi	��D���&b{v��@�f�?��@>t�M��{n��3?�@��g>?����G�~g���[s܃�Q���e�8h���FWz�Z�_H����/�!R�:ZG�6�{.���l�\C"9t{��x��L4�0A��ͮXh�����xϽ�Ǉ�qW���[ۊZk> ���;��r,>���!���zD�8��D��&�qlRݵ.��-�y�@Z0@�X6��s���9%�.��:��v��hTή�k��%US�Ǣ>6�hHk��ǎ~����G��=�͘�n`ެc"�ǁ=}q��'�C�;��hl�;c����?pO�}�5��4�bԁ��\�EL�U���Q t�lS���f��s��2���0�׭-ʻ<��������Բn��h����|��ƣq���k�Ǒ}���:ch���y��}�Ô��T �D�f�*X,M<�!��z)�n�Ӑڛ���<�K'�/��4��]	 Y�o���X!-#�\&�Vb&&轴���wT�,^I�y)�!�m3T���ﮊ�h�a���'�p���Tg��%�m���R��D";�ls-F��q�����`,�\���g�+�b0�z�q�-׃G!��s�q�q�=o�c�E����B+��Z�õf5g�q�hNe��J!���X�
�c5\��nR�T�5�WWP	!j��N�_EU_Z[���I��8zp/�`�of��O���VL�;����?>4�ϧ��o�;���wƻ�"~�tÉh,�Q>@���
a*r8HJ)�F�9�{�;cWX�l2�I�r���sM�5ʺѴۿ�[�	.�6cpp,��6���q�ͷ(��G�/~����c�����nO�|�������x���⎷����O�/����O�ԏ��������e���$�)�L��C���[�Xp�Z��}�Ws�0�԰WB�u���S�w����~������Q�}Go���!d�H4�+ȵZL�?ա�8p�p\w��c���xǻ�'��q#j�B|��H�ߎ��r������o�ݤ��v�Ѕ�[V5��iv�
�L3�]��y���3�ߌ�Ң���E�V_ �����7e""�����=&T�GP�%�����:�,����˂�-b>�_dy�Ĭ|�؉������	����&1HN�ִٻw2~�ӟ���=�ߊ�{*Μ9��zS<���c�M5�݌��x4ξ�R\�����?��''FAt���.�(�ƴ�E̬3�Sw�ʺ�d�N�@�VG�� ��@��V��U��!��^pn`��~���u�"Lg����n|t(�x����kq�����������0w����ܿ�����1��V�E�y�,�gjT�d.�ᚠ-�7ص����S�E,n�=s.N�|&M���:��N����A;P�����<�����S�[a"��o|=._��ϝ�3g_�\7����q��{��x���As�8����(P��E�v�wC��G�w�kЩ��v���Sqiz:���م�XZiD���V��Ǿ_�����_�j|��ߋ��1���A��p�󷴼
������s��2�	��Z�ɀ�:p���yc�<���C+�$��y�.4�&}���7��o
�����tj���M�C2�m�{�>7)���G�o(��1��AM�RU�q|B��:��A��2]y��c����0��@k���Q����XkhK+H�\���/�Vblt�z0�F&@�s�̩�1��`�z�}10��QJ�70_�Ʒ�_���O��o�f\�#I�ߗ��\���HP�]�H�<!LL"����Ȫ&D��~�U3r�NIJ
!�HS-
&���~}9����r�E�r����%�����Q�]��ݳ?�����>��� �����[�ֻ�E
�Ţ3a�{&�Giy� ]-��e�x&Sp{�Y桪j�x2�v�jVZ�RJ�-�����O�9/�9S��I`�+ܻ�ˎ'����S��<D��w���r���1><7�8��x9~��~;>��/ř��pX���ŷ�ͭ�Ю{�V[��6�,1���V!�'ĥ!�x�Hd�j��_I=Ϟ{�9ɋ1:6��zd8�Ԋ��`O�>�K182_�ڗ�[��z<��y��'�҅�3��t�������o~3�����4Lҥ2�v��qst�&�5mr�4B�A��zAw�ݡ�l��
W?�,5wۚ��xu,�g��gD�e���DR�{�\��LĬ,�]Pn�蹶��_y�@f�3��������]U����B���tp���A=�$�Ql�xչ
!5�T���7�h�&i���/͢��x��+�,���4455;�>�<����r���`���0�D�s�_.d,R���D1X~�(�:��LgW;R�\Sts�s��2���'��l�9$���F�`�\��1 ��`�/R��y����<�f���C]����qin!��/.-��q�S�݄ʉd��@bj����ә��t�܅��2gk����5>�⮢���_R�T��瞋�/̣�vL����ǿ�H��o��x��簵��Q���r<y��������O�i|���ƴ�,�L.���!]��ú���4m�v(x���r��F�%�D�Ŝ�h�b]���z;evL��a����<\5�?G��E�,�������r<�������̅s9�v��hLc���C_ٿ?F��A]	�n���'#w@�E�WNv�_Q�vx��|����S�%�|¹��s�
�<����;�sQiB+�����L�`�����n�C�޼Q�:u*�����y�%�_U���2`Q��4R�w@��Dq�Vzڝ���c���/�D#հm��
���O=/�=g/^��/��c��;�1���K���}7Ο?�C�G�A",Zz ���+�,�)�g�����q�̲�9PJ�7ңQ�R���p���?��X^Ng�Bc����8p�H�ADg؞�p1+k��H��%��b2��f+GǓi�t�T\D��ܻ�=�XS�������\>@��?�yWX��Wb��c��Z�wˠ�>������}�������v���_�r|�;ߊ��kХ��?���q���.��;6��xS;x$�����C�?�L:�&x�<]��I���dR.�$c��7m\��ո��c	b��(��2I��V�����G�	��5����>1��z��DL���p�ޯ�3�U�Hu|�����؉��%��:68�C�9 ��˥��@K�^j�~���w�_]�W�T���.���}�(3$L��H>&�>ϟ�ʿ|�y
C���W���2ұ�tH��j�j�D�F!+ڮl�Җ�S�݂����x�`���,Y�y���ݨzߔ�N3_gI����K/��4p��M�z��/�1�:=q��8�J})�����%L�����k�sm�2��t�Mq Ǌ�]�_����ھM��K�cOO�M��WÚ�J	�랷U���M�p�X�`pO~��dh�eNP�1�d�Z�rc15C����qʠy7=;O?�,�Ẏ�	a����kngP����P��巼�'RB���7h�d�h��LD�_XL�8h~a>���ϟ��?�d����_Ư��_��|6\2�뮏���-q�-��U�ѱ�t��O��}���p�])�&��c SH�nW?�Z���`�KcfH�*'y�=�̕c��ٕ��<6:�����h=����o����8X�A���r2p��0FG&c�Ygrw���=0�E��K�G�2�鬏�c��J��@��@�_��T�s^h�DC�w~��g�(��j���㔐`i�=�n���eΞ�w�u�����2���LĄ�µ��-@(���W��)h��NWW���:]��@ݮ:bw�[;l�)�R�v�=i�W���ي��)e��/�V�t<n'�����N��`�{&��k���{�PGR�C�Nv����Q8�&�v���i�*�����a}��J�~�䯍Fmp2
b��N���D��؀��-ì��bnf:�x�x�߉驋Q����w^���R�@��O�����O}�)�����s���31�'F!�As����1��O(�J#;!�@���M�m�dSs1�#&Q�s���n�NVۦ��Ӌ�<�'����c��$�ԓ�i1K�j9O�f�����Lu���iԇ�Ehi]�-)�t�u49�?m�7�)מw���y�9'����,������׉h-�r8�9T�����=~�e��e�ce�bdd?��x2���y�s,�85��f���2͏ ����4��R�J�N�|W�1�g�q�n���L�����!��LD͓�Ձ����u���~�W=�0<R�l����d��LD��f�s{4[��|pTc��i8+�[�R�,Lff�;
!q�մAQ(x�G:d��� �G�]]ƄH�'�k�a�p���_r�d���*�ڥ�إ11�}ۛј�A�l�R������x<&&�B��������sP��c��������`�pYO�f�;���0��gO�e
���R's	[P=ܙ_�_o�,+�VV&�	�H|��!��=1+|�[]k�X�A.Q�V�,��̥��)Ηa.̀�C}\�ȕ�V� �
HO���j4��b�oVW1� �*�PS�I`K��⺤d��iX��l�p�D'8J�2`Ȅ�yV�l�vTI֩���L2�G��[�����(�V��E#q��Ǩ_O��<�yy:N��������Hll��R�l8�|�������X����V��x�^�Z��-�PL�,�.����-\��ی��om�/uR�pu���c�^̅�VhW�d�h�=�����j�5fr���s�<x(n����E��3{�c|b$'"n��vk�����I�e�6��^i�bo`�.�x�HZ��Xv�mit2R^� x���}�+�B�؋��WD�m�g,�%Zi��W���K&C

�dV�N|�O[	+�y�$i�@�6��v�AF>���,��'�7�
\�y����}^Ba6���dC�[T@wr. ci#�O� D�Y�$cz�����:$�Ac�c�֐l �d��m?v]����耝���K��bzn>�`*�N\B*]��i�PU�q-f��0�ֳ�����3��o�h2��ͣ�u�ڕ+�.���j���ٿC#"p�w	�-��)���6��Q���Xu�jgĪ1��Cҙ8D���[�� L�Gc���Tk�G��^�9f�צɷ-���Fa��I�2I�
MF�Vj-7�0n������R���ح����ypU�e 1I4�V����\\�<�.^�3�Ϣ,@��*h|��k�����[hXh��h�IGq�1Al�o�{&&N�7��?�3�_+<Zaf�� ڐ�[���K0_�д݇�%qK8t!LF&Fc����t,�tɮ��!�ɾ8|�@<�/��^�ػ��}�r(�z�� �a�b�+�9e���	vJ'�.�Ԑhp"mCl�M�w�<�(���XT ��0���"��*W/cS �Rk�|�N��P?XǱ��.��j�8P�LfS��5:�Te�`#{�X*R*C�x�Z'��uű�=�ѳ�5��� �R~���q������]�A�=�~�=4�$ ���|v*��\���3Ѹ��Ӎh�.G�do�-����a"��ٳ�#�u/]�E��8�vD�
d�� 94�A��A\���[��9-�c#�Vü�T�Tql��.,-��sg����0��\�xqy)+˱��@&51�m70mK������y���l�=ØA�����D�`-M���r���q�[Aެ�n�E�1�̛�Zi�@d\�z-��&3�ĝ��<��
�b]WC�AS�!Pgȥ-���g^|&v�+1
���݌U��v�7QG@G�  b�ͳ��-5֩��g�(\)�U��[:����8(�Nά��F�/4�t�~���������q���E�\<!�xD��O�/<��ܙԾ391{���e,]xktd4�?�R���fD�g2/Je��^+�&�zu�:W�׉�zv�k�W��xH�K��h;��������<�7�7e"n���c���6�ғ�Ȅ�T�BX�ׂK�2WǬQ�\6I�[�Jvg΁��Ű�rbb�������p[�#�ǵ�_�c'��,,,ƹs����-���?FjH	W8X��m�q`o?y���atlm�/�����\��^�+u�$a�n$ʣ���~}�bj�6vZ�&��Q����������t����:�LF��5�;|��EpǮ(O �ug���2	���^6h3�/�G+Fk0'{� .�9Z�AN4��.�
C�B����v�n�Ɏup����1���4�(dhp0n���8~�H�|�q�m����7^{"�?~4��{F���]�N.�|���x�m7�GFUs
�2�:ه�
�E�_	9�r���WK�,�mR�͹���+�Ǆ>\��DB{>|4n��ָ��9?�0�#XZ^��_ ��˧O���z:��8��cq�ͷ�w�%:�>;iG�'�kِ5R]���2�������2HM޶�mC�S����ko�{�k�_B�#$�YS^��v �N�l�`"jm_˛2=��{�d���6^Μ�S�+��"o�o�R��'7�����  ��IDAT�nǉ8���\Pّ�c�����V��$��S��#O<ϟz>��3�g�ػwo�q����w�3���x����w��#E����c7�R�U�l}�E�蒡��i����Gy�Į�կC�s�D��	Ɔ�1a�on�c	"��W�սV(��SF5~���o������k���;9�k�Btu��P�{�q��������������o���`rh@�5�v�I�Bk���`ѧã�+��H֣�%ۉ_�2��8q����Vw.��cU���CG��w�+��-q뭷���ߘ�w/���d����0��A��z��w�w�vK��N��W��E`����$�
L߉�?T�
G� �Qps�~����L�`Л���!����0�"�맸BX�>U����X�����{P�*�-����V��btb_>k��N�w����]�2+5�]�S�u�Ճ�:m������_uj۵��4Wb>��g�f�㺭��th�D�xS;:k�ޔ�ȁ�?��Cʩ�Ӂf2�6d%@��Q�U�<^�1YS��J|'���ꮆ]�86cf�+��H����� #@ܿ���s\�fza!���b�����b����u$���n�o�=����8q�5�N��FXŌ�pqJ���)��a�1�_)����js*�mj�?ag�#�k�
u�������uO���S
"�n��ػ�`�Pn��0��(K��c_�s��Ѹ�wǽ��[�G��f5}��G��˨�bal�x�;��t��_�	���ړ�̻	.cR[�F�<�M [�ɑ���W���ht�0	��e�Ļ���D��p�;t ���w�F����h���>3�V�4-����&�<�=�
�0q.{!Hye#�M��uid���y%|�u�<W�߄�ݏ�fҍf���Czhׅ��
·溭.�=�?����,���tV+L��:��%J(�4��{�Jm:��v]�q�����0�	/�Ǽg�>$�O=J�9Әsi�������k�Io�D�@�c7�vlaU��iB�s@Vm�jO�b�"?T<�(pDd��F���������pB��]G��&D3?�2tE��d�'�և��F����"� 0�V5TsS�Rcvs�L]b~~)ܒ���ŗ�����(ru����O�a#��i��p�~�7tع6�3�����B.V��9hlGg%ұ�E�A�W?��6�7���ݧ���D�()��Ȩ	�on#	k14:FQJ�9~D��i�-6�?��Yb;�7�I����2P=�0���dᲄ9��X�K39 ��R*��73�*�A�L-nę�Kqvf%.-m��&L�o8Z0��VwL-��3/���_|9�����qZB7�#:ua:���s��sS�Շ����دY�W���sn���5�t�v<��g���Z|�{����"�;�ǭ67���_�'�|2�}�x����Ξ�'�~>{��8sq:��D��3q��{�0��t�ƽ`�]���ޣ���F<��3����^yﴱ�P����I/\�z��fO'������c��x[����&�|�z��|"�w�F%���j����G�
��Ć���tz:W�nl�pZ��
�x�-��R�Y�L� �z�% %qf�n�ܧ��T�v�����Y�,6<��s�x�Y� �Lg+ư�����r3��xa&�������ҩ�T��Kh$�����٘�k�"H?;��K�J�1fA�eT��E$HO��v���;x(^8y.���7���h�v.N����0^4%��k��ꮀ�dJ'�:�h�{�t���B������F3	o2%9�8�$Z��<�aqy&��O��ꇈ��}���s/�ډ{����Y�|U|,.N�Ƿz,�f�Ѯ�����-]ڍP�wa��I�䶗�%��P�N8��ܹ�13;CZ}9�n赕F\�|)�}�x�Q�ߏ� ��^x>N�<��.�K'O�w���x��g⡇��^:�Lȁ[�/;8<��,L��O���C�?I�9,�nJ�JX^�!��a!(��V2~��{�띭�����^|).^,; �)�F������s�攈�.N��R<���'s,��S'��3�Oŋ����ŋ����K٫6��3>����>�R<��������\�vՏ�f��'�Tj|³�mWhM��e��vlj"��D()�m���'y/'Ҟ�@�4U�n)�$�8��NaPPlڋ	��T�sك��eo�3~�H�I� ��'�ɔ��(/pc��=���۟$��?��8���n�\�C�	i52u�a�w�	�i��� �[F�Bͨ��f"��7�Js�<Ɔcmv�l��*Ք%�H�=���^a*��18����-h=���/�E�f�4���ٓ ��#[�Y��5H�֛]�z���"�J���B�Cq����>�k�������q��k���t<���@0P �N19���ۼd�Q�������xI��6����lɱ[q�����c1}�<�Su�����z��bm®I�u��Ȣ���@�"��q�F1��s�'g��z��r�߈���8p�:����1���f.6,l��'�����"���fg�j��?it�.|��r0����(0�E�`Ti���V&:��0#�P�o�-<
T0���w}2^>9VȻ�j��N%p܎�puL&H���
��\������*�j�A�'|�G�q� ���kntN-�N�qqN=
��{�}ۡ�T��G:�v-y�<������ؿ_<��s�݇O߉�c*��N�*]��R��@�v�רo�8Z�L�4��Y��A�ACC��˻�0�-1cC����<rl�;&3!�̐ۼ#-8�ə֎F^QS�5�/��g�^��Y:��&���2$�x���VZ�m���s/��j�ʓ1��I�,���g�e �Ә"����L ���S����'ْ�@��� G^�I��S�<ʙ�z��^)a�Dcy1�ٹ �&&�X��$��0�ϝI�aan6\�O]�U�ak�u=beq&V��(�:������s�{' ^~rd<=��z�œq��fMo�b�o���29��P�o9-;�_��j���L���cy���⸉��.��l�Y�������j�ų/ǋO?��:Νz1N>�T��̓I�>;��I�OƋ�>/=�l��D|���C�I�_w=<�Y$��2&��j�G��A�qC.�*��#tO��9r$�%.��,��f��6۳������>���.�٩ L˵�p[��X`�Ta#����y�Y�:�F�c"���ݰ¦#?��h��:!S@Il�0��Qm����n�Y9���5����v �[|T`��h�2��m��m8*X&����P�/��*��w��CYaHۛj��<�c+Ɔu�ׁ�V���`���Y���ڤB(���+ĳxE[(��6�AX�K	v�2�[���>MB[�����R@L�,�ᷦA�\��.�%3���	�&���l�3j"������W��}̆ Q9���iϏ�B��t>0X�R�7~�����h^CYy���͞����)Qˡ}�+�)AA�e�x	�^xhd��Is۹"����{�$���@5�z@n-t�w�E�x0S�F-T�i�A��؁���,�hV�'Ȏ͏jC�0�WT8kS�4�g��6�����,�3o�4}���!cJ'�7����ѳEr1f�c})�V�s�DOk5�V��0�m�+�H��K�����l2Og�*�]xG	���4�r+F�.��b������D4����v���b���z�Ur�v�bù� ��lv���ݨ�v+�<ZM4<7lB[���$��ڣ����5G���dꎟ���HCa �r�p#����E��7�v�uy���ϿnvB�P9�:w��o�ٮ K��/4l�Ǟ7q��l���d��=��G>���G��p��g?����3~��k��z\��h��@jGЍ��Vcq��F/,�E��˱��۴Ph���K��s�n����B����ۉ�Fƫ��w�	�Ax�&�>vN��W�U�z���ܥ���#O�,Ě�� 梉8*C�r��&a!^O�e �����)��s��5�L��]z�N��N*G�H�'_WR�>L�N�e��r�;)�����:���J:Z�G�
uxdx FGr�����@��H��M��bdp�}%������uѭ��z�S*'OV#�8r�B���::<�������uFk�%�P~%�S��L�Kwo,�n�J_��k`V���+�����7\7`�p݉8z�Poo!1m'"�[�'�a�������WZ�Sa��TM`n����NOOs��̻Qs��Q�!j��Y�6���95<T�MW��i7��_����+�����o���uG��}qם������w/����O�m�荡�Q�d�h�Z}$.aB� )�+��@�jaf�\{�^���J|�k��PNS�����v�8��z#6��.-Σq-���H����8x�@N;~�X�s�=�гH����Ğ={��'��9�?r���\ѿ�RE��fc͞��Um-��� 5�HSC��>G���(>�}�T�Z��a�m!Y��O��ҫt�N����ү�w
e�)�A�;�L�:�N�+�R:��By������'��\��?V��Q�d:%�O���:�OMȱ	�s�Z���h �är�5��J��;<���#���B|�S����'��~����/��9���?���g㞷ܧF�˨�-�"1���Dvw��v���aQ6�zu�F�gS��Myr:�\oӑ�[͵�gkR��,�tO]��z$�5�>6�������/�2oy�}��D<�����o�����S���/���$���)L���'�h�H1�LU�y �Jwal�����0C�P:����i���]��^��!�Vq܅�)����D��w�+�<K�Mn����}楗�������7�LN����9���asw����L�T�Iә�J�D�6�$S�%z;�By��o�?^#�����uZ[_#:�r��<F��G���?��|���%L��~�;���o�s�g���186�[�V` ����Ss�Bn�n��ؚR/�q(W��w��e�OA#(t��-%�C��
��}^`Sh�N^:N��t��k��u���vG���Ȣ�+���u�������x��a�o�����	%?כ����,HGi��������]h�ќM���뮋;�z[�/nĳϝ��� �8sf*�}�T�x�q���Bx���CdC����Ǥq"��I�5�W�O������rԁ�M�D�UW���{��\���o�������Lh���vs7Ҹi��'���oē/��Yw�p�r��W�/^�� o�(�H�L�-4;%�څ���Ǚ�:�el�5M:�tA�R	��^��l�K���皋2G;#VG�zf��?���Ws�ѝ����}'~�x��L|뱧㷿���w��pԡ�cC@M7s����R��o��-TJ�!,%���M�/�CH�H�K,�.�d�
$�0�u��d�kׯpp�s������ů}3�����������/p�D<�����O������C����Vv����cmAН=~j�2?l���$��LاV�唰��u�F@��3��^]�+���=��?&�>֩�Ta"�g�M��oҜ�$���WrJC^y���{��B<��1�p��A@��C �H���Ms�oJ26�ۥ�AH�
�|Ɯ-�=ޭWݚ��؝V��Syb�8�نDH:n�6�l׻_�Pv0\��]���ގc��@Ľ�G�G����8y�t<��#��⍏�ũ��⩓�nmd8�����ºI����B�����Y��j���>�RpkM��2���^�zd������R7g7�&Þ=�h*[ј���hd��zc)�~�x��g�We:�����C'췐�^>7�+��#���K˘n�w+�f�@h�G�m�M
��_�6������m؋p�uX[�ba��)rҟD3V.��~���uSx{>\>����s�^�43�Ҝy����p>f��؈�/�Fkn�9:1�qCoj��x�2�F�`�����jW	!�M Z>}b����y�x�f6���_"�94�^G��Lr�74�L��v���ŵ���|��j�;4E[��1u�cf6�C:N�S�= >�U� ֟g�k��%�	e�,����D=��N�W�#/�4P� l!�*0H�2�-�/�&�����B;����B���e��Ro�3�A ���}W�p|�h�h�~�K"��Y�2C�(Q{yb;wq!^<}){�d,�8���T#E5�]&P
����d �qA���y]��wErH)��0�1��]G�i'&�|F� ���@����3��CQ���F�X]�*�z���S����s�V����_���%�؊险�
���ﱅJ��t	ڌ�j�[�b.HCE[�+���J�-/�m��6Z�i��l,�Nv���|/3�q��166�.����XY\����X�̰�l�w�5x�ҥ\��)�s��`<�DƬ��C��鲽�M�{b&2�0�n��m���׍,c�m3렆(�R�R�</2�|��j
����a���5����	�P�T���-1¬�$�0aF��36}���^X���ze�hQ�W�Eu�Q������C(.Ǡù�����8V
.
�f�L�5��c^�^�����ċ@��h�Nd;����ތ�řd"2�{nk��m�[n�9n��Ƹ-�����Gcbd�x#.�e���#1f7=Z�s/�d._����5%�ೣ��Z�T�R.��L{j�9�.ya�w��v�[�Y��\��	�&́�x�(��s�5۔ۦ!�Ɉ�y�<���
r��!L|���{)�a�h���e��[�J���2O&��X��p�+Q���VQ�xIn�p�"%ȁI1�Z�n]�pk�y�֟ ����?�	�Tzc�:l �v�]���?�q�=��[o�;o�1n���8�4 ��L�4j�W_�}q	Ɋ]��9��Tv�:ſ�N�H���v�-V6 o�L���y�䪰v�g�y(}����ώڛNR�F|��} >��O�;���8q3e��~��������+PD�4*��F͡��+8:��mE�e���&v��vJ��Bt*��}w��6�Q�8\xX���@��q�#�ݡ}��a4��p�m&u�]�ď�ا�C�t�������~$~�c��O��'�to�1���A�n_��NTȩ�6遀��a����~C�In�x�h���آ׊Xz���Hd�$���g��a���d� ��H��};��R��]��J[�Aml���t��z9�/��V��w�7�u+�##߂	�<�_Mz��"e؎��j��ݔ��Q�����8%�PN���a�ޛ�;�\�����,<*L����/4u-:�2�4�	o�D$���kc߾����Rr5�7���9�{͟��H\� %3�� "xEE���)���߆0��{�r>p�����;��P-k,w��P�k���3��3����ӟ�d|�?��G��X|�3�������o�+�ص5bJ ����_�yʵaN��`�/0�l��H�ڔ�D�_έ�%n�O�T8�2��i����\4V���k�Vi���`|���#'����hԇ�S����x���xg�3]�"&Bb��C_��Y��<��t�bw�K��g�
�n���E��9���^Ɨd�n<�m M�XWC4⍒ػ���q�[��}�����/%~��� ���o��ɉ����&�Dca�6B0�z����u���l�Emkm.����2y���Y�bf�z�`�5?�J��q	�R�{'�K��Pv���$��#�GJ|ai6N�{)�z�x��G�+��з�瞎�ѡ�{`o����*&+8I�5��"]�������zĕ�(o2b��U�CG�!i�}|����I���h�vz8��c�J��l�l���	����8s�L^�)1�rK����.��)�"����8J[�P}(�$
5jW�8���%\�i�D.<T�q�׮p1�[07V����8z݉���x�����/�^��������o�7(./�����xχ?;�=qn�"���!$����u��,�a�ˤ�st-W*��D�LN�R�N�Ҁ�Z�j�~4�pT�-��>�z�F��Uc�V'&�=�У��/}-������<'_8	�oƞ�ɘt~��+��4��@L�= �����w��T�Ԋ��<2�d��/�Fͱd�ԇ+���2�wd0|�Z���Ƈ���P��69�C�;�!��.A�i��s� ���F�k������6�hz�oږ�r��&F�b�^$ǘ�q�u��#u��Z�ؖ/?�Hɀ����׊{a�)�qeiތ�&���`���Ŕ RkP��67\�3&���;x0~��:>���l|�#��ʳ3�q�̹�yd�9#�) Er�q?z(����⎛�'�C�̕�xߎk#-B(Do�:�"���e�7���sm��:w��$���4u���4�n�T�P�l�u��"�B�����ڳk�n8�\<s�<6�FF:K�'������ب�.H�y�]�@�2r1Y�D��a���6z�Hk�����ECB��H�C�5#@P��'�F�@�<F����ll���]{"n��XA�;�>�����8t�`�߻/�Ny�ɧ��C��w�����G����S/`& P�����'�S*k�<n)�e-��K	c�s�S�s���z5W �=h�%����.�SE"ا��>��8z�h��;r�p������s⹧��%L0{�&&c��C12q �,87h߾�]��}{c��E�aߘ"�V�{/	w�8�Z�2W2�������sBx�]q�u�s �R}���)&��B�F��C���H���5�Ph����SO��6�g/�� e�V���oߞ����T��8)�~�d�uU����v��y:�%���WG�SeowL�&�o������?�&'bvz*{���"�I������(�KkJ��+9)sfv>�^�q|���G�K��)�K��X�gh�p:��wğ�	��%μ|:N�|�� ����:8q��S6���]B��iD#�Wϥ!��"�	�B�4�߰��%���I9b�˔�`�vw��U�����5G�sU�ap�e$ƿa��M�ÑDx�FU獂��F5ϩ�G_ Q���9\˜�i��x�s��rI�$�&�l���wh�|�}�R�{c�C�U ���@_%jH�KH��~,�� �p�{0�?�䞌͕���W����7P��H�v�N��#�V7s��.Թ}#��O,��/�B�嶛�\Hh��G��L���7+ˬЙO$��\�qn�GG��x[���>��rR�+j�ܿZCvC4���O�S�*ZH�u�)i^�z�T<��c1� 1�E~2�U�Žfu�>p�}��?��cz_�3�fM��<v��Gr�-��~^S�<���s�v ��O�}g���qם�ĭ7���r��,ɡ��z�������}8�~��8{�48��.���/�cܻ<?����2��8�R.[�E:��qs�v�q���]�7G+���l����mʥ3Ѳ�^$�$>���RC��{�[���-��� 8��u׺E�&�>!���oM�o�7�������p�v��p��� �
̗2�}�;9����]�^���h6k�)V�r��4���5th� ]�����W�%�r��L?$��ZCQ�ua��/D�E��a�v��XL�Dx�8m#9|1q,x���2����N���ry^<�~���'N�:�R�;r��"C��-�ђi�g�HC4$�U�V:>�?>����}o���(�2'�N�*����gsU���N��H�O�|&���~���RR�^\Z�y1k�s6�݇�{���'>�#񙏿7>���0jy7eTd�[�I{^��hR2�6��1r�1n'�t?�#�Aط�T�=s��^�^4�nn�@fc�9������H���;�^%�����E��黺t�b���A=�ǰ[qN��ƣ�&S�Ň���UJ����K竦e/�K�q2|W��(f� LO�tiz&׬]�ޢ�=b�=6y &Ў�:�_{�zdp���"�#Qq������et��f�?0�:��t�&tE%�M�k���Q�L�4����}6D��!������>h�}&f/$u�L
7�r�n��A{���ٚݪ$ۥ��v�֐�:���6�X7�6]GUs��Y���16<�m�y�ـm��ց��5�֊�%�G��M�+UL�r�k�ynh_gR Kgi�YyO����k��,�rz�L�����:����^��b��H��(2�����aTX��X�����g�Cu� ��� ��DL`f���% ��2 io��#�ouz�^� D1PC�m�]�]x]�I���������[��n��]�����[�vl��ǎ��("�wS�-`	���
��O�Ĺ�3����[b�<Wp�z���C�Tz4��`V�D5+``${,g?Hw��f�����l���" �zw�7�Gbϡ}�>+.�ȳeT�u�Y�k��#�l��ߴ�2w�.���ڟ�A�¡�Jٲa�`����.
�&rϣ=.D{>v��9��e�} y�6C�#	3�fa1�ю�&�M�2�
�:u`v!�O�ŋg�ǋ���,/��B\8�Ly ��cK�|k��p-�
A΁"�\��0=}��Rv&��06g�[>�ub��3�s���"3�Z�S�&管�9;�{�S{З����Ls�Ә_�}�rKͯ~��[������������ZLM]?I�v�IPHGR�����9B�Y�%DmP�,�%�>N�� ��Kp
+a�1�^��$!���z^|[�h��0�4m�y��|n�{��w��)���.-�L<��7��Xq�HfJA,�~����D}V�}m�I�8��yG�(���x� U�d�݅�h�d$|+Sq䠎���H��U�v����Cza� ��0�M���ҥdp.�:����s��sO�#�4���C���~;���w�ѧ��G�|"�W��I&Ml[Bs��:�dtpR���#h�N�yW�@Jй��e�I{%��)�LH�wT�e�ܛ�s�i�l��A/�um���sg�_�B��o���������_���{����G�����/1Ν:YTc��LT������@2�.��2�=��9��s�A�[�n�̤��s�;#u����՞��32{��ҟ��'z�%�I�;u*�����׾����׾���W2~�˟�'z(V�\��H�t�L\��𾽱r2{������-3�Pozvz`�:#e��lt"h�>��R#L����5`H�oό�+��U�"�;)O���/�m����A/^����<ͅK�t�t,\x9�0Ӷ����G�'� v��e���@�X
�>L0�}v�*eZ���aq�Z�A�E�����)���-pDڠx�f����*��13"a;P�|�a�^y?뙧������h[�o~�����o�������T>�fg���
��u2�wru�R[��+ڀ���YrI�%*�R�� ���C�l��q��v�Ld;x�@nK �`�H`#��s3rD=����_����<����W��������x���c��U�E {���uF,�`} ���"�[��-rg��9Ғ��&�6�ܶ��mơ��������&�����2A����/ga�|ݟg��x��c����ܘ������ɓI�k�����>�'�I�rR�_�C���`��&K�C�N���n���v!�}��l�>�ZϺ=d�e`8��C`����{�G���q���ޙ��A �7Hc)g/��� ��r��v0��[O:�85$�`�n�իo� \���,?�v��&#�^�Fż��#��)���Wis���h<�څ���N��Jy�킏f#j��x�'F0��]�~��
2��Hg��M�#G��4�m�ҫ'�C�����6.i��.���^;�\�MgE�:�֮cj��*����h�IW���Ǜ�w�&�w:��~'CG�)�I�����4}��6|o�;#Z�Ml��ǩ�����c~����_��;������- !�ˊ�Y�a�N��[�|(@:�K����Dk[�q!9��G�L�ǅ_�)؊���h�=h'��3qif����R��a�у��M��)�寘�Q��󝖞2����Cqh��}�bM�رCq��Ǔy9y��?��x��s���O����-a2
#�$C�A���ذ�蚣���7Sv&���gcav.%m��`��Sˇa(�=
�AZ�l���q i}�Б8F�'GFc߁}q�����c�HՈ���]{���q`����C���X�����8�L=!K�i�,���I�M��J��j3��xC�~�a��阝��y�)WdW;���s���o�)n��Ƹ�����[n�.n����0��Cv���ػw"����n+�����đk0G�;��PNk�G_�n�tq)��q�%(Хأ3�_+�8�N�+�V�������X�_���` �m_2�C���uǏ�M�_�;�#Uo�����������k��k9�����'r���}Ai�;��o�災c11:�p��W������OFw},ֻ��&��E���BH��k����wh#�Ϲ�C�Y`�f�2Z�� �)(\����Лi�R&���M�x����8ܤ\2���7]s(�q��\л��~6�D#�Y>+H"W¾Y/�m��~��_~�+qzf-5�C�7�P^�W������
H����I���2��^�p!&mqْ174S$T
���X��.�(pe�W���a�=�˟�����p�.�ģ��V<�����w��2��U����\��:�T�J�-1��ŏ�wb�a$�`4���ԵV������+&�̶�z�/�����w���&��:��s�[/�Vn�m��m�{�4c��F�4���;����?�]Ҟ{���?.��b�8�
{Ɛ���G�O�ݘ[=��K� ���V�b���m8��%�V,����}�[n�&.M/Ư��_�/�)�g4*��gg���"��E�(T��sP�~����]��?��غO=�4�#h~�1>>7^cN�w���Z���hǄ;8��na�����fggbM�e�]�����SW5f!�w<�@����Z�9�B�տ�w��a���,�R�cn+MwC)�n=R��߉��gu3��_���[�h{_��7��3���}q��^L��8î���ĝBҶ����jm`(�_����V��֐&��E4��s7�`N{�����_}>���f�(�Ȓ�A{N��ځV�MA��H�(�:�ġn�
�8�C��Hb�"��):�0��p�2��HK��+�!O�ceC&�6Iz�����~��P��|M�*(�v�-ty't�zE$�4J��:c�7���s{s�W����p�	i�x�&0�T��v��j��tq�4���w��K(}H��rza�F�@�C���!��u�<L��?���ǧ>�����~:>��??��??�s?��K?�������_������L|�?���Oć�G��uG��B��1����t��A8zۧ@�e���`�ֆ����Q����ᨏ��z�u�]c�hoD��򎫷;3��(���Jccq���؇������w�����8rͱ؋�v�㞃�b�=�o"�õ�Ť;p�@j �c���(�Ġ�+s�i	�4�ڎ{Y��W�l��0��aN}�}#��;2}�C�O���:���췪���00��r�m�ȶz�0����W����������jjB�_^�W��2�3�'3���rk��v�A=fW�c~m���e8�����XƱ;�����|�;RO<�N֫]1��sr\zО6:@�=~�|Q���a,�Ihn�އY�	�/�v���:��s�E���b��	6�u��H�p%��e�7ֹg7�{;�F��{��=����a�V�/�n
S�y,}tB�9*�h�h�I���d-�Vƅ�������.Ė׾c�rV���=��'���\&?�f9^�D
�MJ���Y����S9�^�)�D�bԤZ���L#�,�3����
�R1�l�C(�l�v�Ђ����-�S=魦}�ء}��?�'*C�Pe�g����x�����r����v����(�V������#1r�xL��6��1�˘���.���D����F#FAĉ��8C�]I�/V�b�w)��*H�
X����2:���~$�
��c�Q+0���2De��]�[0���Z�@�*�H�e4ɻƳ�&1�ފ�-��؀�m�7�{�A�j����{����]���j����dwң�gi�3}!�hp�{'���_�kbIZ��s�G�D٭K�ނ���!���O�5mi�-r!�K��&,L��K�j^�H�7-�.���X������r,.mҖ�ѫ$��а�����R�jέс�]j��2���������2]��g;F`��*�h�=hH=0�m���q�0�������X��8�&A��Vs�s�/Ź��<������xw-+��g)�kwq-���Y����(���nW9v����DU��V��|tZ~�84V�5�/���K:��`��b�o����q�$}w�.�n@ب}�τ�B_2�(S ?iQ��9�&��^.��`�A��m�~�W0+�1�xـ: A�����J '\�!�����C�A�7�D�.�ѩ��p�S��{@$��u���({`%\(9��j�d�?�؉A�Q����5@�.�AP-Ԯ��2Q�H�"�����:ҰA�.���!��<�������R�X����Xٮ Y�ѪT� �}���zQ+� �Ѿ�����X��"�x�n��nM��t�S�A�m���c8ԮryB���WDl`������=C��"�Ա��7w���F�R�sS�켆���ߌ)L������_��ӳ+��Nô��0�`�&mK^U���g�f����׋)R��q�#��Sq��0:~aK_�{�*� ���
b�PGg�f{+�Ю��fbff>��\�����;=g�^���fb�����X��W"�`$s��6�zKG*Q�vź�5�pkM����s��LD��A�P�d9���@^��W�=���.Qĕ��вa��he5���ۉ��ո85�i2g/����v��,���g��"�����2���x
��g_�Ǟ|	�m�E n /x��N]�]�_ʱ(��׋��G,�Hvq)�����;X2i��le�c�n���c���ti�f���Dg�L�"6��;��1�f��;����}��Z��}�+��k�JK�f��h�Scj�-��4i�	ź�RU|�B�f����Tn�g޷��[{��67\	|������*���<"5ˊ\��g\�޶Ep �=i��c"�6��&pl��_��	בl��8������Z���i��D�sg/�4Gy�
���sq��qv6��)�<�O�i�5��`H/7VB�\�a����2g�3�ҨmG����Uf�Vⶌ�G�o����j�O����8s��8{�t,-��BMW�Z���Q�sg�ⅳ��8�{�N]:��'_~)�{�y$�4�~���)Y��q,��,��ׇtΕƹW��ל��H����`��U5�s�^��	�0������8y�t�p��@96$��kɼ��1������Z���x��*�c? �h�,��[j40���-�J��T�U���k	!a7�?W�C���g�(�*���7�l�%���sl�Ft����xE��lM4����7�?�'�� �yif1^x�8�4�n����Jll#+#���ׁ�"�y�|��3����u���U�{-��,���Ͳ��#��n*�ж�mbo�=�2}�����4]^�:�4����)�_n�-���A��t��.(�v��0'"q_�(�Su��$�#p����HSKB㾞���m�����Ĭ$2"g2�"ㄍ�_�a�F�d����5�A�p�!��E���'r����������grck=׃�:*�X�$���O��| ������3?=�=�\<���c��<f�6�}9���<�@�����r���a����-1�Z.;DY�����%��V�8Lz|bO.q(��a�?s6.�?و=�q�M:+���8�}{'cϞq�^�ᜅpO�9���`R�!��A�Hi?{� �b�����H�ǌV�}�e%#T�H7��Ǣ3�h��M�6�7���CG��,���ҁj$�>'�V��Sǝ`J̮��f}��LP��$4����8�+㒈��q�(��sNt���@1�=����<QH鳱m&'��T�[i��Lkh�#c�du~��j*����ā}����}1�I봋!�ĝf3K��6x�p�?�xCڢ�.�)>�Z2k�٬_	-Օ�u��l��2�IZe:�8��ş�=m�x+�)ǿ�Ax���(�i>g�*�IJ���� ��Ij�����?w셈H�  �C���H�m�S�T�2�ULwY���&%��W��֧=��@�}T���>���k�'r�������=H#%�,!�m���46n�]^�}bY!�	��}{&���q�ر8x�H";q,�B�N�[^\@9�H6:�'���J40'j.�B��J�>���B^Im4��d2 #@ܿw���t��pLU�X^�i��t��ڝ��V����H�Ţ]k SD&�,R7ʞ���R�={&bx��_q����2�A5�aF�Q�@ׁ�^�=��t������X6w̱=��Gu��s��-���`�ю@!}yi���&��}�r�����ՅŘ�p)a�>�'���F`�#�������Q�6�&xb��"�沂 �f��:n5��ͣQ���zNYʈT�& u͸{���@��r�ɔ�����맒��T�+��YE<��w�lL-L�E4b���аG��E_��r}q�ڣq��7����&��<Z!��B�;����ޘ���V`Bi�`�A?�xN����nW�uo�����K^�H
2��#pr�4�í=���]0`q����Qp�J4ؾҾL$y̫���a���.\7�v�X	 ���)�r$#R��0锸��H�~n��G�}%? ��֑�8
	%E7�V��p�c��G�Q�d��Xv��d68H)�ȉN ����G�����0u�R,�F;�X��ɱ�_��b��'�#)�?��cv���;��}*5�AT�I%��QA��ђ�HL���ĬK;jr�,G�������oT���s�b?L�h��"c9�is��l�s��jl�s3��)��i��A���#Gcr�~��/������	��k����-�m�����3�睺؆\Sf���(���3��i����O�]�ݖcXlk��\]BOM��D�^i4`��9?ftl8z��S�s�8�7��!���ӹ5�h7�c�,_
'����&p%�OL��b�.Hg���� >++E�v�h�1�s��Ļ�;�P�7�M���!n���a5{ڬ����'���TK�xf�"�߈a� �p�F� �b��zi��jԹWCzU�S�*���XA�s9�-�s;*\2�B&�J����S/�ܧ&�K���:��
�P�G�by)H��s�A��|%�I�H����H}�k�0�drp��l8
��u ���ת����VE"��0\Ɉ�F���\F�b[v5���wJz�;�s�zJ�z�"���H㠦��;�=B����pC9�\'��iT��ڽh�4~i��t^��^�ŵ�X�\Ŏ\���!�H�x�uq`��\����˩�X��$u@ُ�)*0�*�ј.����~��wTR�����]��q>��۹���8宵�����Z�Nw���X�U���a��#z�*t����H�=��/��@��P�ߙsa�vӫ����ֈ恔����˕���b̞5��+ ��0�^�6��v��|��9zrXCP:�f�)�'�:��E�j���T���)�&�m�~-�1D��=�Lt��!$kX($�"uq�N����5�\�D��6�Q�؍����qH *���`f1B�����y�+Kq�x��E�&b��靦8	�Ѷ��|;@�z�c�x4�O�����o5��cu���&���;����u�c|�ٝ�<��4��؀atbsq.�a��[�Q5/�&f�0��ne��Y�f挜Y�Q�n�"��DG������A��Oj�7e"w�
�3ys>�%�"�eT��\��CP�.�x��)�[ e�c
��ݹm�	�!U'u)�v��4R+q���]���]�ѣ��9n3�JZF�=d�٭k���l�K�Q�]�cص}0�@�b#�\ �zQ����q�ȎM�j\��Xg7f«�6���ev���Z̰�P�4�$���ؒD'��t{4�E-�8
:,�N���1̵Z��T����\{�'��&ѪFSu]C
�3�z���u��4w����s���إ8a:j52�2��8���7��v"�wc�co<���a���ro�1�8�s>*.8X�ŕF<��3��G�g/�K�VR #�6Y��K!�MS{B�+�!c��NN�z>����h+4<2�&Y��=2�f���\��q!��,S��ٹ4����J\ʸ��:��z�h~6�ip&|�� ����:������s�Aq�A���jCc��&��\
�{}0�^�
�!L`xcy�~#58%�uS�t��9S|��j�5i�rЊ|��r5:�E���J!N�:����ȴ�O�������ٟ$|%�ː=/5�rC�eE#)���9í|OF�	o�DtTMҘCCCi>�C�F�phq�=�:{gJ͖��~mr����e���"D�	s �!F�)�3C������
Z�Rl��ۜ���7�1�P�W�gb���u[�y�T792{�U�9sc�S���^���]d�W�:؋
+�9��9Pх�T�s�����%>hnv�{)%�$D�����l�U�s�c�z�Y�@�TC�g��k�K��]u�N�e�V�`�qC�A�j\�i�J]_z�d<�"Cԧ�2����F�H�4%��� �*Ϻ8�j!I]���>�l:�V U|��&'���
p\�+K3eKQ�-��ڼ�sʽ�1#R�1s9�$3Y��y0HV����i�]"�i�_��n�'�T�}]-T�M�i���iW��9,���;�u.c280ι+���H@޷c0	ȉ�p�؁�wQO�"�>1#ߪm `�h�Dq��
�����u�1}K��[c.Dㄷ�]��XɊ��\�W[h���bvy�:/�4�,&�L����8q���� ԦJ�S���[�,��M�s������5�$Yh�o��4/�YRuq-{�t���]����)��}��-Aa��j�2���ې��j�1����+o���xS&R���ӌ�"r0���rO��:�8΁Qq�o9���^e��[� �~��Կ>���¹]�}�]؛Ğ�u��
�i�r\�>�8,9'��D��wɽ-lEW��DZ�����@�.5��q�ҥ��==55�fY�x�ƚE�<�2v�b�h�v����byyƁ�9�ӡZ�.e�Y����<�Le��l��U��e���/௯et�Y9�^��M���r8�L�ƭt
�5�@��N�Զ��er�����n.\B[9��O���n�4�4v��DA4�R�P։޳aՀ��R�|�Q�f���ݎ��`�g�j��o@$��e7��T�Y�s��`k�orm3�tZ/�y���U��0�|�b�M�����hL_���g9��%�󗢲���F�Jt�� v t��T"c��旋L+�)�/��e��Z��%(����iSF|�|6�K�t5m�x�vҍ�\j���ċ/=I��Lg�x�d<������B|œO?/�|��8^�Qpbc\D�L �I�	�j�E�W�-uQã��~�Z�f:l��:m�)}�,�j�2��������.=��,���!�	��ŹJ��T�v��2����?�i�˹����;0�-2C*h��M�:��o7�&�Y��n{�]�2�Զ�aK��\{�y%�+;1RE#@Ů�pU��cK�]_�H�%a��pw�դ���:��8��,���ɗ��ًq����p�|�;s6N�x*���x�x�4�/L���cuF�6�L��K�9sL��~S1ɼ.�c���R� ����S�>���h^�n�gI���ч3ӗ�����s��rO�ܖ�����*�����s����œO<�N�L�Z��CUb-�3؎n2%*��0��?F�Gօ�4��^�G�X�7�/�^�u�Gq������� fY=	��q��ٸx�\\>�q\��]����/�8f/�t�(�SgO�ӏ|70����Z����d�B5��	�����2\gi_� �4�V%+́��}n�� XɶM��r����TƱ��p-��N�:��{�_���(�}�hy�K�?�^x"Μz&^z���������W㋟�������x��_�&Lf��7\�/��v %�C�d�H����Y~�e��xWo�C��anc�bg�:�:mS�G-�F��Ӕ�;$�G��?�3���s$��Ҿ�}y�~�W�WL��� ��$`�V����~4�����x�,�F�U2�
�;�c��c�C��r��t�CS���x7@��lƍ��������S�x6>��/���\����Ξ�a��{�k�>L$򳫕pg3����T����$��z�\<������/}�g ��pO�kr�c2s<��@v������8WBgo?����j<��ӱ���nű����%��&�%W�������G���M�)���'G�
޲��B�!��IT5o`N��g?����R�*�~�>��?�'��#{��rH��v�����G�1���}�rd���ޡ��#iviu��?����'?'H��'�����C<�������P�#<��ȫ�˔x@Y�iS�\�����Ϳ'>�㟈�}�Gc�J۠b?��3��s��T�1@p�;p��v�k�;��i��0gw���
��h���*+N�\ߎz}4n�햸���Hc3����6������s痲�%�"����:��tœ�<��6rs�0p��{G�o���,�;�m�2L���9�1�e>J�e7OGp���
�6���
m@ZdQ�m6�{�!h���0�^sm��Q�����/�7������Ř���� a�-��[;�M�{{b�80�OM��4�v����n�mP�s���{մ(�()��x�gSEa�Ѯ�~������s?��80�����:9�XLİAY�z�L�w�����g�cS�u8G��PT��-��JT{u�@D����X��%L��J�7v��߻'�����G���8|�`�A~*�FG��g�������x��Y�Z��ND�	`�d�7�#y�+<C���ڌ_��O�D>���X�:�����o}��d �%�9��M�윥��^g���	��s�u�3 �A+bz�<�'n������W�	1wZ]������7z
�wB~~�h��28�D��V�H�z]$D����Z����/���ZLdq}3���/������^���<�d FAD�RZ:!�lW	18�䕡������>LL�}%:��������^<������;O��}AL�-��Y**����̀ tlV�Uj&�)9R�œ��?}���*�5�+�\�7C1a��ި>5'�����ۅݽ>�{�~ժ�1e�)8�����c�ݞ}�_�n�����;�̈_�t����hBSX	]��`�A�j���Y�)�p�������č�@˛�|��c�JW��neG[;*��#����1@}e�ٳA�R���E�sT���/L�ʼd u�����2��_���ܟ�B��=XT��B��GK_	��Ai����:�̙ˉk�E[�,����o�^��e��#��k_E���D!V1�]@��`����;~�'chnn������8�	���8��?����c�cY���d�y�[o�w�{GL�T(�%��Ѱ�Μ˽E�|��$�kN�����w��.���J��q��Hp��T���9��o!����R:��Z�.�^K[Pu�;6����'���Sp�F�S��bC��`��H�@`t��ڡe�ԍ ��GC��H٩���������P�C� ���Z��^������W���v���UP(�Mm8�/=�s�\ԆtE��ހ!�#�_��1��E��@=�V�k�ә��)�v�V��LD�]ϻ��9ֱ�]f�sסpdk��9�~%���6��ˈ�yi&����?���:����Z�LS����ݝ�<���	P2�u��J�;���3��X��O|$�z��i%��]�����6}jܴGI���gy�@������ʠ��p�ZO���-�&�~�V%������?��S�3��_L�T�
�p`�]�%p�[�7ω��'q�����/�������6`N�g�S�Xt "f`��{�$.MG�����m�gԳ���[`=�_��*0�.��x�s��/q����G�2���ǁi������D(py/�S8[~L�kH}�28�x*F�~m;��Q]a��	�.�qU�������J�!�~�����qx�7*]g����H;��Jhn�lA���/�������V<�ԥ�ȠB쯴��;n����㦛N E�!�i8¯
`�{�������L����[o�9j �Mpz0�i�T�:��ce���������RlV�ba�76��� �1�3-]T�'>�����S������iO����d�y;HUMąZ�f������:�$x��H�d�IP:��cnq#��o�A��_�_�� D!�j�K ��S�B�� ai�d_;�+����ƣ�K?��x�o%}��l�2��t�ps�0���s�����ځ�a��=:4D����YM簰v����6|W_|��ߏ�����x��e�����FW�dYpH�j$X�/ӖYv�8�o������>��|F "J��߭+�=��A��	eC#q��乱�4���;�;�O�lQ.W�O�
�z�ŗ����x��'�Ei�oئ�-)sa&�@=�hʕ>{�|]��V0�R��>��]q�聘����QG��~;�q����r��Xk,���X'� u��M4qn����R�r=Z{B��k���f���~2���a8�04r��mj�-�x��+l�ը�.`��fo��w���Sڍ����� R`u��&Ny�i
�pv�5͙��Ȼ�3?z[\w�N��Uq�i�+2#�*��̩�N�~��s������/L��-`Vl�G�3>�c��=c�1۝�_Q��̐C���DC�{�K���Ȳ�E��p|_�is���עB!� ������[������XꝈ�ޱ�A
8�|qe�r �w�qc����D\s�@���^u��^���)A��$�X� �:N#U�D8�/#��{����+�;�%L��������yCC*�6��BB�(U��^#�"�E�2���Kc�P^�T=|x_|�S���&Q��&�%�@x-4&��=_:]�M�)Ã\˹(z���I�u;������'�5V6��Ź�����{���RD�^�#���1��!�]v��}�V|!9ʒ������cr�`T@�^P�J_�x�ߌ7^n��O�%aaRm�,��agԪ^T��`�+�k���^�mֶ�����?�-���Np���˱rι�BΑA0�)R��%K�d���k��=��zu��x���dK6ER#@ 	���\�B�r��r��������ުP��ϚS���_�g���{�����ٴB�S�lR<I$2���NoP�F��������}D^4
c����U�amm��]�ӡ�����fY�B&�U��d-4��Z�0�l�!=s�2��>���8�TE F�V󲠅�ó�Jx�ڨG#�`Ʈ�B�B
�h$���|q�CI����S�P��(�
]$Y���۷�����6/RyL
hD�ºk���kU�w�\�C����C{m�	�KV����?q�-�벢�,U�1�y�c�E� �<�\t��H��1!����M�+�Ϋ ���w�����o�f��ڼef���}���SϿa�s�VI���T#A(�z*+�R
Ҭ����|��������1'�/-(�,B�����ɂ��{��'��xK(==S�<��b�8s�=�gfd�����(\�
/~
��S�ө9*��+(bD��?�.�"�!�Y���V�Z�]���sf�i��,��yқ��Z����Ytf���l3���&#�TTJ�%�M�J��flDn���+�Ky�5kJ�BVm���
�t@f�	���H~\�D�)��UV���\�jv,�d&���v˵5���p��I�c�I�޿���##s�R/�ե.�&�s��ɫ�����1�&�Y ���_� Ls��W��
DQY��#ό���xf	)8��]t���U8S���"���x��iV<8�3@n0	)RT����&���!_t�T�H�0�"�LF�O�فdVߦ�)"E���	��	g~���V�I(7�z�*W�@$L�,9_�Uv4hP�����w�&�����-Klj��x3g=�|8�׍�*	+۟����7�Y��N���kv��^cJ�X��?o/����\j[�-���)�ts���H�N�?o�ī��WO	�E&!�2C3lk.ik���W>���_�gy{�����w�S#Vjjv��ѳe	$B�+�3^�
�&���i�V�z�I)��ȃaJC��B��4�)���ƞ�����z@<&0�II}�L1	!�Z�ޣ�D�"�I����Jt��9��{	�X�«����.�@L�˙Q�h���)!�C/ *��5W>�C�0�^�3���f)S�CB�b�fz���Lb��&����d�%(��RK4#p��-��qͯs�|��q��ͫ���0P)����j��*�)<E�b�O%pC��O^�?��I�=�BqƓ��	Ѓ�p�l�<0 ��%�t�/�v�����1^���,�o�='���'s��*�0F9�Z9�H�}��^�%��H�x��q�-^4,`<�P�$h ��נ |�?ƛUR������1\�������֐�FY��Z�S�i�ǠbL=��fu���7�'�_c��Ϸ�s2jU[�z]c�fȇРPW&Ȟ�kF�8���]����a�A����H�Y~b�N�����S��b������~�{`�]����[�<;#�����Ȟ}n�,���~��-Z`j�S������kUX����ۅ�	�0�Hht�]�sT��I9�!�#7ìl����
WB���H�6���%䀙��b^	�9M�x'����d�`��a�93��o3�#����x�(����g$(���B�C^�F"��?O��҅J*��`	�o,_�u�h����zu��8�ј��� 5M�L���(o���;ҧLH�-�ĩ����ς�^��s�C�t_ck�8ilT`�~M�DR��Jɛ�1�S��.�%�2�����*� 2a���2��d���?b~��Ǜ��Pa�2�l�I��X���yy�X`�v�"{8�s����dv.�yN��2!`kY<��v�(PS�������-��B�$�+{����2b�G��e������$��WJF����x� `�3"��:[ݻ��Q�~фlQGI����o��o@�=�7�1��z3Q󶍋�J��������� ���
`��&�J�{�Q�ݩ��E��f������ŝ{���_�P��+iV<g#�Cv��q���m[6ZNV������~dC��g�Nj�O2����j�+����ْ���i{��lp� ���3"ԔwAIӦNH��d"* ��0�����>m�2�s��B@�&Kr����{�r_<�"�蔰�>QGĀ<x
�����J�d���T��q�C�a8ذ7�@�!��1���g^Y�b��0�߁I�� �Lk�,D#�BP�NoN�u��]ym�a>�rH,���>k;@D�&�Z�ӽ��KT�[����}8f�ufc7�}T,��f����ɣ���.���\,z����i0x���|<�����q�C+�Y�2O,=�W��-�VC1<���]R��^u�^�4�����r���,�{h�1��H��1C��/�F�P:_�����u��q/����d����`�X��D�C>�W�>*~���-�q��ϝ�W<��~�y�/ J�
r�8��6����\g-iy�����O[�w~`҇��
h梲��57[�^@�`S��iĒ���ͧ��x{ɨ���}�7y�V���b��<**qQ��INJ4==�L h�i�H�gCh-+A����J~i�(�Yތ
�]�zZ;,+��W(.�B�C������/���r�E3�S��g��,_�N��L�<��bU
/+(=�J2A��ZB%W�����F}#.���z��%X�/�c�j��C�>)�_ �[��1Uq�&��0,.e�)NMH8��8��K�,��Z��Ufއ�,lZt�y]DQ��v�j�7̿�r��S�S�D9�R�E?�Űb�W�B�������ga���%nlxa1)'���L<��!ʞ�^"l����wݖ�+R.�����������&��yF��_���԰�8nM���(s�P��BZ��F���P��v�$^����k�3D�
�x���I�ѓT^��4'9���*�S�pE���S�W�hUr^�%�i[>�Ee5m�괵$��-��lR /�B�_�xU�������.��Mxhe�,�
���F�]�Gd�o��|қW8��M���e]��~���/al2�F�D%�F~=�V�k��z(���������Ĕ�a���c_j���d��A�yʲ�Y�0^F�Ҕ����%Z���]Ͳ3�I�������%XLz||Ҋ����I�2c��i�Y��{#�c�X4��2/��W�샄Y£��̅��*�ç��}A�.J�8v�\.9C��0�!n�.I�(���F�F���P�p[�='���@�k�e������x� I�S3e�L�X[Sɲ�qk����,��R�z)���z2}7����ly6"��8�������)���B�8��tAs���y�7�+�LIF2S/��ê�9*�L�sFy��%)�9As�Rud�W?y���o~����>k�{���|����'��7-�D$Gk�+k �,}�Y���.�����o!?��u'�|>�4���x �7�M��Ҥ�F-^��\S�7�H57-�sim��Ik�����h������ڧ���K�M���KUFďQ�9
���0�^fgQI'�B����.# �/�፡��.o�_��r9�͓?I8�0=�1\cM#}h8��k�fdl�v�u�.�ے����HX��-0ɏ`[�HL^A��el�N[�d�=pǭ�j��L��{��	C�b�\ʖ�t��vy�	[��l�W̳;n�h˗�:8]�gΜ��r��r�&�|)���T�{��I("ȋ�O�,�Il�
oi�

8�u��QJ�a/��$Dwx�uΛL�w�_ʏ��X�Mԇ�D`��ޠg���T��N/���y�%�dT�Ju�S̐�b���+�.դ���lԖt��5��y��5K�l^�B�֋y�?�S"�O!15�J�h�V.첥=�>�NR�ptx�u�@У�J���O���~\��K���WFC����F��y�B�u�[��6��J(�A�0ψ�}�����G��6���+�m��^[�|��]��/쳎���L�dŉ�����Rт��֩yrE������T��7��dB�]TLДR8�X����y�i[ؓ������&l~[Җv�l~k���mqw�nܼ�>��{l����@���٦��Y�A'2�Y�?�u9�Q�L�����B;��)z���X"�,��}�*Q�s���=x�	�$E�p$���؎-���UK3����3tJ_8눅��o^J?Zg�<i�g�ٛ{O���o�?�ǿi��a�)NZ�ȴ|r�e��P�r��P���6'�X.(N�cV٦''
��1Vyc�J*j;�S�J粡��H����u���Y�ĺl�f@�
��&��o񠗇�/!���%/4�?"$��H�$�k51�!�ҷ��?"�����hI�w�����we��P��ǌ��ω�C��nHF�Az�9���#bu����lݶ�nپΒQYp�PYN�
nΜ<i/�|��޻����fE��Z޾JAN߻a�J���|��,=�����v�HE�}���yxO�
j�G���[T�����\\��ț�'h�,\�i�}�������g���x�m{�wlt�-���{�]�m�knm�B�h�ڔ<Ȋ�+f͙Vc�4��]��_���ce��6���-�ge��\9���_�W�R/c�h�ˋ��ڨ8���T�3�o��^��ݷ�ڕ�VUd,�0d�������U��%�+e8�g���Ӄ71;=]�o=�����׳
�˄��Y����!�ۍ�6�k� �L�b���{uyFn�I�X��Q/��q���QЀ�����}���x��b5&�#Z$�?�'�Gmpx���s�G��!�v�[-:�����d:amT�ŭ�-k�͖`PiI�K),B�xZ������]V���5W֡=��3���r�*�z��Z�^�u��_T<kv�"�n��@m�
V����D_uEt����U40)��ѻ�k�n#\a�+�>��:y,��/�2��BSJ@C%��#�
`Ex�2m�e�D��>�����������)�����̘�X�ؾ���l��VɆ��L�{~��ri��'cA�{p����cldt\.rFV#�s�y�&�䃷�Z�[)_����Q	�,�K�}���hh�fL9��)�����I���`zOMǦu��C!g�Ⲽ{zl���6���6�]l�ްѮ۸�;�����H����_�W��W%g,�Xtt�ؼ�Vkn��޽�X�ȸ
'nS5z<�Sdn�kP/��d��=���P��yF�G0�ⴼ��+�}���F�ҮP{^��y��?�,�����9�'�;-�a�S�T�Jqђ�F=BN<��۱��ԃ��C� *��{^.ِ��ꄶ_,�6��_ROW
ɿ�7�$�vOD�Ch�����Tf��	J>݂�~@�CA��FY�)۽�NZ�=c7�r���>8J�SQ_�RM���vXqNa#s�>ql�"�u_�m6m����]�'f36\�7*1������$-�l�щ����~�Q�#���� ,|�rK���
�A����)�Y���U1C�����BW&�����3X���!Ĝ^�t�r�E��֙�y�/Zb��Q���7�R��FQ5��ޡ���P������R�7PT4�m��V��G�m�VYIfa�ko�_}�'�֑A�8�|�֥�,a�V,Yf[�l�@w��Ĥ�_����B�Z�c7l�d�D����g�Q	�,~�Z+�P<ў�%B/������KC�y���E:�ct_�Ra��[�Z��Tmb�b�l�u-X`���Y���e�����o<n?yu��=~�.�����1)�y�ڸe��޾y�-�枃v�¤5��-?�zA��8��A���{+�y]�	i�򡯯��o\g�̴&����|Bd�����WbWg}]�$Hr�\Ѵx+O��Д���V�.�ګo�c��1��9��Y_����띃�'�~9A<1J��ҕ^����� "W�3 �̪%����H�b��Wpoc6"�����q��	۴u�-X�"?c���Wwﳷ��]�r���#�썽�핷ؑ��'����ؾC�������3���C�G���{�^|}�,�!۽��M+�Ͷ�Xs[�N���^�e�'Up	�E�o	d+�����xRa`T�����i��D(����T&l ��VV,�k�4 D3]iʺ��vێm�Ź;����1֫��#Д�1��]��մ��O��M��9�_�D��4�����~h�R�3����D�S�b�u��᮷���}����vr0o����⫻d��IA',�I[�<�>[z~|�.��vݦն}�����и��2��R"�����p���� �	���e�|¨єH7r�XY���n��m*x��ڛT�'d\�-#O5N���s/�c��U����ь�D��-N�#zg�V,���v�`�<�o%�LH&�/��5S��~t)��2��v��U��)e��L�x��;p���Z��%�ʶ����7S���^����:yʺ��-�M����I�����^�=���G���tQ`l�/����";�<����$�͒���ˑC6���ؽb� ��MzN� 2�nٱ��D�	��� Σ(1�t��\��g:�ۛ�O����v�e{��������ヶ��i{����@���!{��)�s�;7lG������ۅ����#v��	;}n@[�9~F1������m�!��r�f��� 5�O`���P�)PPH��{m���m]>�Vj�bA�-_�jK��l��o��ź]����j�e����U���^�k�޶��"�p�J[�k�Ο��	���dI�W��m��o� �Ђ��䅩-T�Qx��ɲ���٣����k���=������ZsW���������{���sVK�X��^۰�O�c혵�f�[�YOw�ϑq~p�^�5V^� 3.��L�ȂڊID3� 	�p���?��IX�pNe�jY��|�&c���Є}�o���_���H��Ǟ}g��'���1y|�\���%--�Q��ϫ�Gm��Ţ��^z�%;~�r�p4�7��_-�$�S����!.<�E�u�5�^�� *�Ж�Qy��^�����d���b�<�
���Ln�c�٬�F ���f�
ٟy�����1�P^ޘ�>1ti���Vя	9!�a8OxP��%W�Ui�I���[�3ު#���Y�b��q�
g \��:�XUBr�����ȧ�k�O���'ߵ�Gmd��Ѭ��"�P�3-�Sѧ����t��S�$�r���Y()yT��--�K�k�	�����!��4��	,���XH&T���K�X"4Q�"O�R�#��C�֊r��$�
?�����}��[�#=�«z~o����Dk��КΕ�� ���Ph�v�w��[�����?������@�Z�%�̳I]OD^�#����2�B3�� �4SX"���Q��ľ���lQ�im���҃��=7X[�j/>��=�B��CVIvZ9�a��o�W@,[��>�������-��=�#?���֢_s��W��/?�SsV��9ߨ�UK*�@�w>��t��7ET���O���d��g����e�h5;p����˟ۙ���f)��bO�\ߡ�I��p��B�ce�֢|o��i���>oٶ��o��<���S��3=듇�Kb/'d�X]7:�,��P�UW�:�3�;a:�\3�ׄ��������5c�6���o��6�\lm��\aܚ��o���lG����<i��?����.�%��r��W�ҫX|�`}E���B��
D��#��_��_*�xV$0ak��К���d:�~���5�'��	����}꾛���ݖ�Qy�4�0��{"8-�t�`����K�H�P���﷓��YX)^ad��ҩ�<��U�nS���Y����h�N
��3P�������k�R�q�2[��ǖ��X6�8�
X)ָP�qA�?�O{/KI<�z�M�&
�U���c�;`S���=��̣�pa��>/Ŵ��bV\!Q$�k�daAG��/��g�mm6%�T����]��r�L��Q���t?��3� ��a��fz�+�����U��-:h���Z��..�x0�<��j��K��^yM��و��Y��T�NJED����cgUV5�|�u�"v4'-9�hY��7��x�+.�'���
��c��f:[�|"! �2�`�l^�<�l�{�$�����w���	ُ�g��ٗ_�)����OJr��Ek�V51�Ŋy!�t�l�V�ڧ>����:[�r�O|��so�ŉ� ��%S
�G@���J���@�'���0Ry���°�)�'Tv��8�j��|��LI�L)j��N����)��P OiN@S���{;C�}~�B�3��v+ʰ�a-}mVy��t{`�T��'�%6�>��D�3���/��y���q�a,���{'�S�ʢ����'�c�RKK�}���eY.�3�WB���+��
�6B�s��šI	x�[XV��f��t�*�c`d%�������mN��\i�3�$B��^l}�f���l˖u�q�j[�z�-[��W?�ikzbLr�|�a]f�*�S`*ZIK�ѕ�!\��:	<�L��X�ʒ�ZAB005kϏ��3�v���83h�N؞c��v����h��\������eY��������l&��<YT6�+�p��^HtP�i�S� /�U������������g�]�I�ZT��.	�
^�O�#�o�:��o#�⓸�L˒
d�
�� �������]h���/�����@��P��_+a���\(cc&�S��u��_�.��I�^��[e��8����,��ZD�;���O}�~�^��h����{v�>�C�� T�T,w�����Pd�:�'�DF����/��o���&�@�&�ġ����mh|R��<���Q-�ރgE�.`5�XT�'���q��P�x 4��ͤB$��E����A��pY��O�D�R�!k����7��$�9��X*�`AO�-kW��[:�4�t{g���3�|t;���BO�zt� -@ҿb�$V�g��r-b'Ϗؿ������e5����o��n��'�ᳯ��{�X1��&]�W���W
�H����_o�\��:r	)���\����.@��?4jϾ��=��N�K0�n�i�rEW��B�0w���M\2������Is�ђ�>y9[6/��S1l�=����η�d�Y�������e�tF�Zv��f�Pݭm����6oA��������^y]
��,��Wޙ'>��\��zP��� �(:��DA]����7�V���=�D�6�]b�q�]'�M�;��b��o�7Y+�_Dy`63z�2U�cY�%���m[�ٍ7\'O�dO<������)�q\^zN���R�Ej�>0�ቈ�F�� �l�O���bť|I��U�{[K��:{����bc0c�P^f\g���B.�~d��R)o�-I���>f��u���M��W$?{�N��T��g��ْ�*S!{�i�HB+C8�W(?M���J�cT��K`_��� �� +2��aZjۙ���,����!��usLw��Q����J�D-m�jFr�PIc�|��=��^�w�,� �F�tN�����) ��lx�u�Q�l��b�}��ઊNX8lQk�}�{틟X�S���}>_�V��k��+(�E^nW��\���h/�:j�}-�/�����a�������?|�&�����&�(~\��l_����Λ�
ڊb�v�+��
aӤ+���L�S��T�칟�l?~�y;32e�D��[YB�,�Nj�%��8q�3C[�6z��Q�2�Cr�l�q��뭳��^y�M;}����I��\T)#C�^Ϛ���L�Y;#$Ne����mL'�Wx�� T	�.�� ����T��*<�+�����@�Q��p�3��AdN�׬O%P���zm����"�y��lL�3}��C
���Y2�CB�K��ɓټy�+����m|rT���J@D�O��T�z��?$���S��_�f�K��+���'K\�mldT ���Xth�
\<B#x2'ŀ���<�{y;�|�X�gkW-���a;~򴼲�$U�*���"s%���$o��_(a�D������P��HT<�m��a��6�b%�]T ͺ�>g�ʙn��z(�ߕ��x|Lw�D����Y�%Y��KW���������(!���A��[��c_�����.���8>d�l�%ҹw���K�n't� Vi=0<>%z���0j��w�}w�b񪮥�v��۵o��������Ā���K�x���Vœ	��ô�4/FV�1c�ޢ<���+��|򚴄p��ESaڔ@�& �!���m�Tg�>|QaQ����&&�aR�s����S61*!�P#�T$�Pp=�,�X���� B�p��t"Tc��J�zX'
O��Z���Ö��=��o4�e���{��5>%�@�S,U-��P���3v���O�D�#�l<<��_& f��u�L��0��`�m�Dޖ@I��z��%pӋ(�:-�|i���H�Im��q��Z�R�3��:9�6	��f�t���-*O�И�
Le�6��mph�9f��\��9#�#R^��Z%�eP���$<�P��_�f< ��I�h��sʈ��~G��6[�Ph^���lN�������z�1R�Ј�b�fe���({�`
���0W.��!���1��� "�9��m^<\��"~��w]=��^��f�˺����6���k��@/ca��bی@�V�Wv�:����u�6�'PH �w���=|\�|Z��V+L��ά��YG��' n���C���k��3;��/�m?{a������8g��-!�)�MKq��Z�a��G�*�I�dEl��;c�M}0a�� D�(�*(����M)LIP9U*[r.����V=7SR!��(|a�>�53�s?����� 6��R���g�/�r&��M������T RL � "2�"��i~6��5���m��t��ćfyK3�i��&$�yK���b�]\|�R�ѥ-�|T�H*��J�S
q��	�Z��I�7B�Y�/a�n��('�C�,����J�h�c�<������wV�V^��/גz,"��GEe:�3[��xj3gY<�i
�/�朼@f��f�_"!?PyV�y�>�3x�>��䁵r��c�/���v��$U������8X���\��W9%��6j��)[��,WmxT�o��A�Ek#���$A4��$C.'�e�My�<�q��HWd	��+V���}.�q�)��"�q'���A�X܇�gxt�v�s�N���z"�W1/�z��nҡl6�Q܍�K�k{�v�[��YB!�z��i���/�w~��7�:3��B�M���g&GlL
�h�|�	�i�-i�N��S�֔hG�E����By@%�	زQF�f�&d�����%�햍U�=�T��̒���Y�$�7�l*"_�*����f-{t/<�9%dIf%`4;����
;�E�N�?�'��� ������\���j㘅�������ڪXt^k�t�{'lق�z]f�G��W1r�	�Jx�`�	�ג�E=m�i}e7��t����Ǖ����yNtC�{���t �S��I��=k��UD V��E�۴�׶oZj�WϷ%󺭷�Y�ʭ4��ӫ��������M[K�fz[lтvyLuPr Ϥ�ݽg.���'��]N���s���%�� ����y��)�a�*���7ۣ���n�u��^�L�ͷ���А�KK_	�ט��lqWR��eݵ�>��O[����]���\*nq�Qp.�mP��/	#�>��/�e�_��{
��hk����6��t6�a�b�;��t?��F���:
�A.�=�N���������q{�Ճv�����la����~����7�g�t�\�%�([�u�����v��er���g/�j�|�9{e_���;�mӪ��\_2 ��ŵ��{�M��_��-m���������k�̛��/�T�.�.�C *t����S�5[�6�3�{n�^�c�uu��;p��=�ʛ���E��*�M�X��⤬cٲ�Yki�؍��`[6m����'l$_��¬�by�Sb]B,+�(|�l
EE�E��-���3�0�RAxY�;+0�ߜ��KxoܾZ�&``z>�����7�3/�iG���MLH$�X��%���i�,���؟����3v��U�9�j�s���1�� ǁ��$o��{��B�@Ί^�'���+a�ub�n^�ľ�Gl�N�QUq4��S��dޞ��s�䋯{��O}�<�zwܼ�n��:Kd���~f�?��M�^呮�
�
����$�_yL�N��{�a`c�����_"�Be\(>�9�>fj� ���E�i�Zy�
q%T§��m&��c����'>�57߸���[��K^H�固쯿�Ӿ��mR��L,k5<l�W����z>�!2�gB���yo"7��|���p���5�dzM��V�^'��e�fZ�Z���7m�?����E #���M�v�p�7:�I:����3h|��p栝83`}����X�B��б����C��"��#ʆ�K}�R<R>4����s��HN�UQL8S��rkɀ\��b�&�zT�;6[g3�S����w��9<�Q	#%���R�E�������ꛊkg
�l~��v�z��G�2�mK�γvY�ɒŋl��>N��##���qY��]�a��u�6�������֬Ybٖۯ��ę~}$m�\�<Ѣ�FJ���&���6vWK��ބc��\?�������uد��#��7ټym�Ƭk~�%�s�ڴr�2�:1�/dؚ:�^�k�ܱ�>���ͷ_od	c-���F��C'lx�$�	�����6x	���z�,�A!���xHqbI	.�NT��laG�~�K��{n�j�uE;?4.q�g��e�T̖�MfA��tR^G�mۼ�n�i��v�uv�7ق%}>"��7��{
[�m	 �5+	(����[�B4zv�FA���=_��5�7{�Dt:�'OH�sU���s�}B`���d�.�S2��=o�ʌuv�[W[�(�e�ӕ�m[�كJv|�V�]o��_?�gް�?���m�_��)���9� � *��:�A�9TC�>D>��67�m^��yhC�hqZ���n�a�Xf���a Z��3�K?��v���x�|���(�+�N�=o����6�)�sښ��y��P�9����Ν���hX�L�D��9:�o%D����*�{n�n��Y�W^��.׬<�y��f{�3�JEf޶괵g"��O?`���]v��U�r(?�����7���y�l��$R����Q�/ ��]7�g?���(�e��.��N۱3����G��7�=�����3b찂���=������|@j�A $�{a*���H�G��������;p�����,DI^Kk.m=��lD<��M׭�O?r�]��[�kc��R�S���O_���΋ڰL���'�P�n�Z_�K�T�SN3a���η�b�����G��Gi������=��+vBr��̿J'������|��m�����+����=����o?�S�ɋ�,��d�ͦ�%��X|��@W�%PF>�5�,l���0���D't���x�� ������fk�v۱cG�������/����9eǎ���\��欽%j�����+m����d�������	�}�=��[���_��G,"e�.`4�a �6j��Iʃ�6ɺ�"y�vߕ��U�7��s�y�2��9�o8}3��$���ƕ��C?=����ŒURcSy��̅1�ŸA�HK
W�f�.�����U�:�q7��f��֦8b��>G_�<_����_�L3B;&8�T��L[V�J�heҶ�_j;���M�c2Co�9b��ɂ%�K��&Z�NFȋDW��0i�o�Ȫ��g>�T�Ӳ,��uؾ��.{����Α�r����
�f�*[�d��~�ݶ��,��mSь��ǟ{�~����W��*���N+���1ɺ@c\òaY����e�f
��Fyu��aʻaq��7/��ǖ,�q��}牟ڷ%�/�9&�bںzHx�}͓y�m�x�"[�r�u/Yd�TZ�({�'��>k��>��tD�O �}�I�d�J��F_+]ƺ��[x��������:[.�ZyC_��#�v�|�E��g��'^�}������w�޸a�<��BǰfsR��)�l�/�O��{�%��[v�숍M!d\�\m����׽�DF��u��1�Ʊ�Np׽钇u�{!BN�;��f��G�M߼u��+�|a����Ǟ��/����ݾa�B��<�f�y��2V3��.��?��^x��9f�%�)#pa�R�O���L�@ 1�V{؋!����;��t%(��~�� r<o�l+�鱊�E��[�H��
�:�8�џ+� ��?F��I�~V���h>oYy;vl�[nXe;6̷�m�>kI�0*�$ �j�����
[$pM%��&-.PX+E���-v��U�୛���n��U��l�
1�GRZy ����!"$�ٷƤ��R�tu�դ����~{BV��g޶����/�o��%�wj�f�)˶�ښ��l�Vw����y������~�%{y�I�)[$٢�׷������ h�S�
ۛ��37v�.?��c�!m8��-�ْ���Ĥ���-{��v�줝�P�?������`^<:�-\`�TR�����q���������#�NKh#-�V�/e�7f�t�KBxB� WO"��~��꽅%pԃ  ��͔�lA_�m޸����Lڋ�챁1�+�-Zjv��W8Mڔ�v�P�'�؏�}���o�g_��Ol�['��P�F��\�9)��g�e#��9-���i�=KV�[Zvh���c��eNg}P�=�8*8f����H�M��y�;w^ d
��޼�*��.)�*QmI;|d�{�����}��?U�N���#��	��:�»��%�3�Q&!�Q���P �ȗ{VQ���%ӕ����ޓV�jL�-�$���W��Dq<��cZ �lt�`��)�l���/~�~��>k����?��'�����w�l��uY�mjbʖH�?���m�҅�:1xjkV����җ���o��������o��k}��X�j���0������L�G��`�2�&�V�r̛�@e���������^����춷
��s��"K �G�Z���}�	�_����������}�i:!��EJҬBK;�UsqjB�ֻj*�=n����ϘB:�Pi�A�rJ`����0TP�cqkI���l��y_oI��Z���.XdrҲs3�ܦ��;&�}��=���i��o�`ϼtL�n�T�U��6W��3.��%�@Y]�q�M!����@z�8%
K��Pr֣�7�ܪ'��k�b�?:�Q��Ղu��to��V���o}���|�v�}J�o�t�[�A�T��0,�Y~bț�sr��W�L�zP.�}�9�$E��Ǭ- 	�Ȓ�i�o�!ꖁ�
��p	c� ��<j�+�њ�(cUk�I
(F�ɟ}Ͼ�wi;_z��N[�8a�Z���Ik�̈��{C�]ӳ,,&H�~��-�鯷�����:5(|C��c�I�Ӑ�_&��h9��j�!q��x' �5@��'\�e��;�I8� s��){�G��l�L[$�a-]-��aIIN�b�L[�5�2���$E����r�`�J[�t��^�ټKl�u�n��~y;�d�\G�=��^���=��Ԕ;<�̺2L
��C�E���:������JRx�e��9dy��f�-U���\o�F@@�x��9��7�i��ۿ��,'w5#�I�:�r9���T���83C̬�̻����B$>�T� R"�����B�|�w�5I�,��8:�euX>o9�|�L�m�����<�����ډ�,3��\�@S�j�I�g�]�L�F�b	%�r�#Wil?G�m~wTB����̘��Lҝ&)�IE�\o��1��k���e���G��޷l���ml肥�VR�3z�f��+;g�H����ْT�:c�#�x�P�6h,�"N����T�z�裶�Me�w�׈#��Hx�4��OM{�����,.ښ��뵩!��1�A�FGX�Qr��Y&=g{[li_��r�e�3�\5���񂤠�2pT"Й���q5��>윻��+e�s!o���/�B�P��\�B軂��5*�I�"^��u"A��SO�� �	��Je{��vn�l��8�/�MXk�<+ʶ�Wm`R�SM�h)f�ը���l�2g�ODJڿ���\�6��%��eZ�+�I�edei"U����{����g}�z�4��d� 5#4@�E�U�����Q�u�-�[J�4[����A+NMȲG|M+���;�[W�@A
�������E��k��k�W-97m�XYܛ�~ �#Q^�8�b(�%#���Q�%��0階�gC�߷韻����j��	wvv٢ŋ%��f�N[�hoO�YwK�>��l�<�E�;6jN��Yy'}���O�	h�3Q��،�����+�f�M�C8"Ԕi�Aa{c��Fz��*a����}^�V�V���^�A@(��pc�-�Mن�v�M�l��%�&���c�"#�j�:+-��e��/�N�,vMޓh/Q1�a$�el(�{��<���u~�S^��7!�!����)9d\oV����o^���v���b�mikUܲc�=p����!/Y�UK��V-_a��ͳM���7n�U*�UKzm�e�k��y�	�R�����n�yy���S{]�i3����-���ǐO΅��*���A)�xʕ�z�����G��߰j�]�}��@�Uu�!��H��k��9��t�R0y�vzp���~�^�����5_�b�<)�,7��F���Q
}An����2/4gڹ�T�����fJ6��;n�d��}��ufm����k����~�b�4���4'K� 1�R�rYϻ���[������k��׬%�D����v���frb��K�;�|JQ�dx��~�t�K{(yX�xΎ��g��cg/L)�j���ZT�b�Yy�h�ܸ&u��^ď�����. �ߣ y�G���>�m߰���6=2����N��}�$�B���ɱ))�V� k�0u_�12��:q�~���v��@hb�kN z�*�NP�V��_/��!l�؅�� Й?"�,@����ۿ�k�F�$K���[��S�qq*y����S��fZ�����{^�<ѝ��c���=eϾ�[<�Y��2�ă˃ߟ��U���-RN6T�+��G��ʒ�h�>����O��f�����Igm|l�8-/~��o�Bv���Z[[e��7\�I��������3�gϞP�+�S�t�kmm��M��	 J�87� ���'h��/�7��WI^v�㝅pN:�$�/􎁉��_y�n��ߺU�U�3�<�ʜ����4S������ȸ��?}�^x㌇t�����y�a�(E桀�[(�-T|�AG�+E�?�JI3Ɋmݴܺ䍼���vq@nn��ʊ�g�,c��Gȩ�> �9W����<x ��i�y�f�������M "a�������  d�e�}�s���l�[+эp�f�m�����۳��%��^��2C�֨T�^�T���}���Ae�Hn!�[#��T[Kܾ����CT4�;)��t3��XP�U�JU<:��T�H�
��r�������)��\����������P�<��@�HXt
������Tߑ<t�J`��W/s��;�$M���B���mv�7��9�P8�8���3�c�XN�(�\�f+��$}��)�d=���ny)����'��W��+��M�H��mW�J�л��"}�PU��U^�X)��O@N�_OW�m߲�V�s�ꤣ✔]\ ��3F�{;�-�
a4�Ң�����J�{�=��.;}���/~��뻤�����l�R N~.A�Z�#��W�F ��Gh��J��G�?��;�]j� ���"R&����X�dUe���������'��8�D�~0#�< �"aNGj���:��aA(�cѣ�g�V�GE��5B�� u�Ƽ#��yG[�P�s����mE�"�!�Q����u�<�V�h�>�U�'m�ʥ�[��E[��W^�hd�T.@A�G�� XG�bz�����m�Gqay�������I;}nLy���Tޚ�g�f+3��S#
HPD~��;� _�+?�U��d�ݸ�>r�m�۞ �}%��<A�L8@��]"AV�܉h�֬*��P,���i�ˣ����;���S^�23Ǹ¤�z媓B�_����᫃���d�IyE�;�}X��e�m�,xV����� 
F&�<��P����O��O	�B�|�:i1�Ze2#𙓯����AD^4���a*S�W�A����($km��By~S
�E��@��J<>�E�(@�;�+��{�Ɖ�af�RA4ÿ�u_����{���\�������]%s)y����'����\	e)%<�X4@�A��+����b��{�+��-#� ^��D@C,��I��%�G�\�?��s��ދ;	i���SW�N8�5���y�z}���఍�NKh��L���R>җ�ar�Xs�vi��n�*vg����������S6<%�g�y.��5��lOP�"�p/Ȕ�2�D�ްn���t�`���\��A��I���=���M��',�RR����E;qrP嘖���T�d��>iPS�����TaC����e�v)���6�ŷ�-�3�Q{��3�v��[��υ��y����㙚�H"�f~*���."���k�^�g����CO��@b8nHK��Sz.���yGR �ðy��SyX�l`	y�E��	d����Y�RD�$��T�Nݏ�Ȥ�̂�L�L�&��e���o� aD1�K���L�-�{�[����0}&���Y���u	h�� �@n�/��5�Y_�E{�+~�g�śtu b�9��H����"��K�t�=F�S�ܛNS9wD�ˏ�w�@��m�܄2W�	�&� s�D������Ȩ�9x���oھc�Ōr���5�h�Xw6m=��u�l��u�f�J��������'����6���T<�B��즙��\�о��G��˙"�"���+69U�'�y�~���6\P��R��Xcw�f�RF.�`�-3L�:�yE@�7�i�VOC��8���e���C (l\M�䔰$�1�hA�O��f��F̲�6�|܉s�&�r	0�� "A�C)�zR�o�yD�h�n5�)-ٜ<����>b�'��ct�"��
���y���0"�,��^�x����t;d��	v��/^J� �Ы�;��[J�:}:&�)�Oԛ0�FI�*��ug��{y/uP4o{����E�'t�|��BI3��<����ˁ �s�<4�"x7��%�Z���e`e�s�8}T��Y=�����<E~�}���]���i�<���<xcx!.�zBn�/�&l�fG@=s�+��+^���@�����y 4�>S<i���{���o=`��S$��V�\o�	�^U����I�.���]��G/��XQ���ȍ�hM؍[�
��R�~��ؼƭfJqSG[ֶlXk�o��Lϟ:)�*Q̬)�)0�,[bw�}�bHZE��x�K��]�z��r��Y�7�d"���Ӊл&�M`E�*4bV��Ҙt�g�sZxX,��@���c�&iy&̩J?Yr=�t�>�Y��P��I�D%��9 �
	l$l��w�RA�/@Hݲpx��ʄ�<�&j�0f]+Y��d,8Mx�jx,�A��hвh�`=�W�qϨ�����>�Kލ/����5��8� Ky� 醕!����>R�<�uz�
{����Q8C����K���J���jԍ)�TYQ?EȜʝ	�����@�g�<�[�1֛#��3�6y�[���H����$���tW�Tphw#Q� Ө�I[�	�bI�9���3Α�<E!���1r@}�1pT��
��/ �_�]�|����~�o.WWO�G���}Prc�6 ����� �ć0�w��d�Q��G�� �$��F���N�}΋!eY�����O�е2e�V/���/��U��fc�e���peEXB�*˹n�J��h�JaB�͸M�v�,--y)�s�roUP�&�s�~�W[��$[��Cǭ��s� ���ƞ$�!Z��SxU ֗�-Pìm��)&P)�;�h\&���4w�A�G�����J������'��x����E������¨�p�w\.p�QG��P�&���u�+P�%"R")>9�ޫ}œ����f�N�YX��^��~��2a�r�9)15���\��/}Wh�6�{�|C����Kw�mh�&j�|/��JM�S�gQ��h&FI�h@"�uxU��B�fؠ!��������9��<xG]y�S+�P�����KD,�A�������4��r➩_��o�� �xd���[�m��hs !��H�,�WI�w\uӿ�r����zw�Q~*������[�{6	@�gE�!��$��ZZ0�8	e�%k��6�c���7���f��垊����KZ1�j�l�M�$l�P��\��������}�ٚy��6[���Mڛo�m��ߴ��ߴ�Z��Z�@,Ax!�cy�DH�C�C�ρ$ ���%6�:	�(P���@E��{,7���a��ʹ�`��ޅ��נ��:O~a�_+y��~ϻoDu R�>�D/��y=��{8n��^J���6l:�7���w}��N+?� �����Lz}�����������>�J�R^��n�Gd��;7��.��֋�;����4@��	��Q�J���t[Ȅ?��~��B	]~�շ��w���>��:�(��A�)5��
��l�5��m�M\�����n޾�j�I=:gE���w���=�Ӿ���γoُ�8b'GK6!�(�"t�v�}w�d_|�>�>��Z��K%,���pގ����}��.Qq?} ���Q� R�5ćd��wE��A�\�]��
�ke�����q�M?�w�{�&
����Y0��/5����rtM�a��Ľ�J��.?��S���!�}Cy|�=�,�؜�@�U�frͪ�YM%���@kJ܊��N�[~�%�s��W?=�=��;���^�ت����Ȫ�S���B���5�}�m�E����#�C����߻6��ѯ��K����J�=F�P����x`B����+:��V�7�~���o"�}���y?�Zc����Ixqx�����/y�ˎ�d�R�H�J���ST��u��u{���.����0��%�@����/�f�{�y{����i;r�8t�gD�%U��
��z��#����~��?煕K��<5n�V-�-�Y�V�Y���U{s�!��0Q�ȼ�꿴s���<#AeB1�K$٨�`��^�5��gK��C1��3(��;'=���u�i�Fr�J��3��+�踗�}^e(��4����^��f��f#����+S�T:B�a�^v�X�\;+�3P�ȋ?��n������PH�B7��q��Bt�+��t�B���>�����u�^�;u�s��~^�W��6k�Q�:h�C�.�/��W�k�`ǥ=�����tI�~Ѥ��w��5o=��P9��FuE�;�v1�IWK�n�i��dC_-�Z�'ޗ(��/d�c7=C%�uv�ZwW��^P{�ʛ{�?���:7��#��6ecc3�?T���ۿ����?��w���'�@�I���7�>��ݼq��4M[�:a�?�8>h�
q��!��dI�j�QEP���,��_ڠ[�����O�<��-�<�4l����F7��tb�K֊c���b��H�pX����D��q ��-������y�O����sB�a����^�ӱ�)潾�n�3�f�@o�M�\a�>(�m��@�Y�������C�-���C��96WQm��:&B��y���K�?(]��{�ڜ�����[��-��7�� �{����/��R�{9]�:m��}���e
<uK�(�n�aᇦ� y;�������P��7i�����{�<���9���k�$,V��Z���b�^y��ŷ�gv�|"c��h��;쓟{�֭af�I��E�81`Ã�X�� ��3*�����7 ���zR
��L�ַ��'u����������Vk�PT6�&��ػ`_�T?}��<l����r��Kms�)���y���m*K�.lM:f�Ĺ���&|��Nj?�}^[I�н����N<t6�)(�{邳���N�����s�����z�B� �p�d�x��-+܊k��`�E�ɷ�>���~�
1��V��al	_�`��̳Q���@�	�g�O���Q� ���[��ķ���U���o����U���E���.ᒧw��_��W+O��r��gj��M������s�5g�dܲ2����$L�J�|zy�B�T�B5j�Ύ�w~��=��vN@3�/�۴�~�W��vl��Ԭu�&�K�NGg����������y9��6!»*���%�/o^�TrK#��C�u���m%�X�Ʀ��
���Y	�2��;���A�0?��_m��.�ب�	G:���'݌��H{���HAg�*��pWX�H�|�� ����Y��>f�?��90����)���n�ߵ���^�c"����ػJ�Fl}�|*};&�`*���g\=����w��:S���*{�<����=u���ɯB���FMI_B���H�Eqj��(������ �⺶mWm���/m�~�vՓ���H��	oS鴥X�қ�u��H��%�o:�H1b��WQ�cB�T�r��60Y�����R�'�>�-.��ټ���7b�҄1`,NG�Z�.�����S��7��\ZV�ٮ߲ž��G�{o��[�X[G�*e+�B�_L&��RQ��3��Uu\]�I��)�����Ǫ*�^Y
��	��$��T&nF1�JG�!SV|Ϥ¾�V?�کXyF�
 ᜾7+�d��H2�M�4Y*�&�Y��-4�66)�D���I{X`J��R����_,E�6��<#K�J��TX�{ѯoFya��Yn�)':�*씮��Q�;RQ!��*+g"���< Yk�G*�WE"0# �	��A�n�k�9�ӏ����>��b�����J���Xͻ��7hڒ<���N*��M�U�|}�����V��� J��U^M�5���^�@F��t�g�ױ��<�9�Ug�[��$7�^�Ɏ*���DE/�PT^�,��w�r��7I>j3E���o�DT��ԬZA��XV�M[$J�C�F>����wk���Úh���p�A����^+/<#����T���6B�F���ԟ��]�Bhn�~��X�lFrI���a�������"�vd,��j��Q��/V��G�ȉ~���W$}�:��{2JwުO��h^��]�Ȗ,�a_�E�n�dLބ<��b���?��"n�z��c[kζ\�I\��dŒ�.����;�?j�0H�Po�UFɰ���`����  ��I��<�\�&�a-)<r�ku/�-�&0] �k0_����\Ǎ�a�)�~��O����5%}|9F������T����A@�g #`�䛞���l�U���~5��)z�̣��}b ��+ɥ�G^8�{��y�L���v�E��)OIr��4�M�M) k�4Zg���qL��%��I -��
Y1�)��Y}0�v�����7�PB��iџ@�~P���ݍ����X�~{g1!����xPv���{X��3�T��iO��,�o��� ��y��}*�C}Kߛ��p�}��� �!?d�������ҥ�/����;��?�J>��W\%���E}v�-��ʯ2�}�tϻz�6�R` �%�v��^{�9?fLx<8h����[8��vl[k7nYj�7.��o�h�l�l]���9vJ A�q�K�Og-)������3��}������I	�2W.X��-#�_�0dϿ��O���u�p�:�(H��#9�t4P�P�,&�)4ӻ��3�U�@��lJ�i�:���_�A0x��?��
Q �KRj�����lФ� ��
g��}�p/��K�I����p�U܁B��y Ga�l��<e���%yw!@jnR�K�2�Q��)��|Zȓ�	$�/y^�qm6�w!@�!M�̯B�ǚ�~L����˃Rٲ���Y����Mʫ��
�X�,=[�T%oIy�фX������f'���8n Q�,:�-���������yI>����*ɋ�����$�s�y x:��..#��Q񷊗`DYzn't�q7�/���S��5��Ը�����K�_:�?DD�x�g��"m9�G��������G9qwj61����ڞwNY���Y�)��'O�[[{�uuuY����e[Z�(�i�S�7��ϾfcS����t^ ���+IW�\,���36!o���ך;�,��+rܕ���d�^}�*ƀ��-�m��B!�=l��Ȩ+F \PF��ܹBѳ0l��R�����J�P��'��{,�
"�v0�ΉD�B�ax.0�� �Dﮯ<���iY>?R5lb�R�+r�h}Cw��Z���t\�s(��z��<�XGG��pA�U�&�ݔ�:�Wh����@+�f�����J\��P�y���uψB�X)oY�L\�*!]ܣ�\���QT-)Z�:i�
3�f�7���֔�B=}�e�/�)� � ��O�q@�
�(��MR�ư�a&.oJ����ҧE�=�&t����.ʒ�/��ݴee�X(mN�=K�)E�$�QA�����A�Aw�{95Γ.�����+����<-�yI_��q�zy"Wg+��>����I���s�ȱ!.xH�x�B%��ލ=ےS�=�k���Zq.i/���v���ʳ�\��d�Rj9��5[#V����X��x}de@�%�K5����=��^�3.�֔�rҼP��@{]a4Ȥ6��h�3]vńF�1��
2��
�����r�[D$� ��8��y�����������V�%<׸�d V�H(�	�xt���(��m*�$\�w%��\6��0XJ��CfT
�x����r�I4O�B�7��5y�E�p� Ш�$�N$�M��-h�ڍ�V��=���Ͷ,_d��w��\��gm��^��b�
s��,a�rT.K!� "@ݿ����f�}�:�e�F۶j��t�&[�f�r=k�CÒ�4��RH*��ަ���Տ�K��7�H�-g�s�� s�)���s�0���0�15Yy̕% �9���lK���g��%�pN%�<B�ws��=\���f]�FV�9=�'���?,]���q��s��ȼ.��f�H�"2��|g�("։��4��B�84j{���d����9��U+�I�tF�������6���֮]k˖-�����7��1;wqԽ�)y!�-�659�/��))q�f���"�io���lӆUv�M�X2�����}�{O��d^�d��"UB/� ���3�� 8���qd�<�,�8�ݖ2z(�]������xŕ
�R� E���Y�yi�E 䚣�z����/y8zJ׼iS{o6��	!
	!�G8�Gm����
��D���a���!�.� EB^�@a,iis����"ӥ�@�E����}���9B
yv���,t5巪�yk�̞G�Rٸ<�?}��6���߼�>q���Ӓ��,+��5�+�S�15񌽶����c?�SCӒ�v�&�36e7(�����Dºj�RyNI�)�Y�E�����߶�����t?�n����l.k�´�ސB�S��k]9��᎐@)\g3�a�<=j��!Y�v[�t�)r��|ъ.fh������Ԉm۸ڶmYo�V.��ִʉfv��
��yy������$��"�D�o0h�����_�+�i���^�%G�2�r��}P�t?[��$�KX̀B��=�Z�z�&�����޾u��w��Ӷ���^���{"�  �7u��P�٠�����0)-X�J<g�640l��Łq{�#��w��mF�M�KJ�D7���VJ��zsQ���K��ڪ���;{��8m�>��s�^|u��L�;�/sR�HHO @���uÙ����9�4���" Y\� ����{ƸFyy�n��/��Nh�~�:��w�n���[g���!Տ�;l�K-~�PpZu:k׮���}�ݻu��]�ЮߴN�Z[.�lA�mۼ���OOkO'�k�W��#k9Z=�߇���Q�%����ˤD=�B�xt�9]���O�,ۜ�� �d4/�u�K1s��u�@�w5[K[Ύ�9g���K��/�YR���w�l�|�N��2��'���,�$@��Ygw��={�<��QXcf1ʞ0��)苼<���%k�6d�Jg�]��,*�	�m��g��~�ч}*�Ç��d�Ų� Z�+�-��W��	�We�xa���tZg{NF0c�׬�/�;)h�+p�DW��Q{9�z���/�am�����?,]���q��{?�Q�����pF�A��xO8��� ��tv�.ډӣv��J^�1c��&+MZb�h]�e���'mjx������S��\ޕ��� �]M�!�������J)��Z��|!��gN��c�f&'��ae��)���AP_A�8�^H�i�=>��Čk�R��I��~3�IsJ��䨥��ã�2��M�X@/rXH�=(�	�3aќ�-MY[6)�v�XS<V8�#�Ϲ��uE���CL�X[�1>���}�!��/�d[6��M�7ۆ�m��c��u�Y�r��m�v��!yv��
�nܺ���>e9yV�O��'$��ю˒�E�ӣ�|�֭YjǏ��bu�GDa�6��5�Q��A�ǆ��bJA�٫��خ����w�2;���b�z�R���ʼ�|s��ײ`'�W��n�����X��A����i���������:�?v�:+�SY&�Y��)Z[���d���{)�ҥ��r(���H�oܾ�>/>�]�i��%{c�^�"����s�c�
���+�f�2Y��I>Ǌ���%�欍�N�K�Fb�f:�����C�����B��.;]z�< �sL�������G�7�/q�{@�ן�?�HCƜ�\ox&<Y�3��L�h+��=����|lg�������r/gl�T�h�#�v����u�����>�Q�놭�a�B{��[�;nSܘ�s�/��_�{0�j�S���`�d2�2Y�����#�[�*,j�ѡ~y7L�(���$6R��� 42� ߜj6E&��U�C�Z����lV�Y����ﴯ:O��T4�K.��ͤ�**Ӳ�^e\VT��N%�=qD��*!����y"5`�<�%ZB�B�β���F���/��2=��F��0�ތMLLX���
��,��o�3��r�,��c��i��۷ؽw\okV̳�z�����'�o�\�u�ۣ���.`9�vap�*�
7$��N?��a���+��&Q��|�,1]�لB�x��
��X� ��Z����;qfȊ�}��G_���^�c�}���׿���<;j��}�`�W.���N��o{����"�,E4Q�WO��L7������2.�))���W��7l6���97`�������2N��e�2��?e��/WID�'/�m��;?�Ǟ�i��\�Bz���ɳ��K��>�3
����%B��d]������-�`���Z�U>��x���o�~��y���$?��{׭k/�oF��k����N1I�X,����t[����(��ي}���/|�>��g���~�6�i�:۰v�w�W�$+N����YyT#��H<i�XƦ*R��f�z�V�����#��W����?��m�r��F���{��b-o���Q0!/��q��:#�T{���)M��l~W�n�n���o~���?�{����c������T�1	j�Z�M�����햛�+�R8&KU��T+ؼ�f[ ��V/�% h` ��qHЩ�
 !�
՚<���k���Oط~��o_����o|���{?�o<���~�t=/�� ���m�VR�^�QyG���sQ��|��V��ԊYZ�T�]�3�#�&��)E)X@		�����+����|o�^� �k�	.�ܧUp�Y�Q���6��Z��uYl&g-1m����s����ğ[�m�g�����6&/��������Z��Od�K\��r>p3�M��&9t~�r��ë�8Ͷa��&yE%y�
'� ��20 �.*�5ۦ��;6YE�|��Q���؏��o/�`O������M�Iǌ0u�8�M�+�/e�8�F���˄論����a�}� ����{ӵ���ɟ�?�J�
[ �p��	�J���h�Gcn o⢥3I���f1E�1[1��浵����/855�W��Ǟ{�.�mN�"�S�����RZAX܈B�6����ß=g;�9k3V�`�x����=l7o[%�?%�r�1T$:�@���}�f<j�CA��i)RL�Z��v����_�����G>r�mݺ�>��#����%�O�ךR(V�d\VIBzÍ���Η�W?���Y�]�<*r�˲Vk��֗���K�u�j�P�p�͸��]�%	"�u��JF<�U�� ���D��?e?~��ۯߞ{�+�}&̊����IkN�,�(Լ`�N��MW*tX�r�p~Z���Ls�p��L��J�)}�%R}S���V���v
{��]{�U%d՚ Mߍ���ɻ�S����.�V4���R��j���M:e�������u
��z���GP/�|J�}���e~�D��
#�S���ӑ�p��Sw4K�d��S������kN���T�2m�>��T>�g�/(]C	�<�bh���D�+R�M6V�ͥ01�|��$N5�����k�׷p��;��r
]Cb�}څD�4�ҳ�9ER֙��p/�'k�m��������ڋd1�-6�j�Β�8�b����uLp^B[���u����o?f����s�A;;:h��V~�ч��m��E^}$�U����L�'Ӵ�U����3k�|��[����%=66����b�c�,��<�Q��F�{Q�ϳR�HՖ�\l[�-�[n[o�6���'��֜j���m�{�q�V[�|���@�v"U�� W	/�G"�_�;*�%����IYKT�ܲV�����E��\S��&Fe�+���:yQ��~U�p�|{��l��vĔ���M�H��r���R
Ѩ���²PVR`��h���)�7��Qc���}\�1�2U� y�sY
���h�V����3���Q�-x��TԎ��g_|�&�i�����U*�G+=K��^Hl��/���0�*�Cg¤ ����r��*���s�1S7�
D����#��mJǾ���J&����!Q�y��-9� F}��eO��<؇����}w��Q�����I���4���t9z��I~��hq)��.6�)^�? +�l�R[�p�'�J��쩟�a��Oځ��>A}/��ƥr���S��;��B�������f�ݧ�?x������-�p�4k�֮���u��er�([�$�ӻ�0�	%u�)" X��Qy�y�j[�t���v��}����?��N{���G:�k�"���EW�抢SVp�;m���V��lͦu�lQ�0A�ԥ��C�-L��T�!���ᤐQ�CQ�M�\���*��$!7# �iA�c����%��GEߊJ�-	='���P��b����<yn؅��[���7{��9F���3�Y0��KE�հ,�A_ɡB�Z��.č�{������G�<b�l�<�lR�*�a���MY&���QBn{�����]��~&d8��I����X�Y�Px�S���ل�ވ���̿1o^2R(�*��e�2Jɝ��h��@��7�ؑC'���Q���orE�AҌHn�Q���t>#���^'����PWDm\�ԥ����0� 	a���@�\����� qԠ� BB(�_���j!ҧD�g������Y圬M�^}�=��svaD̏fee$ܳU=;ms�������V $-c��͚B��ME��ԭ6]Lر3c��K���reϟg=|���kQ�g!����i����A��LAG{��_��y��io��d�~����;��tȾ��˶��y�V��"޼�K���e;u�����n;?Q��7�M;�Xw{V^��|�%�7��5�j�~��!�:�������)(,��mh�D@�b�W P�N�OJ�XmM�P �,JeD5y�m��|��B�6=]���V[�l�<�	�l�i�n$O�i�%V�0pa׊�=��AɅ�@.�nyO�X��.��_�ă�{��9��Gﴎf��� �n��T�ǌ�-�,e2D65U�������%y*E�_0'e/�Zs��������PW����ЃT`!Y, �)7&��7�k��"�A�D��'�I���/"p�/NA�� Q1��Gh��c7:��}?=W&� RWVx�C�N��l�+��}��}���kÃHx�!�n�˹D�x8\��Y�0�9�sD9k=�i�&��7����]�ڐB=#o@�&2�P��yQ��٪��<+X�����@gaV �)<��%0g���������I�I.c9Y	��Y3敠> ���~�X� �$CLPKȚ���u��(��*��v��h/�:b�%�G�~��a����ʀ�m޼yv��wɶ�Zs"e����sچ�>$�v�m7ڒ�m����R>z��ʠ�"�'�s���X.��	���m���PZ��_@�AhR)Q�����ݴ��ܶ�:$�RAo�XB^RY�\��g�f�����ٴ�{˚e�럺߶-n�[�.�N�aLޜiWY
	%(,@�1R�b�9����_#Aoc#�=#�1�b���rv˽�/���v��7Z��)n�U�9-囑��lj�:N�ľE2H�V�q'� ���(��-?Z���q+��gB�!�8��Td��)o�օ��tߥə�1[?�P���t��3z'癍ݗѓ�'��N�`Aԇ"��4��>�Y����Y��6�����YE<-)�F�9����S ��vz^�ɥ��8U�e�?����`T�G6�Z���X�+�QV�&�z'����1�X � �>J����/[���rޛ���7�LL~Ozڀ�%5�|����Bxi�X��d� y^g*���X�4-@���挵R����(Kz>%�W�-w�er���R���jҽ3�^ZC ���/�mo���~"'�7���o"�e���7��b(L��!H�d�Rxڒ��qZyB�>������x�F���-m��r��^��
��W5�8e�Ik����m�N)����4ٴ�_Qr���}茘�9j���q���6��?጗S�r6�]a��+_�����Tx�$>� I݉��:&��Z��Z����v�b��%��ͷ/~�Q������\�b^�"6�!� OYa͌�QQ�����UjlW�3=?73-\�r��6�PupR7��:��Y-�r$,���w2��.J�fuo��W���SRxh�x_��<�����w[F2èZt�gx���Kۥk��X�	���&����?�?���h��΄���2d4�B����e����WY� -e@��$G�2�<ғ���Boj4O��q�S���=釯��oP�⣰�I�p\�G�2����|1y�Z�=,@C{�p�֯���-!5�ٸ���*6���~�r���$ݍы������Р,��&ѳZb�ri��t��Ƞ�T(ċQc��f	WZ��G�$׹�«*4��D���Ȉ�=)�[�Œ�3�FL2�� �g�6o����K��`.bCG��@@e0��d���	圦b)�����X���s�楶a�R�J �V�O�.yYg%�����e)��UK�\�PTz��=�9�Q9I��F+?��WKw&���n��n��3o�e�.3�9	wD�OZg�	�TV.�{o�a�ηY�D�t���Mg�M���sMֶ���j��lS^� !|L>�A� ��g�qy_IyLqY��w�f�i��'�{?{��M뻱�M�,��6gf�d,&��;����Xo�|�~�{�������Y�ZѼ,�����$�pÑ���`y�_=%���.���U �Th���% L��B�3��
%oD�Raȸ�t�ٿV.N�#���3P�&Y.�o��L�ݤ0=��,!Ħ�;�y��~z���0��A�]-ɓ  �û���S�@���!�i��(�Dg<�A���eƁ�e �v�[�G���H����ҭ�`e!��@g*���?��8wֺ�,�[o�ɖ�uZW�j}2.�����.����\K�])оI.�,MV���Bꔕm6?l��������i�Z���V2��W$�0��t(�|p��wIq�m���3;���D������*((M�[����h��2�Z�ù�R�z�/�u6I�S)�^��]ȇ����pN��]�����ꇞ.�C���B�c���A�g�<��"uT�'.+�+��"��?��>ve���ޑ���/��LFe�I�5aݝ�?���Jɷ <41�`5 �q|�^�O\|��$H��^��_x�����׾��8qц��e: A�Qh[��oѰr�j���֢|���=j��9y)rM�&&� )�T��x��k'���S��Z���pM(1/-��� H ���/��6�p
Z��qv^�{��M�_���#q��"��&D�x,�0�bU�9(��Ë��r�-�2����7��1,x"��~O]�E���?��P�=�+Ao�y΅���(�o���6�	�hR��m|�C'��K6{Dy��e>:0l���~�v�򣟴�n�fK�▪�J�-N�]qҢ�E�4'�O�S)����OY�<i��|�i[1/c�߱�>z߭�6	K������~H�	�V8`82� ���M���+çܪ`R1)�P'��4��D3����#�C�ƵK�;���N�Mm)�a�U��%p%��K��j��W����S �<w�7]�'J3��ۇ�O�����juFa]�
sNn���+�90֭\f;6��Y���?{վ��'�/������~�dD3��<O��$�WF	^���	]�̌�����L�f��h�4��H���I;tꂼP@s�r-L܃'����.𥳐/��P>#��E����"iK��ָ�#(���C���se���[��q6B��[�������qL���½3�ɉis�ܱ}����TV� (��G�k�lb���F�W�eXAU�6��f#�Yn��%B�4:F"�J0	�np�6���r���}�ox���&8# .�������H�m���A$���M\�Z>[�>^�f���]�ցs�li��n��>�ۗ~���}���;�ٍ{m��۾��6-i��q[����I۲8k7�鵛7,�;�_iݳ�>����K����n������셝o���$T(�)01l!��Ӎ��f.+gR�Y��9'�&.�MKT���H0�t�	��-�δX�\����x�A۴v�,g����gv�cO
�r
b6�b�P|��2;��!\�⿹z�v����c����(�w��~��^{���6]i���j�R٪���J���Y�+fc#���<a?����w������O�h����M����lxP�{��U�%�G�B��(�FohZ���	�Hi�W-
���kі��<w\�����5�	P�E�ũ�C60Y0e���s֑��-65d)��-�^�X��t�pJ
�jM9T�Iߠ�[n�%�o���wz�Rm D��Kx�I��qI^PE<��bZ�ǩ*C�S.��_�®߸��rE��-33��L���x����

����])��͍
�=��I�n���Wh�F*�8�MϞ�:x�w�K�8l�n>H
�B� 4�@�m��� "~���s�ߢ��v9"��H�{s�q{�ɝ���r������q�j�������w~�c��_y����}���<j���G���k_����_���������W>k�����_���춛7ZWgZ��o�CxV��ҫ{�(���X�שw&\���]p�x� R!���\�,�,LJ�1��[J���Ɏbv�̰<�!��Z��;n��[��ퟱc'N�w����7�o�}��7$ɦ�I��(<�������8���M)<�T?�@B
��_YBY��h֦���/�Fm|���4A�=)o.gm�=߼xᬝ:v�&��,�X[��"��M*��QH�Iʺ���aX�Z�������f�o/m:���$��M���Y��֢p�c�h��c��S�$���1+&J��z��y{i�>����K����f�-�y-[��٪y=֕��3d泤���Zi���L��ti�k$ڂ:꜎�|㺶����M��y]p�':���L�k�����ڇN���g�,��{G���;��)o�ikOV�-+/J@O%,!o�
|Z5`��pe��w��1��x#�9/ٜ�OD���?����س���9��eE�BO9�R�B�"Q�~�R�.�OH�k
"�����YP�D<�L�0�b�����?���>9`���ݏH	ۺ:�������vڪu��ƛ�ڝ��h7\��V�X`]�����j��fk��lg�M��f��v���=���6�W(��#&k@Ů�sD� 4�Or��A���F䎎Oy8S�����\Z!Qiܒ�IY��uf�֢g��o=���8?l��.[�l�%��{�`G�C���d:gO�����uu�X��:%�� \�B.��G�9���A�  g*�V�0�%Aף
�R3��L�3S�䜼��,��SQ9 d,������r�s��`A�%���`Y)[��M���;�$mނ^Kd�$[ޚ��0��
���hnX��n� �����:(ߙ��ݶ~�}�w���G����;��/��}�W����W�V�E����G%z��>sݷ���,�^�]w�v���������?x����lՇ�MʍdA�,�F�ki��˛��6�<�-d�7�(��@��� �>CǨ+�$7Eܬ@�F���<'����[��������mX�ާش��r3#��2k[�/P�i�2��j%Bx�D��	P���P� �(�*�d��_o����uץ{�=�X����.k��2�,��y�6\k�</����/��|x?���}�M�����/8�X��� ��҇���٦��<&J���Lߧ��eZ��f{�#�Wr�_9r�f[z��h��b�9Y=���˝��+���d,!�IoY9��ͤ26!M.��h���˷��o��i{����y
�����ٺ���mdE�cs�9g�a{}�Y)M�z.�{�]��|۪͌Em���y?����{mL�IA��\E* A���t�"/��w�Ꙙ%�-�ӊz>�B��qXuP�^��i�gpS��9�pOE�6����%+���LX�VY���w���I�5E�zo��I�����M[���u�-#��nѻn�|ѝ�� �4�� �Cx�u]�0����A�v��@?V�{�����/<�����j��u�=x���C��C��݈@����e���?Rԣ��쉟�f�F�ֹx��_�ȶ�y������n�Q��۹g��?qƘ�..�����+�6[��+:ri/�i������(���	���)�0<f5�E+��\N����I���[Q��n�Q��>��Oگ|�c�����mݶ�b*���YT8b�&K��l2j�D�%�)���w�^�z��;Wt�W��߾׹w%��O��ස
� Yl D� o��P��u��{���L� 9}�����rHW�'B
'C����ia���t�v�}�N���>�{$��L�g9;uq�v8boPD5MY���b-�VQ�X2k�H�V�o�Q�M�Z�@��hٞz�u�Γ���/���N���च������.��YW^��9O����e%���4:2�}֯�`=]q��k�
�
����ح���K������<+��"aO���kl��>�yzb�Ξ����@+\I��� `{k�ۭ<G���7N��=3��
��i�v:'"؜�� �/��"�?^�D�,.�Zgk�nܾ��m^�<(��~��=va�  ����^[�x�����w��e}�f�J[�j��Yk[6��ֶ��d������4T�Q��.��V!�!pWnR@B_�=]�vݎMֱ��J�Rg�<��8�BH	��Q�s�����;64� 8�p��Z6�\8]��x6���X~B�0+ّ�9|����؉s#�i���6���B���ph(�Q�����
����!O�$C	B���.[�f�������I_����s܋W���E�ť�w��۰��\a�lֆ���ۇ��=G,���:��g���T@�D�F�
��V�\����P�%}�<��j�TH����P���>x�$.�zV��¾v��Ƶ�,�лK⡑=�GB���%X��M�92Y���O��[Fܦ�R��i`M�"�1){�f���])k�e������;� X����qY��C��:eo����^�(�M'�1�d�2���3"<.ʵ���*Na�qi�l�V���1�T��H���%3M��O�o_��}��U�a��{{�ivA!̿��o؋o�d{�M�v����W?�[�T+���609nKW����K��5����ǯ���h����JRGquFV,��/�����B0��!] B���7�-��Yo�`))KM�~�%k�W.���fU=5U���������hfKV��Gn�l^e�-MʕxpW�|�&�I(�/	|_޽���~��ɋ���)oO�� �	��7q%!��PD�V{s�nޱ�֮]-o5��=99aEyJ����{�>r���;��<��3���;u%�e[�i��Y�H����Y�\���G�ځ�G:���x0��+�V,����%\������gD-M��m�KuF�\7[�t�mX���&
2��m|Z���؄r�`+�/��-�u5�l�@;���v���)����1�蘧�S�J��<'���d|����~֕�j	����$��^H��NdO<�2�m]�a�B �K�D�R��>Kn޺����i[�Wh]��A�2z@�4�� 2K�`e~pl����v�cO�a�Ւ,�
P�$�.����$w�cj���l�-��flzz�2b>��$�>؉�NQ���@�3�`]���Y`B����K�����R`����)�������R@A�>��������l�������w
Ĩ+�{�ԡc����Sϼ�8'�(e��i�<i�y�&�ؽw��Ž&G�JrOK�����V�pz���?���q�Eeu�t.S��{�O��w�<n�G�`%�"ԅ "LND!�����?�q��G6Z���J�@*^�O�T+�GI۽k���?��N�z��+���w�d�Ηg�����ZY�F�*��l3�މ3���'���_�+�������$�(�*Ҫ�P�Ʊˍ�#Tv�a`��$C���ޗY�c����iUr�2�Y���ڤ2�2��O���<�V%#z��8+��{�"iv�.]u���O���d�9�k+�P�ʟ�^��^���$ U�������(��>zX�u��d�>�ɦU0kf�2mS���oZ�Wo3
�'����.Qή�p0���y
WK:�~�o	w�\xRgt�����;�"��ĥ{I~g�<�����9V��$�C(O�P��̱��W�J���"0�����s������C��Z
���lc،����B��:D�j��= �s9��E��GL�{��$B%�A�t\,aA�����h�[2C���ڳ��M��P�7+�uj��P	M��SH��Ks	u�:�r�r��o�r��PO=o��>b�Żu3�O,��+|SW/Yj�����6�a�_ )�˯P(�Ρ�6Z-ɜ�5Ef�!��0�A�
��s�]d B	�!����oڴQ^�*�$C���4�ʖ/,��it�v�k:x�hn��XBߖE�A�E����iI�D m�621�p��>z�
�,�1)��:YY����3
���-��hX@�Χ�O�Rp��A�H�KD�Ձih��>���ʤ�W����޷ӭ���H�5�3	�E��q\���l��T��z��6 B�9z}2-����-<�P�ų�\U�"������juq� �*h��zIPb��H��,!�dɋ��}Ze�D�~Lޕ����N�֒
�f;_��8��in�݃�j�uɌ��e����My�sʷ�H�r�Z8���Sx��?�3��f3.��Eɳ@$"or��%�D>c+�쀈ʓ��� B3�����O�gw��´�A=!��a�2��-�5U	�(*#c4;2s3t��2����XodN���=S��B&���&Q��0�7����GJ@Do�>D@Bْ�R��
�~Қ!����|P�)���%U芉%3		������s����F}LU��;3���sY<'0�ˊ&۔IING:��B<�R��𓿢�<�MY_��Q�0W�hU�b�=g"e�DR
��j

��8n�����'��#�զ�@���JĨ
S
���(��)�d�uˎ����I��MU��Y
O|��0K,D'K��,u��Ro��,%�J�d�b�<�J^���xg���E?�YD@a���%L(_�e �z��0��J��ᣳ
U�U��
���h����ȕ��+*y���� N:Y��rO��2b����/I����aY��)�I������VF!KW��o�G�i��ʷx�H)E�>p/4��K����@+5I6��y�oʡ�Q(=rEr���s�tqx�}�%N�,�6�M>�=!ΔBFBΘ�����gl�<@�����z��� Gol䥾g$iY.����_{��x猬u"BX���ν����E�t��r(I(h:�\wvp�idJ�(�Kұ���j+�=S�йI�0҄�*t)��,�#����3��$)�yF���(��7Wj�}T(�P�?��W��VU=$HO$H�aJ���A�
O�L�!Mrt� Up�Q�},&�L�y�ȅd�U:+������rT`��y�?x���9�n�� �w��2�"~����*@@�z?͘��Ba�@@��k����
ʳ�� �P��K���*��HuX1�M���ŋmɢ��ͤ����v��1�j��
���o�(��{��lQ�H���~<7:|1]�O�$)%�O����e�&Ҟ�@�V� ���)�1w�tH�'&'�e/�ٜ�
�n�Ζ���$���{J.|�&�&T&5�Q�L�+z�����n�uS)
y���k֭�����3�=&�w�zr��0����;J�+�_��2
ł�Rty�@xkz2�Π�_Y�?�$�Z��CN�2�� U�J�(�x�X!_�pT�rU�<_�6ެ�p=/��L&�ǓyE���*���/���>g�:�iM4�D��+��Xy<_�w��o~��}��՚�},IT�*ʆ���| �}H��z8�%�����׿�u���F�@��P(:q�f��m��y���S!��XY��G�2x-+����3Ai��HȦ���C�P
* aʑR��hT~sK�N��cq�X�&����7��� �H�Pؘ�I�� ��=�J�^圢����Ŝ�Ed%�@� �L{��K�G���4�B�BB �QyT�Ԁ���(�I8��BR�HS=�+�#>+�#�|U��\"�E�Z�>���N�>�YJ��bP'�ڜ�������V2�<��c�DY�7<"���50Jy�v��\(W<-Ŧ+��I���1
x��TZ���5e��g�4���k����bK���%)tsK�{-a0��0/�tY�����r�hmk�o6�v/Vye2��up���h���*��GG�y^b~��&�|�#걨_�p�HI>}����A;�zCZ>�[;<_����^99fc5)�d����O"���A�(m� g����>���E./�3�����GIa��ﶬ�/O�Q[ғ�g,��� "~~�.��k���S/�7����,�X=*�}?��Nc����(�X@��;�S?��~��+,�G�v��laW��q��}�V��h�e<ے�|�y!T����d]��d�\��.T"͹⾡�̥=�y����@���,X׋����3�ßB�u���<sr�j����Gy �KAa9��&�S��C�lB`�(|��|.'���QO�˃�/�!J09��Y�A��+ � S��#��Y�T@h��P�n�J��C����:!aa'ǧ��P�U�g ��^G�	)�.��F������X���#�bX`��,�ʴ���1���JJ��(oyS���c�"EY���䁑g�6 �й�$�%�"o����
 ��T�30���w�)x=�����
	� Xd��� �:��<0�Qpy��9/O� M8d0cz�*�+>�	�����_��o�ɡ�ޑpo��{�ɚ��D����`@�	����HQ��`�٩�m]�������O��35|��AD.�T~������C'�;߶�G.(��"L
���(;!�>�'#aҕ �s~����S�y������g�"m)���9��>e�{�~k%>�H�`�
E��
"��#���T橠+B�Д��)<ދ��5�z������A�^��V�j  ~,IDAT	����Rx�m��R�5P�D � �=�ý&۞7/�F��~�|�:�"X*g��8�t/��:�侩d_��@�F������ĵ�E�<(!x�� �h
n�1��� �]����/�s�苼C{"e�5
��J<���U�RiN�E%<�R�)}7��S,4]��:0��3��v ֻ��ޫ�z'<����̜�ub�;��bSb͠����ȃ���2�!�1�-����(&��P����C��YR�B�V|�;�E�����I��$�	��� +tz�7���Mʫ�$2�~G[�����oٞ�u/�4[`ұ]�R^�����u��7L	)���"����������)���� R�u:s������a�ѳoر��V���)�.U� ��Rj�H8���F���D��[�>�����ʄ��?�����}V����²�Ϻ���Zgje�]1g�+&֨��(!�p&CA �}Pl'S�0C9�CB����;�@����N��TzK�ދ����tЧ���KR���`I��q��U
���!��gu��%YgB�I/^\{��J'��w�^:���Z���7}��J4������
t?���a�v���z�� ��Ť�0Z�r���ʡ&υ�hy��B%�蓜���Q��A��E0��t��6�Va�n	��xot˖W���h��>�9@_ @���>�%�И���0�y�Lg���P����E��-T �����Yyl��<%BXf��.��x=�/ڤ���0a�'��B���-�eX(�m�������mѼ^�HN�����C#�_�����uXF���d~����D��_)�	�+��� "q����K���ö|~�2z!#����᱉1��G��c?�iG"SŠ£٦P�vDH�Z�R?� 
ᘓd����Bf/g������3���+Kc�vY�����l~g�f��6=5��K�I��$�U�����:=l�Yz?�#tb�
��7���RL1�w��1%O;KS&4r��O���b�H����(�Gape�#@��b))X��^Ǡr���F<���{�9���{d�9�)(_�S4���.��%އ+�����<f�R��4��:,�W�+���TN�:;��>�	_iJիd���Ƀ�&_��
Rz��R/�߽ц̱�ykڬ9�x5y$��衐��/�sT�C�V�Y�g���"k�<C/J�|�����15I=�@]OR�E)mU�I�	xga�X�/�_�j3v���_p���zGss��tt90�twYg�B*�z�,���s'O��ѱ1KJ!��5�X_W��ų�q�`�H�Nf}�2ֺ�$�h~��v��i4	��%�OL�c?�e�����!z���V���m��O~��SC�|C�~I���mk���~[���:OZ� ��a�04n/���~��n;rfԊ3)+Jf����hy	I��.(����/�[����n=3��L����Kτ{�C�re��k������l^g��*SPj�Kvqt�x#�4AKxS̬&����KIE'���]���ũI���S�0��&ܪ�J�+Z��y־ֈn��^B'*S�O���6%���#�I!7�g��X�愾����n0�E�D���X��{'P֤@	p�@�wxA��yV��P,+�ݶ�F�d�f�<F�ô�����|����!܄�Z�io||D�D� 	1_��`��A���y��o�ӻ4��C�!�Z�łOᘌ�R�F�5.:
L�R��*��L����غe�,�Ix�������R�"^ed�s616ngΜu	bRm�p��d���+74��p�⚷ꄥ�v���^�J��ʫh����ɰ�q:Iߙ�����o#��n��Y�̨�7���꓁w���<��'ģI��={�	*s�kL �+ɪ�
��K��'�^���E{_�˯��6o�����?Ѿ�$�%���O��r'��F�� $�;���ҁAA�t����<���١p����m�@O��g8O���_{۞}u��?>`�������\Ʌ�_�.����M&p��TR2����{C�1���K)<�2���XL�I���-a���c[��ˊC^�}a`Ծ���GN[I/�(/x'��K��9YG�ǻ�@ر�F��-�f3,JF��Xe)N�APE{�1kqpD�2U.�:����U��d�=��z�[��J�o�)��"�JN��
5B �G���uN�R����*p�lmm�V	�N�s!�bI�0. aI,����EYՑ��Z˛��д�3��ު�w2!��������#.>͉��5�P���|2�CA�^������I�p��s�1�$�n���X�ұi��d�"yy��p��E�sɢE��:��<��z{;m�ڕ�);�?nCE��r��L�� �,�o����3�ձ�ɲ*OtĬ�J>-B�G�c���h*��ƽ�V�B`[�O�[ �2����E��@-�K�NZ�R��B�_F�CH��TR&��d8 G�/�N0�[s�H�a�r[�l����%��Ç�
D^�ɒ�>��ӒӢx��*x�x�p�Do��n��@��<E;���`|�HHH^��r,��=Ҏ�S��������˿�[�N��&�jx����e���g������8g�����W�)R���p���h���g�������Y<���� ~r�5~#�����������3Q����)���>��Cc/,EHSt�$lN\�bK���4[�B�V�����*ژ��{*��\�
�oVde��baJ�g*�?�2e�v]���6'K���N���n�@�A��w	7���H K�����^AVz����;#����h��of����[��q	�Ȩ�+ؤ�����ڹ3�l|tL|��ŤD���hU���I�sRl�(�M��nuh��i��~*6E�[xA������I��eݡ�&ޱ1>G/�@)�U�0=1�;K*���#v���0l�C*Gz�JI�D����Es�n������Ş�B��
��q�_�ڄi �&�@�P�Eݽ/�\��y�nD@9�0��4]��4^���deJ���!��S���%,��3����E��Ȑ<���664h��c6��	�0JTV��%C i�(�Yߣ����#�y]dP2�l�z���P�"@V�$�����D��:�{|at��������6偢��,�e�/7�����F/$ԙ5��[ߔ�[�a��E}�v�M��"H2(?�e�CA�9D�Mx��Y�/+?U�3��,�{{;`��T �+D�_��{@���G�c*�jd�׻fe�wu؝�ߤ�B�,/��.�����zfz�z�����
��S�"�q!�%&��f7	JM�S�d�%(l�2�Ѣ4kQI+���&s��%���!�`>N*C�=�#�3��	��D��w	8�&���|-��B�$��
�*��I#ʳ�����89��3"�*�ɚEWD�C{qj���:'�n/k8% �˪�d�gl�0g|���z��{Sc�T���������Ґ9]3��! �����h�0�h��e�Va"k<3�':�?�g��9�I�4S`3n�I�#�V��忤��ȠIIGǆ$wq۲}��X�B��y��abT�S��F��)yC�(���7]��
�$y�k;�O9/���c��� v�h���jq\��3y�ϋ3>�8�j�ʰْ���K�0<� $y��G�	�ҢW�j+���X8^�-�E/T��[>�o�T��vtJ�6��oT��=n�g�2v�!A��s�z�J����6� ��g�Sm��� G�Ȃ���:���XGVߣ�魪
"��Kk���c���,���yeL�����(D�0$�=SJnh�k�5��/`=x�ҧE�2��^g br?�W�bRq)3�������]5֔����Ha
RĲ,/��Ԩ�WA#ص�&G$�����&䖠�M(����)6'O�*�Z���� �&^�;�A@���$��b��aN��y��FAQ�Tc��4��s�hjB` K�}�_^��fn���YJ�?@R�H��V�Մn��;$��"m(qh Х��W~�  ����Z���tK��R,�B�� �=��q����&��p���72WQ<OE�����^e��ib$�ΑL�����������O��>�� �oH��ȉ����2C��u��[�����AYX�c��'��&X:�����9�����Ĥ�kڍGU|��U���JA�(@Q���CR��vّ�
�!���x��L)=�!�x�ԹѤ�]��/������i��4����L(8&C�ցS�=���~��Q#���$�ʨ��GFSz�2�[�t�.y������Ɔ����h��`�-)�~�2�n���7����pF?!dxt�9n��m�@�&�@_�-�LŃ �x.�o`�H~*�*%�?!r��@A\+6�#�{��j�vw�M7n�����û#
9�vQ 2LŪ\���Ŋ�.�;�xF�H#�Q�@3!33ѕ@�&y9{ڟXO���r��[E�r
�b�R��N�fU��t�ch�񘛃E��ڸ��@�&r� �M���L=�<#w7!��uu
#��S	*��U1x!�rD�}D`EIu�5�	 ���\	�����#g����!�4un1���4/�MxE�E&��
fʌJN�����u�L�޻� �w��0XD��%���g�Ц'Ã�â�1��Ͳ��E��� �I�Y<�D%�VdR�D�ѡ�q;{a@
D]K��AO`�X�7O2d_
 ����\<v�B�/@��Ζ���*Cc2b������ GRB�Ό� 0�~*�5Ys:!�#�QF^'2K���k&�W��J ���d FE�Kg��x#����[r�Dz&)˦S6&y~���6�/Uf���R���qO_4���	�B���[��S���H�u A���S}�[,מK؎m�m~w�d�|y���D5.�)T8m��RЉ�M+�g6-<�����>2�Lz��Q�B"<��(((�8${�&̜u���֛6Z[�P�6-�-)�W8#oih(��S�A���Eeͣ�&MXC���6!�Q����"b��qG\��f֊���/�����E�M��Y�$�,II�w)����Ϊ�qI%&�
hDć�x��U�����҈�x�(��Q����(�g$� `�oYv)[w[���ۢy]�r�<[����u�Z�\��͞F�(s\
�+�cf6	]�h�闷�cS����+�2P���w�_���R�Dsaj��Bsz +B�9y*�,�M��D��	)a�
F�nm��b�}�z��5� C�GB'��[?uB�����M�R����X&V��<���h0P<V9 W('�9a�~�':#O�%B*�H�W!�À ���p^����5�MEr�J���n}�Z�-���!E�y����t�okSf2&�!�")pY�d�uvv����ϐ_�S������t�ɖ,�5+��q�`����=Gm�8g�L01�����S��妿ށ�u�*�N�0��#]�8<��,6�K�v��Y�0e(�%T��T�6��>���ct��s5�BԾ�'�ٝo�ޣ�uftJD
�f�Tx*�@\��%���E�7��,��6��z�'��?r��h��rC�oK�Mٚ�]�/��7��=!kB|��G��c?z����ʸ�ڰ��W
��
��ԆWU�)	H�����"�#G�K��}1)@����;v��7w�Y�3�,�`6,b,m
qe�g��L��{�ik�RM��m�J��w�g)beP�y-��(em�U�q�e�#U�;�	_uM��t�ٲ�����=2*��fr\<���jQaM*�B�d#�r�+sv�ܠ?u�&��ꋦ�,jW��:{�˲,Mk�l׆k�f3w�)�=�=#"c�Ȍ
�:+�V�H�hx�PK-AWK�j	��x�BH�BK� u����ꪜǘ�#�'37�y�6�|����{FEf�8���g�g���װ�ާfAbN;��Yؽ��X�0
_?�}rl<���瞋�e��i�mn��2�f�ơ���!�f".#ُ����Q��T}{���5-���ÀH}��>;���5L�u誒鎕�-�f��`���-�$9��E�O�I�;��T|A���ݒC\s��(Tڶ��A�ܖC_��]0����e��4}�܃�+1��(���E|(�b�>��ڸ�ΖN��!�j=9��6��ګ�G����"W7��6o J��>̣��}�(�o|����?|e���~r�a���Ǐb��J@6TL��[�q��l��rQ8�������"����|�B�2��8��X֊�9I(2]��>��#|����������G?<�M��JK�u3W���#|�&��$���b��>�ŕf&�9��-�s��R ���s�"��V,����.>���p��;�$�	1�I�"�@��{����*L�������ݏ�v<z���n�bޣ�:�]�
�iw���6�ǭ���_3���W������1<��X�G�o�dC�_��n܌ׯ��~���h�M�Lt���t�!�['���aP�E5�����aN�W�8inO-��
�}����V1���C���}�v|��߈��_Dk���`�}\�3,"��"��%F&���m�z5��딧���D��2�1���#Z*f�ʔj�zc ~B�t�"�K1�0��[����H_v~F�](��vG��QC.\��A��%41�5���P����kht���K_:��� @9u+e<g�:z��PŴt���'<ǵP�%A�QC�_MwKsz�u�&H2���&[�[ 7�y%�N�@ڢ02�q��h�y$}��r&�u;�2��11����6��P� `t����?4}C��K��Y��~iދ2Vf5�m�9Nş�p 饾�����\�"����~����M����Ae�T2��T��&cx��eN�ˁ��2�� 	V#�,��� �'������H\�<_�>��ny��<>qg�c�,E��~���T�/���F,�V �����
�K�Y]��,�����ʓH�W�Z�\,e���4�x(�r�r�q��##ů�x+}FMF#�.����&�`<����D9�� ��n��%��ͯ�׾�F<�F5q�Ŝ]��0eA�23еT:������ׯ_e�Ly��Yh���@t F����"��!A�q���yd��@�
�;��J-}蒈�X+�pX*��������fܺu+&&��>��)0���oY�;�r�;�&�}�Eg>3B�7bwa||��'F�dF�j���%�^f���&" ��rvt/��ub�b�m���Pw'�i���g@:��>�G ���a��D�-Ly}��s�?0~9��m��yIO�B:�v����l�$�)����!��B��U`�������ASW's1$��Ba��#X�-��\+@���m�̻q�@sk���Y���#��:���Lm����^t\Z�=5��9�-�Z��ut�V�?���s0��)WW/]���i��X]Y�����m �H���%�S�2�@�V,�\���u���v���'`���(�\���f�(\�#hu �=1\Ǖ�_^�1� ��Bjj�6Qx3;7	cԞJ�D#�@�ph�S�,]�%3�e�J�e�<{�U�s��Ry��D�35{h?7ayu5�0�_��Ǳ����Y�К�5�Z�e��׾�ݿ/~�5:~��-�ZT��P	��Ro�>���Ǐ31�5&d��|���?�V�������xd�J^-��}�2k�fة�1sUp7�"�#�{�e�;0@���=^y�����/��rLM	 �d�%�Ӕ?�i��bj��9��Soڑ����x�p�f��җ�+��מ�ݵ�pwh8�%�Pσ���\�g�� `y4Q"hp���Α�\�&4wM��v�C�a��������Z4�Ї~5������;b�lW��O�� uuhh�pE���!���lujf2FF)TZL�3I-�,�0�������L�aף���O����e;b��29������]�ֱ���&bdx�zd�������.��2�%�؇�ъq�N� ��]_�|'<��-`��=�;gv���o������n��"�[G+ W�7iMY��O�Si�KX� c��YGe�Nж\$��9�̺�^�p�T�a��|"�HE�Njm�"�F�:��[r=
`�@��W.g�l5t���9��l��b���n	2��<g}���T\X�k-ߠ��y��cttE�D��eںV��P��l܎��믾������Y�����3�/H(�NyvB���t�W�7+p�]Pq�aui%����ΩXG�n޾����`�^n+�kܻ�9��/&�� ���jE�Ӆ�͊؍i�	S[w5�돾��� �ŋi{3'�	���2�������0 ;��uu99����P������4�W㝘�k�f�����F�ʻ}EђOb�Z�!`��;���E��y�V�	|j�
u�E�vt"���z
[[��<{ ����e܁阺0W�]��_��Ux5fp�qm�''�a]k:��XX�,�A�]��p�bL_�NF���`u�_@�?l�mA%Qף%���#?Np^�Oպ
���P���'8��k�M$(���r� h=+l�*Hc���l����5T��Q�AS�pzcq
���*<��&
�*�=�G@y�I�j��ף��k#����,�$p��1V���=�$A��7�	�����S�X�r��e2^�b�B�9��Gg��{k�;b��"��I�6�3&�����]qqRY
7V�0�,�B���	�~���اw���F�[ͫ������_}�맃:bS�_��Ǉ|b���\�e����_�����Qz��:ei���0�S�\y�C�f/z�u �
4�4#�0�u0h,�l���~�@��fW���� 5.�k�� �>��fr:�DfX����棼������! U�~�>�����-�-wA܅�@J�r���F]�� ��GaW8�heu1v���<s�%�l��X����#2�&������0�^�V A=���2��o��/��:�Ғ�r�*�L�z�:�8�չ�!Mh�bچ���[������������2q5~�Kc�9<t��Z��.�Q}y' ��Uֱ�n� ���\��m���ך����w`!eLG%�$?3�ͥ2�3<<��`n�8�f���6�z  t���R�V�9s��L��r��/ݼ�n<]#ְ�����r���*
Ze9��)�a��k���+<��[,*UI&}��U<�*�W�W:��A,�ax��k�\niu�څx���耾�A��/��t,�(�|�։f���0�
�扥!/r��t�??=���=v��3]���^WFk�ԯ�*D�3��_��7��I2uZ��h8�/�t#��N�6�����:�n� x���o�H����߅I����m]�t���n&�a�Q�u���兜4u���%1��@�^^/�袜�0��6���4��eX����4��d�S#��z3R�B�l� ��'C�8nZ$2� V�4�#��l�A�[!S���t�0|��6�u �敘�暝��.`l�\�kkc-�a���샇1?;k�k��8��$��Z���=����1��S.��� Be-��h�^}�y,�(
�a�9m��y���sU ���1Ͼ��	���Ӟ~�����Ҭ�W�Ԝ>�άR����;c��}�\$EG�ם�h7i��\�o��d_ �������^-�3��o<�����3�ZY�S	6�T�D�F�/3197n܈K339�/Т.fE�#���<����Ϻ��Kh0
W�w��⭦�F���j��$ϟ�1h�hb��U����T�P9�Ͷo�t_P��Jв�ôM˨��t�|�ĶN���S~����j�P̛}����9ddkE=��y��[B��\��K��7�ٰj�@���4�ZV	G;�Z� -�Yg�����x~1@�����W��pK���j���Ǚ[@�)e�{;0�&D<�1�J¿g)ˑ
�yk�@���:u*D?6֗�ʥ�x���-aR���q��7��g	"�[闋~F�3��>��?�i�ķ��F̠�K�v��Ɍ2����e{J?�s2��-���#����2�ƜINN�/��4ޭ���0��T���s��5��"��>��סNX�5C3S��$L��^�-�JR�5�Y_�ܤ�եꡜ��+�3�cbb��2�����R���63(ۋ�7<6�)?�+�i���� ��#���@
&�����+�~� 7����q�m�DwĘF_���'m���J3���fx�_���`�����`ث��;�S��)]�����H���c�g��U���iu%Ĩ��ux-1��2SR"�]K��V �tw
w]-.�D�׀�X�Cd�56�QnƝؕW�W����A���
�L��F�^�"�qv{�4{���䜛�Zǫ�:_���L�Jˀ!��V����$�,뫫�2���3�ʯ��e:k�ߔʽ0"�e6 穘�q�I�9;�c��FKb�spT���3>>�'���B���M]��Wc+�ˢ���]�,tc�)��=���u�v�k��7��/��4g�R/�[���G��#0��k$+��~3Li�/[���N��hz�{��C �8^��[/���D�� ���3;�ZkZ��.�|�����δ���0���ڵ�q���C+w����~?��M��s���[�l�&̸H?Z��$�s��}���+7�. ��a�+�5�n�� a�G����6����W�w�aE�M̴@������_�� b �5i]@V#�R�B��~�l��a����%�h�/�Ghtd4�yXW�X��TН3e���̀��k�[��1Ņ��{��zT#,��c.%����������F��@i��(���/�n���*�O����V�
��x^��~k�|aˇ�5m�V�����2W�*��VE�'����j��޺�l����w����~f<��i�rK��z;���\�ZP�A�+��ן�F�50���;��|A�1�2�y�BS�A@8 ��'�������&tƕ�(���&�&�nnp]p�"�W@�![M���Y2r���o5e��1N2�s�Ƶd.�qp4�&ݤ�K�%}��Zݜ�	df���v|�!0������v�&����9�F�yu#��)�����QHfe�e�#;)��Ϧ�Z9�<���q�����;s���ML�2���'(��������4�z�]�(��7�i):�Ց�q�뫱�'=�irjD��y?^�D`��e��I� ����o��z��rD�O������Z]D�M�u��}�u(���2ƌF�����#�����
�#�1	@����)VT��& :z�������u��xʱ�IK��s��R�Z$�#����nlK��w�L���������5��|W��P]�VɱGl��br�ܾ�((���B$d�r��y<}�֖��"�swK��X�'[���7�X́��1���ۘ�{0�`����̧0��1���:�B��0�ʗ'a��I:��E����
�> c��N��+cv.&��:<7����tI���f.:466/N͙�ꅐʤe1#�+9��癹
0���f�����4g����?>eh�@�榌�1��2���>	�Jsk3ݴ�}��o�`�k`v�Sȏ��)���3.�Ok�_�)w͒�3�_��@��&,y^Z	Z���á�A��K�`:��u<d���5�{ ��Ð���,����5~���v��Xez�������P�<� RG��rQ���N5����>E�y4V]�#�y�� ���֚��7�eُ�:��Х�s��\�ga;ڠ���r2��B�<$L����h�ׯ�-ӮY@p-��Lo4�o� ������TX�u��ָ���|�UU�R@��n�1�W�VwSݝ?��<*�S�TAyeף�y���5)�Q�E�W!��y�}!I�E���!ZUH$��+�� ~Wփ�?k������:���u�ӻē��x��W�9?S#t��/})���AW��:H�T�eT����0�"ڨ�f${{o'̬t�C���Nlo��V��G?��������`=.]���}�wieF:��BG�1��4��Lv�Cˣ_� P�p�����J3�Ef�*��-@hQ�`�@-x,,,��Ǐcee%ְ^�i_Ѱ���~m&�a��[��E��(�\qHQ7��T �L����n��] �������B�HW2Px��͸|i�΍5�u���[��/�k�:�a��tж�mv�a��ͦ���PP�3!����h���]�a:���ģ��X^^J�ϥu�W�*�B� ��9矂h���}��D�^�	 ���mԋ��|�q�J3�~��S|D��Q�ƴvd��
ɕ��{���O~��uܻ��,ց�g:G�hg}��66�5�
0����Xۑ��S�c7n�	n	 G���e
/h�x��p��weIk���\��x�r=l{�ocYgS/*����@����U�*K�J� ݭ<� ٓ���-���Z�y_�Ym�>�<N���� ���*�CPGXq��Ӥ��`bNf������k> ���l"4���wɘ]����9!����������5Mo7He�D?Ba���3`k�{�C���5����ca�5�ې@R��25U�n��ON��:���w�QLac@Ŕ<i�zj�݄���G��H<x<<�ri�2�H;�J�\������ƸN
9��ô�΀�٣���L>P }���Y���� ����K����@�����"f�\<�_ ĚX#\�	�e2]�M@��ދ;�IA��Z転�^K�k	s_k��L`����~�l�X.�h7��mYw陾>}G?��_�[���v�䘱V�]�p�ġ�FIQ����X�.�.J�����L��GZ�#�De��X���k	���
t^�֔V��q�|�ֲpe48�!<�K��Ү\�źs}�F��l��5��9S��"'�e��ja��*��������W���恕ɲ�E3���)?o�Z����w�FY�|8��s�3���rq~��VU6A$�TS�.�g�m�� }Q��!��ϣ�6�W�/7=W@q�{��셰 +���#Q�j$L.�Ƭ�F`�v� ����x^g֪�4фZ#��^�7�c�_�Y5\\	L~x{������=� �Hg8*Rز0�"cW3Mˢ��d\�����	_�tH,Ž{��ҏ@��l�h����,ȫ9d�#��6n�5�����n��͌��܊���@�Q��rD�:fBu�-�Gr���Bti��u
����=��8�d��j�����c_���N���;)�����LI���Ԓ�U��e@��0��o�U�����믡U��*�=*$�M���$���8s��T�������D~
ܹ�-�����@���[���e�*�e�k�rmm�_�����'��\�˗����x��)SԳQ���`��)�c�]���'�ٮ"I�F;�^pq.�kr�|���*��oO˜�s�*�CK�i�5"��J����V��s�r�hO�d.���1�DS�
����^����2Xȟ�s�lE��*yʗg6�5o�h3K:������\���F����(�
#'�S�Ө�Ӂ	�W����˱��P`��a����u�-���în�����5�1�z���'i�Cr��?G���p3�M�	�d6	�ze��k4�2���4G^���Φ����]�w�t�<-�w=t�`���u��X�8�B}���b<EuQa�ĥ�P(L৫��fnHǉ\V]���ه�[��pmm���g��<�˗�`�Lc��f{X(�<ǉnjM���6�؝�G/��s�y8�1����|㝂$��^��~?��ƗL��/�f�tO�o��"ew~�k�*�L(�GF̋���im�gj�AMv.�y�!�-nL��h]=�i�	�Z�������HT'&�d�^��QB��W���-7��O*k�4~36!H�C9��|�f�ڣDɠ&RzF�tƯ}��F��]�A��=v�*!0��f2��jI=��z�5�|Eo/U0Lr1)+��
G"ltf~� *BU����qKy�b���;؎����y��~��ߺW�`E��8����$j=]_d6c�`-����s�#W_z�[k.�x�dН�fl��K�ǽ;�'މ�w���{b��\�,,���F47v!�u�mC1}�R�0uO��w�K�Z@>� 0�����[v~�_@�c ��.0;���ζ+��4������^"������k���3�p�+g��|j�k����њg���&�����
,�ĩ��t�q��P� �ʯ�}���u�
Q���d]��0V��ӹ
����h#�'G2�x{})f����#�^b1�� �K7�����Y���S�"���@i� ��bum��:��tZ����u^�'z@w-�� ��=	�5���v��pu�N�������SW�y2 ?�u�E��'���Q4w�]Y���O�mL��&�ᆝC��a�df|:��#131��_��ujh����ȍ+�9��ۆ%v�~�5,��b]u��zQH�=������{���<(X��5��)� �.W5�&}�s���LA�(�9���l���t}�$x�^����G�ly�}�l��!^ ��-�8��T&2Hv�� �7��"L*�<�W@�5O��Om�
��ӭ��s��������t �i�$C�d
HG�����0���n������:�K�řO4��wrM�&@�t���v^��܋uWu�ܣm"��L7�Zŷ�	 ���HxS���+~r�&��0���݀�����=�to�GmdyF�e&��\�R��K>z�+��qw�A������v�<��2��d��[4��yf; �vڙ.ա�Grt٧�����-���\�C�1�W���2ׂU��&���O�e�%�����ǻ�8  ����� us7�DР��ԗÃ�/�)uUYt����]��#qq��*�䐴ny4���\4�v�D�?��0)/o��؝���[k<�����i�γ���}L�!�gG��z�m�C <�鄿�!,�
�*�}y������B&�����k��e��t�rf7�l�,��Y3�����; 1�,DA��?u���|S�1~�d3��--2g3���Fi�!K�|�"G�����ր0\Ո�#��*��P
�>w���he2��Ӫ���`'(P�Yf�T��浥Q,�*�gi����M�+[7F��i(�;[-�:l����"5��o^��r]5�uDp}��á2����u��
���� ������&:���4{ebӫ�)آ:��vf3e�6Df�ڝ�]Z��G�6����ߝ9#G�ź���4i�YФv|ߡ<iT�YP�@��x����R��zZNh�wϘ�'��3vC����ˡc�ts�P�������y��k^�qim�.��4{�������;��8��Ԗ��+�����H�e�'�R9�cZ��&)���@	�j	�ƨ WF(z``-&Ιu90�@��9\�f:m�E��OL�~Ⱦ��xP~U(�s�>�z:��;n�<g��Wo�c]i���I{�e�b�э�;@W��ō�x_�E���'N�/�tt͇q��矏�鋩�u=<c,Z{��}�K���r?�� ��O����c`�cX��	#/�\JN�Q�7��O��S��9*V-)�y�k�Ay���+J�C��/��M�!�t�ԀK
*-�@��2�]�DK$���U��;t�?�J%�<9��7�D'��7"3N�r���C�����)���v��>n&:���T�� ���,q�f�ap63]i{�ō0��@����l]^Y�Ǐ�1�7���+�!t1� 1�-@D�$��m[���qZ�孭�@;�jg3�fD&0�I��Ǉ6�g�\ZV�j����i��nޝ��^]GrX�Hڹ���5܉����ʡY�꽼�ƹM�i֨��@�,�-A#R'�s��)����/����Vt�D�{ց녛t �E�����y�
�Er�:�x-�ܡ.�5�+�x.�L��'�,��]
:�cnC�;M�6ZO��t���I�?ݥ=.�o��=1�+�9jD�@�ʱ�n�
@L Iz�_���� �hcKnll4.��]�<�������wMi�mKD������ؑ_y��1ǒ���#�S-�ܩ %෢��l�����n��(�ؗ��K���L��'�ty � �����<Y��"P�T%H��ݬ��հ9
�*"�mv7�� 	�yU���*���8���|^Kbs�����kX��Il�ePL�������w���� =����;͍�-	��ne_Z���b������2��!m�Y�d��\נ���:�p�fy��呚����a���N�:���.�Eف���:�������j΅������9���+Ӆ �9�C�؅w; G�\�w۠�m��8���tD����T�G�J�0�
��/8�"��f�Gf���Zl�6��_<툗#W�1�E����6��2�cÃ16�C}=�Ph�8EA�����)�I���l�N\%,���xԇGa<�H,	_�e�����TL���r/�Rnεrz���kфT��&���; �0�9�eh8���r\\G�<$ϛST���{������ָ7p]��~#f.]�Y;�NNW���e4�1L;`;���~����iY��j��2���i�Z�{�'��+[��|��k�q]8�Y�V���R�Z��-�q�Qy3��8|��l���&N�,2��Z
�7�f�����ف+[��������h �;ᡂ�Z��'�D���V�Fv���'W|j��y]�k�'�u�a�L6�Wn�ʋ��ǽ�wSp}����L��jn4�楻�K���1�4���S{��7r�vbb�����.8#�U�qt�"�G�)��p�JQ�AR��� �*~�k��͂�Z(�C�&��N6f�ec���n_XԀy�m�rH�
$��W/�D�	Z���p�a3�F5�vbl<��dB�!�WE��vWC�<el��,�\�܋���8��t����+ ���";0/�PN�5&59�l�Gq+�l��2��d0���	������S9��ō��v?:R�ԗ"����Z>jr���B�O�ona�Q�Ch��y 3�:�]�?Vpl�ﻩ���ϣ�2� ��^N�?;����a������q�\R����7���_�nV����,=��OM� �|�bi��b�/��m�K-���_����mg,,.�_����7'�C&]S[W������}À{�K �zZ0E�8�I�QPτ�x�D���4�b}���X�n��^���G��(������6� �e�2�H X�W�"���ݽ��lxT���5D��߻q�������Or��p��Õ++�70Hif���.�e�5(�m(�F�kW��1$4����W��۷�����������d�N�R���3�қ檚Vp-����0����G�I���C�J����.���ݺ`��U��iLG��~ӱ~�-���
���$/�*u��x	�L��Zo
0T�􍥋�s�1���]�f<C���A��70v  V`�`k���}'��A�oiq>�{�����w�׿�e���?��Ex�8Vq��h@O'��r&�@(�e�>4�/�6m�)�\�̯��\S�kXoϚa����Q��s*ݐKj%�:��%�7�D���$@���~ �.��3�L����4��j5
&�ɫy��K�xÏۻ�0�"�;cV���YP/ݧ=�K@���Ft�bqm#>��~��;�lbQ'��XP��C����𗟥}���Ѿ(����>�\bﰥ�-�@r��)/	2*���j�f�@Z��{Z��#��Q$�2?g��
��t���qL�e�c�T �`�e�λ?�*ؖ'W<ݼ7A������Wk
����T�L���IG��[0=�
�T�0'l�?O�s�bˀ"�m��c
�n����^!-��[�2��Ε��@3�5O]�oxd"��M\��	mj蒴�S|.�Ɋ�N�S?5�)�lsg?��3!,�-��E��q뫙^�ĥ��/b�CMm���1d��SLq1�cR���m Jp�GGw-�V6��8��h�*,������]��@�k�j�)��2�����G��F��~36V�bi�Ww�n�C\L]a�����d�V�����=�W!������92*
�C�7>�+|��L��F���.�����&������i.#T=F�|}�+�m��RV<d�~��`joZ�@V2�lL�X�VQ��	����n0[>*h\ё²Z�unG����������l�8[�����eJ���t/|�H{|צZ!u�|O٤?��;�\$���H��B����n<LKJ��e������"��Yϕ%\m�"�˴	����6����&?�N�������eTק�x�wm�m9>������((g�#�g�7_x!z12?��q.\$��זNo���+.�}a;�XJ��N�^�XO��z�j���g���X���,h�; dyw�+��u�!������� 
r� �J�A�{��t|�`5� ��g�sz:�&�iP���hi���4��� k��e���Z�\t>NW�6�;�`5�Ǩ�y<Ƥ>@�� hο`r�Ý�4������K%s���aoA�f���-pf�^�J@�	`��@��(�ʺ����
�Z�o����Ndt��# 2���M��r�ǂ,�uqf�']/ח;��g�;��-پ"��,dP��ui�|y%4w�M�#�ٹ'�0\��P�NS�q����b��dأ�XJƔ�.W��� �|�jm;���hq5>��~��xLGGY�ɲKƪ1?���{'���Z݂��+��SW�wq�x�wu[O��k0}ũ �����3yQ��n�1�{T �ʾ|g�tՔ�\���}.�l�ë���MF~����(�(�rE��A�/�>k��4��ڧ�=-�UQ~�y0���4F�\B�n�`b�ӯo��w>A ,��}ǺCt��.k��2��&�3B���}����j.����`���"�ֆ��4��w���"=�=ߍR�r.߃�e�� �mp�S2v1�w����$�gt8�$ݍ
��>�I��=�h�ת-��X���v����¾Ad5���
9 �>X����yM�RoAC�,�����P��#c%0�Ǎ�Ȁ&�IK���J��o�K/��X�[��������
º��Y+Dbl|�}��?y�t-�ڭv�9���4�^}�Ź����օt�\jF!��O�(��v���ow��G��ڰ*l'�2!p}s=WsƱ<��d{uO��@��>cc� z�k�Ӆ�os�4��JooxZ^�[��������btS&L�	�״rz������P<�`tA��c�8}�F;:�-ң	�iS; �Z�a��x��Z��p*C��3��C�f������<%g|�<�}.�����	 ��$,�Y��v7W���������k�1A�c�5�&���7��c2��f2:䖾9ߍ��nR����r<�[��ݬH��=v�iV��ձd_�������ow�R?x8�g�ɜ�� z&��X�Q��L��?��߿;�����q��� tB�N���#}m��*����I^�g�h�@�I�df3��&�&ƥܴ<� v�}~�q|����x~>u�)�g��e�����繾��Q�1S��������v_r *�� $8Lt8ґ�2Jc���R���1�X7 R�>���I�����]�מ�� ��D�q�T�KW���ŋ31B����?N[s�/ S,̲.����{�{uZ�U1��I��		�����ҥ{@}ݵ&��� aSz��Y�Qfkqz����Q⳸��:��^V9�<BK&c4��k{�o4cmc+�x����tYJyUe������9�#���E*axK�;:m�NO�$�u/�h�y��G�"L�B�^y:���!G�� �-X;r@ONC�eaZv����YIh��WaY�3��;��qP���}.�d�-�p˜v��LF��ي�����=��on^��z��_��Y`rKpa71Ǆ���) Ħ^�n��_��~��_c<Nav�Asu)=�#a<f�	|���ʘ��q��&3�(��������_����8m��>~��.��;% ��H�a2�Zz��j�E Bhm/����:��;O:b��L{A���oJ��E
�5��9'�-.,���\|�����Ν���'���\Y�c���w�?�0c���oމ�ۻ����XH�:��v]"�6�A]	͙�}���SB�abAg��<vN�cL;4m=��܏���� BgW�/ �ͳ�����š���V<���ϕ��m���7r��.}rb
8"��w����ܣ�c8� ��0Uxn�KZf����
�e�R�3,?-��7�¾���P7n�14�uuI_F����� `�H>�rJ|��|i�@�i��X_�������� l�ɋ�1
��"��ʙ͋/~)n�~!&�'i�ﶡ�Z(�6�u�o�v��M�sJ�������4�s�2kǄ3_�%��_��QE�Tk�̽q�Xv���C�N,z�T�Enl�Q"�W�bf9ƏG|��ܠ�S�j >�� �?�sS(�T�C�U���h��Z�[o�
*�^�% l��~��'��tc�t�Ct"��m,��6�
���5����$�@inҁ���M��cj���Pkno��å�嗿~7��x8��FuY-��3N�� ���WO'�Y|�BG��"F[m�Z��U_m��Y�����^���zk-���c�x+k��e��ݝf��n��ϑ��!E�w����v��D��S����S�������Y�`�0�Y��1���k�oF��s"�u���-ߠ�mU�0�2��2�wZ_�[�bm�&;�ָӣ�����w⣻�f��t�6G�x�ב�JW,�N���@
	��Z��;��Zn��Ƀ��h�����X��I^�՞C��*7���+��.���cŜQ���?�Ela�j��d��w�6s�j��q���1sa<3Ou�-���ă��s��g9�U� �K�v�s:�݇�G��� �ۏ��= �ѧ�����C�Af�
L�L���	���n���XO���1<��~.����)�"{Ũ�p�)Т��Lg����չ��%;e��;��S I3�㔖�K-J=�Z�u�U����\��L�F�"y4����[q���4#)���Gː��Z��}�@r��5���`�h���9e�
��w����? @~��^�G{n���.	V��hFo�m��]1�cĔ��!�e�
�>.�Z7]�;:�	k��؈���B�8���7���dF���L�73�!Xl̅�)cc}#Wh�w�{�/�y���(�"�#�0�4sԩ�O���[��XRh��Z��������,�f.������1�c5�V�2�9������� 8��jݛ�����(�/��6���2��V6���b��R�t�������M�2�-�����Y�E��%]_����b�:�����(�k�����q���JHwy�{�^��λ�+�1����bq�J&��r��չ���|�A�--@[\0�}��{�0���<���kv~�&.���/�~�?���E����1�j%c)<�k�Y�ᮬW.M�D*YͭEy.r��Y����2ZZ�$.�a��4-�#��yo��'@#s��]���r��d�*yMum�m�3��Z��x�;12��ͯE�pƽ;����K4�B��ƭp��-P��n] ���U�r!ϗ��x��s~�/�]WĤ��:�T+n�`���?���n�H�\,�z�X��R@��2�����6�9 �4�1{�u*�Z�R?^WB��V�%h�>̼�E��.{hׯ�90���|�����L)�V
�o����<���̉��<�Ϗ N�4�_+�o�@L���Y��+�؊u���)���~r�Ï������9�:�*��\#�Wv:9�&�Ϋ��g�:
t��!W��Z��q���x���r��kNu�!}�}�{����i�s޽�Km��A�ub���~���m��]g�у�uy!>�����G�L�Ӻ�B�G�]{vh�p�ٳ� �`�(�֛
D tU�|���B<��C>�������8��N�<ܦn�U�a�5z㵗nŵ�3�ht�~u�A�woKQ�TOp�B�ђ_��E�1�kY���pL,ӭ�*�}��%�Ԟ7�#ߵ�l-���0^�}1^}�y�F��\*�2E8�/ ���h�w�~+�u����a��/���Qo�� ���PRZ#�L9�l�T����cY���[���L��wu���f\�4���'1V-Owr���}����ƽ����� �f�@�7���E8��)5��Hv�K�Y�(�U�(�ª�`[~k�0��'g���a�|����[1z���J�ejp�趶\*'��-�Ϛno����h��p$�s��'0�39M~s�{ ��F��Vi]��z�c4f���bZ?�����ox���/|�.�������խ���E�m��igj��v��L�)�ԣTMTK��6��G�Y�@I��]m�ݶ�\䣓q���_Ȝ�3Í1���x�d�6Lz5�����e@�Z;鮛>:�e���ccc�vuĥK���k��1@9Zk��djG6�%��Uo�����KiE���j�tt�n��wH=Sf��&m�Ѿ��q��7-v��L����J��iS7�@�1���#굺�����`O�� �/�� V
��F�D�����ko���ona%��?����_J��������bO������t�RP���~�t��*�U��q8���Ĩ��G�t���s��ȱ��q���?�w�o�q+�)�� ���sA�$��~��x����Do<X+ �r��g��ktL,�U b��4���o�ύOm�ҳ���g�Ϗ�5+ ��s��_�����htӐ�=�3���?�g�2>���wq��lP	��RO��9����,�t�@}v�nHcd4|e�����6�akM�{0�����aF�լVKF6oA��IeD�P���)WPR{&��&�������p7�̗f��l~��A�Bn��]NO�ܿw/�o����������i벱���ԑm�1]$�wߏ��ǸnXh���a\$�P9�eZ5u3���fpM7��4h	�ά����P����pɰ��]rlcc%>���X|G�Z�T{�i+�G���`�	�洸>��o�ssm#ip������of^�VU/�0��U.4X�gR����U���IҘg3J;��� 7ehy��}׋�SFv�bPy�Νx�����Q���:���p
9��c9L�Xgg�k�ݾ�B|�˷bb���R����$�1;GuT
CC��銻s��?���7~��],J�g��ѝ�﵈r��OK.��~��� z��@�N���U�8�,4�Kf"�2� i�8M�;���n�vc*zi���9��� b�һo��y���7�/��_��N���K���iK�M!Ҕ*�By��ϲ�����)\Sn���V��O;4�d����_�R�����G��:@�u��;;[h�m:���ޏݭ]�Cs�Ew0�a��CӴ����r,,��"����83Ԉ����b-\���M4���H܂��&'��p:�k�2��O��3�=��k�����Βt5150�ˌ�>5��h	9q�7��rN��y�Ԕx�0=:�C1W��8����~cF�:rT� ��~�m� �h�A�҅��]N_o��s���QAD-���(� ��5�/���7�B������n`���n,,<�{s�F\��嵘�uqi���F�pe� �mp��\5��L\t�'���v��x���1
������|ߕb�P�/��N@ �P����Q@=n�Z8w�v�D�{����Z^�n=���o9ƭvϡ�v��n��I]�#�<iY���8�A��+4�G�Z�g ����!?j1	.���)�W������?���`��>�Uu�<�Sʹδ@����X��ش���D��)��}qV��ak}�C��S7��:��p0��Vcf�/�����kc�������M��?����iW|4�Li�7b���	h�i�v-݃!��'�ώ����Wmy]^�ԝ��0�||������C@d+��%ώwAV׾�M�3\Ys�x�Y��P[K@���C'�}�����ݜ'�p����4�nlmo�V1�*�9���NNL�W��Z�i�HW���1wM��2*D���\4��zfr cSs9<�u�i;�':��%ǧ�G\4�!YM6;7k���	L�rhVڽ���u4�s ��Tt���f�R-����*/ݾ7������n���R�>|�̘�f��'�i��A?�΀1?l2B�+7�Cf�=sS��s7�v���撁��Vcw���)\W�]���n�~�M�����[�"Ҫ���+V'�gPy�-�F	R�ku	���ɱ�l�d?Ը9�_�"�y��7�|��Y�vPI�Ȟn���V,-�$���S��uޏ4:�ʚ(q@����X�4�LQ�E, h�/y'(�@������/����,����0���١v�J�<X��G*��Q[�.�$�|�;��E���C�4~h �I�*lg~�wFwm86V�cf���|/�rs*��6�g��|>��q�	?��O!hG�7���g�n�h4M�DxӝD��[��U̒�˦;㨊'
x��l}*�>������m���?���4��0��G��oo�QF4��(.���w��t�~F�)ϑ�n�Uq�� ���Y����v����P˹:"�:�ܞC���k�`�6AA���ܣ�d���D�IY�2�~�f��`����#
ԡf��7�[���jn� q���}hӌ�3H+�h����,��(�) k�����f���A���ř��}�V��U3GzP�q-�B��C=�����y���*�%�qcCX[0��s\�Q:��;��Qj��N���n��&Y��%	���l�
��s�ҴN��֟�.�q
�.��D����}�Ϙ�� ��i�.��fЬ ���Q�gL��r4��{�󦜽���
�G�tk����,��}��Ġ6|Rќ���ݙB =u�Ա�Ӆ��;���7�*�ֿ���'��g�Ł�?�l;�T�&����|�	/��&�g ��^�O��GU*��,+߉̅��5r�1H_�b�lz�;���k���x!z LW���� B��Ə�3~vŻW������<4N�D�ǽ6��ۓ�fpLpɦ����ꚼ��Y�'5�3A$�������ï=����1����4��������w�Ws�C�$��#�|�P���<I/*s(�aU}�\ÁM���} ��Dc�����s�W5�O��Y�Am�ͳt+�F\��Yi
������K�U�ظN�+@��"�����Q�o67���	��0��뀉�7a�G����c��@_+Ͷ��Tˌ��e΅��D� �C�s�}}� F2-}{���.�E��J�/��ƅ���kc����u&���/�R���@_a��۟��9iL��/\!]��%���g*49����"���s���J7������}(�YFZ���/l��2��F�}yWz�RG�m��.e�&�#_� �Zt�c9'�ϲ��� �Gߖ�'��}�Q��|.���a�G�@:�d��UސG������2c:��K��,���/��g�J�������cWZ#Z�Z�����x��#�Q�O��c+��HO���\����j�X��,����?�9��6��~�^l�Θ�ؖ�i�"��8��f�֞M I��/-6���*�խ{تo��yvl��<w &��7����������ah?�ޏ%äkC�ۙ��9������IB�_B�6.�iF
Z
pZ�����M�j��]�K�u�D�R'*iB�E�zOl��%��9�gh�4��������i�(��H7J4.b�X��	t���BȮy����E`Hi�kr��;Є�����(@#c�hE���l�㒞���y4��ޙ�]� hL=��uҘs+l�	c������1AE-~�8� Mm��	pZ%��o�����hZ#
��ֆ��LK�+ I#�0>�+"��mhk�����̀1�;D-�>8�WZ@���������Ԛ(��( �0�[K-���\��h��9[���쨜���보�c��ʫ`�m� =�e S����NyE,C��^۝ej!�FwAݾ��ǳ�b�K!���-a�D0NMu3�W&��А:�,�����X�@��ë�����s#���/�X�k��B �8??��/��>^܎����9�B��P-L�Gey[���O)~<�I�K��JW潄)�8���Oj��#ʩ� j�FP�~�o�3���X�����k}`��:&"T3Y���w��|�����a>�r���ژ��i%B�M��v��S�N��)�'~��{�$'� ��tN��,��EG]+�S&�:gZvAOGn���[ﱶ�v��4|���U�kI)�z!��j�ߌ�\�85�r����lNy�=8�]8`��9Cغj��,l�:,Y&�I5� a���`J#�0��-����^!}�¸'�>�{����[�A@��E�Ho�w�s���͹���!lqW`~�A7#���y-����#�[[ڒ���g�%2�.��m��R
�#E�rtU4.5���lB׏��ܖ�0N6=58ve�-�Sp�.���rIK�z��H1r˺[������?�'��7�b�� �2�fN
�G  =]f]3����"к������F!�M�f�����������7&�+3�A��ZssU�������կ�A��ù�����.y"��c�"2�>iQ�$Z��eU/@%;�
�1�V�egr��=�W���w��:�u���"�\աQGE5��w�G�I���}_��'����i�2�P 3�VA���my��ڻ��o��z�P��h HkGpIK��nD�;T�-�����`*
���h�X'!�������=@�Y�!�Z%.l�L rB�5�5?M�t���Ӏ->,�:H�@�k���Xk��a���7�~�樔.	��i��g�,���
�.�{
5e��-AR�F=��<"Xd�gz{����^�_ZЄ�*��Rq���=��q�Ij����B���h�s� �*[lK���;�d�����R�1����7���P��ګ/� �	��5���UYG�����a5ܻa�F�~N�����9���:�����]2�϶��j <�B�"�mK����<�f��u���P��U�>F�i� PV1s�f/Ji eՍ��{f��9��q��G���pw��S��3���(����[sgZժ���N�Ü��t��#>x�G혎X&�!��?���H�mD�F�cO
��ڙT����SQ&�|9Ȟ�Kznjhͭ���jV��˒���e�޷����	]�!<����42��˽��=|�� Թ��u����+�ܜs����������p}�>R��(S�ڕZ��¡?k{-�O��h�qi�o65x�Os���+�UN|�a�B���r�٧�ہ!7qm\�f>m�l`],n����^l���	�+�h���3b��kR�}J��Ly����aJS��dȴ,�_`)(��k��D/��3��r�o��*]ݟ^
����n�4纹�߾7Ǫ����jT�u2%$�0�2/����P|R�����'��/�樔���j��ҡ^�+[j�w�G|�-�1���L�2��{#���ٗ��uc\IO��"IZ�|���yD�ޮmh�U��w�~*'�o�l�����汤;����@fgѧ�R ݲݔ)��0��C�<����0����um�j.��� O�u�Ƌύŵ����Ҕ�C@�-7�������(.V�����g72���V��Sq�P�����`E��ܧ��Z6$����E����|���~����N��q�Hܻ^��Ԅ"����g�î�.��CL��P����h���P�V�50���l�@�PȄξ4٧��L��WުF���d[�����*�o��d$�wߏcl���� *� �y�,�����sl#M-t�;l����DdF۪{ef� �%eU�ǝ?"���`�Іu�ƶ�D�� (���/�G��qk��m�*��]���'�<���~Yw~˼2��B�m�{u�Ǫ/��Oe	F)��N&�[��~�+�vS.�j=)�v7�|��5��;ee?���1�ϥ��í�>wH�]a��~DL�JWSJ T��uƮ9} ��:��� Z Z�!߭��!�����-�W+�	����Պ��X$M!�#E��f���2�9/�a�ֿl7{���^'�u�,�NZ����2]��aw8��h]�I:���6a���//��@[����[�l6�\����pg�cgk+Adem3> D��o��y=v�֚�GNw.�Y2�9ZC���X6����y��+Õ�W�[!ĳ�(����G˪A��J�\��m�i����4�=���c� ���t�c}}_��giݸV����3;*�_�����d��۪��#�m���#�X��^�(E�8=��}`5�I�P��&�����`]�%�QK��c��?�|Rq�(eN��"����ԗP��Z1�P�0�@g�"����0�0�f}���'��t�䙾��\�o�&�^.ʣ ���+-Ϟ���}����tL��L}�IS��3I�[��Q譟�w�A9d�]�-~Up}�O����z�YfՆ�Q�]�;U� 9�ŗR��Y�>[ 98@�z(B~�Ȁ�	t����:���M6�b^��Y5�=��a:C��>|���2`��BR�������*��i�l��v����Bk�P�����\��c>��剒ãbp�Fz���R-A��a\�5���څ���������ywL��V}u���E�v��������c��/�@8�hP�Z��y6C�%��z��ڰ4�`z}἞cU`5�㷷���e@�AU����mS�A|:��2�p3(](u�Lae'��w�{��f�/7vQ����A���8���<�Ԅ�u�"Y'��j�T`���Z-�̆�m2���k�V>��=V	_�
��0��b��2�tpb�&VV-��j���g�\�?���
�;
�ӫ�}S�0�e
��Z$�gc���*���֋WS_3+C�F���sRԚ*%8

�"(�����-}���F�v�ʶ�[o	EK�m�O�C���?���ٺ����C�o�X��oi*�x����=�p�+'����������鉉x��U�b(>|��cW�7���TO�'��i�xyO�H������v�S��0����T|d���L��,@��n-�B����Ge(���3�n;䙔�,�к
h{�ɌǺ�j ڀ�s�2S uTR�x]�H7�2�kҢ-k۾���w�{;F8�0{� A���O�{��J�v�̳���q<\j����KMSbkq q\� ]��n�%�&3jf{ގ�F[C�Qp>G���I�\&��d�	W�>�yt�lYH`��PnL�P�+����=.ޒ�l����x,���f���zn���#�W�g;������ά���J��t.��(�*$}k�5qMU��AF�Zc+������]���u�}�#i�v�<JR�F`
pS��y���ip"��*sS���ҧ
�����k����ȸ�Y�.��u+�Sڊ��IW���n
�u��G�R'�GPKf��~�6��^_){ä�c�Z�jt���]����zi���]eȏ���E�ta�!�������<=�oތW^�r��q��G��_�w�ͦ��ڣm�d�g���:��P������^ӓ�::T|���2U�����7w���a߬���w�,�p���.�'���ɛ-��ӂ���,W�p�$0�G���t�Z�f��M6s���C���M�ܓ���������2K�Zjv:J�M|�S�K��nVJ<bw�5>�bnn)��?��q��\�u�G3���50�LDf� ���n���W�*.�?��g6�HFa����$�[뼄��M2��o|�׋�%�R��@�;;�`Z
��,�F"*�Xn�k9��V��%b'x>c-k��1�U����
�-����<u��+I���>��z}֏MaJ�϶x�"i!�p�2�W	tWB�dؖ�f�)GF�k<o���m��f2W����8�-e��Z��46Vd*���(Pn��l�c9.���0�-�\5�k��CaB�R��V���k����C����'?��9�gx�Ih���%�eI������^&�����O7��u[���2Il�TP�Q�۬�י�l���>�w�I��n�~z\�5����ٗ.{)�+�[P��<`�t���斊����M�/Vw�§�<�o~\]��ׯ#Z$e�J���~�Ly�$Ɯ,�[���>
n��ڟ
7�N!T�q��͍f��_�8<���L��!���A&��E�}�go
G���wlv�D��K](�2E���U����z�B#y�D,���v��o2��^΋���(���S�vy4˥�ݼ����
��Π���V޻[�欌�z͓��w)��� $2�1��;d2i��M2V
mLl*��RV?+�)qG86��3�I&�y0��T�9���y��Y�#3�����
��2���u�|��R���
�1�����A�[�n�tvZ�v�S��\����T�����fe]i) ��`��͜sY���A�����T �]	�m�~���#8�w�]�6�6�<^���w��q�q�����;6�Qm�g[*~�[uo�U�~��۳��S��ߵ}V�n����U�^��5��,@J+��R\�����j��<�qⷷ�փ0��3��I����1�d�k��碪!U%���W��"�D�wl6�h����~6H?�����Y6{<�KeQ( 6Pᠵ0[�V�Y$`"��<"��@��*ư>UGVϴZ��b� ��a�YW�_�]�^��n�y��sK��8ϰh��������� �o���̀�2�}#\3�J�uR)P��+�b���o�33s����_�������.T����n]_Kal4Fr��ϼ�ܵ���N@��7�ۧ�I�(�m���X�	�(VV�������e ������v��8�ey��q�^��V�Y��M`@s62�.�r؜���쩵�U[�S���O��s�^����?}��>�{�������k��nU�,��2��V��!]�i)ml�����OA�i}9��s+~t��tt����B��T �F)��K�V?}���8L����T[��G��������O�)����X!ON<٠GnZN
��H$�̼'[�yݪ�U[u��,�v{�N� ou�nkݛ���b�j�����u��´��er�oՉ��h�^ ���S	V�C9�S��-K���U6'����s���9%�V��k*{��%��Z���2�9i���bH��f�k�:tD�zZ_��s^kk�X��q�9�`��3u�+�*�g��U���e����� �^W=��^�@U�WeW�׹yOҖkܪ�g�U�Ǟ�|v{����>��'����ݼ��u�}��j�>�jO�Y]�^����^S�1"��xz�T翹    IEND�B`�PK   �EX5&�ܐ    /   images/3b95452a-4474-454b-80ff-b9153f229806.png�WPZ��<R��b@A:��H��^B C�&� �GB;*��#zh�&�$��P]:�!�˙�w���p��{f��Ϟ��Z��k��&F6:::6]-�u�����t�B	��9]fo������K����!�_����?��ׅ�FK!��~N�.R(_׌::@����e�zVp��phg8��4���_�9�tn�.D���L�ph<�Z�+�K�D$�}�چg:_ȉ�!m�bDJӄ3�:gf�FQy/�Ҭ��#k��фО���Ń&9t��FVh��tj�@�p���8���o�!!�*|����P�_2.��W2N�%h�3�������v�N*W�^a��cJ�<F~�a���`~�׵�*��0�{����I.<�
SE8m'�j�pӪ0�=z�Ȍ�����GV��w�]ef3n��=��d�ޏ�*4�}��Puo�f5rE�v��e�"-����s38
��f!$&ơ�Ur���<�=k���]�������	���+�?s���R�G����Y6D7��Q|y�Fvv�1���M�G�tU9eB���,�4�/>����Tj�T�QQKu�����.O}�-�yle�d�-Y�~����u��8��\�Mwym%9����6T ���$4 R�oi�]f|,*r		�i$��τ�n(O��ݎ����w�Պ����v9=��6钃A)hw�N����g������������96��$�xe���~L��ujN�D��S��k��?��� 6G�A�}���T�	·d_�U�l���P��gDM�r��,%Bx�M٢���Y���Ҥg�����k
/feK=�H/)�r,��
���
�[��tl5e/ӷs��xd[�`V�4r���Ty���~��Q�L!Pt�Fu���r'���;4��dd%V��x	3s��< f�������6���2�\���{AB"F]sCj��}�4��D�*M#$x*�ԤY�{'������6����]���^�-��4-���s��s�%g������2�:��޺���ְ�Rv��t����	�q�ݧ�=���$�>L��)W7[O7B#ߓ���h�#��
m��95��"._���r;[��Gx`�jzi�q9(���ͩO����㻋Hb���Bl2�V|�X��dV+'#c�r����g�`G�C\\\��?r5�6��l\�f�D�4�ъͪZ��&k�|��z�/�x�p�c�i|X�n�o,7+�īU�S��3	h �Uy�qk3��ù�*�����q �(�A�~��9��pɍ�z��Gp�S&�KX�3���U�u�ד74��6�:V�U\c���&7�F��Z,bl�~Z�[g���A0`�-
�g~��^�����)��gM��&L���_��]�_B��H�R�g�	.���������Auk�\yC�9���I�;�r(0�v���q�<�X)��ȝ��'�nq �!J��9u���ي-���D�O!l�G���N��"i���YF9��W�'!���T]�P��KM�sa�a����S�� hv9�
�����E�x�������/
ZZl1LA�'����?�E-4����-��f^|�O���:a/�'=Ր9�Ŭ��dǞ�D����H����91�]��_��ߺ��B��&�JZtu)q䊧�5S�����6&��|��p�Ec����|H�^��\���r0���_I!s���J0�"��>WgK��1}:��F
�6j}����Q>���D�*�<4x�ǒ�ml�Ig�Hd� :�zn��n�b����u�_�vv�D��ӻ����>|�E� +��M�;�ێ�3��,��#ʏ)��߂z�ֆtBW#�{iE��b��~�P��;m���q��Έ0�����[=���?$rʄ��,�PN;�'�!S�3Bs�v6��8�ݒ�ǃ+X�<�{��'�q6D���
#�x�4zc�A��@�V_�4%%e��#(���ϱrziJ���R
gQ����P�,�3���{[A��-�w�+	��n���ޝ̲$��SN+]�/H!&���&���� �X��3��N2�<�_\x���;F6���y.jb"���[.@��R��S�79��Z#/"��c�0�4�M�M������O�w���!O�{���#�w�gѕ�N��o9 ��_0�Řri��Ȩ�����.�+n@��7���gM$�[�i�k����M@�/}��r����O}����Y�g�'�Q�#��5ww2x��ߞ�<~�I',x�����.̳������X���=(x�d�L�VW��MѯT��ֈ�|�e��x����u�u]w/�����  �G���R0Zk�u�P���ɑ,}K�u�4w�K��Y�y�*�yq?g�^����t`�s��,qi��j�w/Q���s-����
���* �ɟ���[�e����ͱ3��fǷFԊ�|)>���b�>!j��>�Or��|B$�N�t�Z[�z4�ʸ����]6L�U�{П(={3��f)Y�E���`�1�?\��y ����!(���m���j,����r��&�A���կC�����S�I�4�\QT\XH��wL�Fd�H^m��5�4l��:�vg�w$�'�č�?kl�[n�	���*U%Ņ\�/���6I@��ؗ��� Gb����/P���ܺ��\|�췸!οJ4] ��f&�
���k�����N&ay=�{�z)o�;dU��E�&ao��H�]����$(��/��â�"�cq+&Z@��I7v��fO\�s�G����t�^Uo��k8�?�iO��1�L��89���1Oc�oT�	6]�,��}n� ����+X��+K�7d��V�aQK�J�++ɂә��4��� ޽c9��::���̷��b�߁m��P%僘d\*0M�P�~���x�Pڴ{T!���H��#|��}�f���k}�X�K�UwP�m��6V5o�m)�p�9h�)�����T�/�!IN�
0����d�a���BI{��������c�G&-��
<*&!P��x�ϯ��0y9\�D�F��j*��0�˵�
4�-^��k�y��5���P{��~^�'��l��\t�E�r��t���͆8s=?;轓�gٻ&�BE��l��/��#Zb+^��W�2q+i���Y��Z�|c���G�����]v
s��f���Cwf���Z?���|�U����������8�u����a�z1?�6mx�����Cm�T�; �o�J��������}艏�|�J��'�\\\�X,��{1���Q 
��z�"e�:���嘦qR�J�8�9�[���b�~kؗ�g7X`bE&_�Ğ�ظ���f �
Bh�z��1��V�N�˦�D��(*b&V��|ˇ���l��.�<�S�9ô�7���}%=��zH٤]-3����|�k���p�Y��D�_��?0��J]����{P��f>~.�q�NxE����d�s���UKA)��AC��_�i���5������̓n��,|ԳT�v	o��l��_�i�@"7���)f��q']p	��ݠ3q��Ȅ0��4�����a쓰3F�f�� ),A+A��K[�G�V����L�C�����=�
W[ws��/�����4�q�y�~��z/�{�e��y�7j3�6����V�#7�ٱ���D>��N�_z3� �h��S��w�XS}VS��:=����GB���[����k��+��~�'�	����������[��N���\�Gu�D�]"m^aO튱�ꐬ�����=P�/�?Z�	q�����tq��B�S�O���Z�f��-�%��!ˁ�@77Lc��e��c(O��C�j�s�ۅ�\xq'����U��O���四�]�8���ԙ۹-u�v�q���ry7J�s���6�j�J³�	�AC��U��c2��ds���~�=\{��b�jiU����7PK   �EX+_-�$  �$  /   images/674f1970-5ad9-47d9-a0dc-0530c1f88674.png�$@ۉPNG

   IHDR   d   @   ���t   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  $LIDATx��}x����/�RH�nz!!�"HB�b��HDP�Z�(蕦���x��@ ��4��	%Jz!���n��͜dæ��߿��v�g����3��dhLLL,�z�D�:�Zwj��$�?h	�P��B��B�,���I�I`}����=z���:���Ɉ�������GG'����^^�J��̌t�˗/���B�|�p:�>w7��{��y@@ ޛ=�VVHN�CQQ.$&��ƴi���+V 77�����R�wRs�ooo�9s����w����	��
���1��PZR�/��"��͛���jK�)�����O=�^{�u����l������D(�������6���}�>�]���`}�����BCCі@+P|2��;=(��S&>�L������G#���ܹ3V�X��?px�Ix����ڂ%��2q��i�%J�\�%��صk�T��o�?�Ah��ʁbƌ��_"��'���PY��A���>rK�v==ܝ<��3�c�XN/���Ӑ��Vg<����FRR�_"������W�
��tqq�f�iccC�W	�Z�?��m	A�:��\A��c@`g��������_a{ȏ��!�` ��t)t�����¢����Kqq	6o�/�����q�ĉ�������:�555��3�}lߺ} �+���53�3�{{9U2���,�Mg9;)K�y&��Ă�7^�3ާ�~
OOOЋ���*�~�W�^��z������Nr�ڵk'��A�PRRB�X&�0a�
�E%�N��J$�v#��>�G�)��������B���ֲHO���Re�����-���k��p��{�q��9�����i�i�ϪOjO>��SHJ�����'WUQ�� �I������	�B[�v�r�t�Z��prtX��w�ј<y2��ӅN�h49r$�Z�Xᬏ� X�~�P�{�쁫��  _gn����SUUզ�``�HI͆��}�����ر#TJ%�G��ٿ#��r��*)R�y�Z�8�WJ��m�=��Lq���T{O?�4BBBF�0*jن1��5������y]	�U���0;���s3S,^":���t��V�����v�����E]Q���WR*�����Ĉ��/���`;!!w��iR����g||����ʪ��טk��q+���`��۷"���x������������`���󋥯 ��^��j�v���j�՛�1`�@&���t�v�0f}�x�?v�v���X��ZSu�B����9ޙ�cmG��/�cX�3'�W��e�.G�C��A��*;�B+Cjj*?K�.ży�����í[��a�����m��I������Y	��2G�Nw��C������Ϭ�3{�:�x�,ꎚ��'UiK`ckk��i<f}���J��ӄ?��qJ�b�3"�2�7�C�R�Ī�'3pҤIB���ƺ����ߒ�<�^G�"4�Q���ݐ�5�J�*���¤�c�q@F��q�Ɣ:���`"1��J�!z���
K?~�kXq��i��*���+2�
����ag�H�}7YS'��1b�);v,<<<��?z�� PJJ�P��5,ژ��~yF �3�����������l20liN<�nn*D��|�4���z�g�Ǔ���@8�`+�W���G� }S.�u0)��Q?�Zd$\����� �����r�W$#�{v�ŗ��
qBAa)U6HM�ann:(&.��y����;�$=y�$�w�.�!6K1e�\�r��Yl���⋸}���-,昻�8l0���&���;6n�H�w�P����#��\���u��S�N����ւS�0mJ�s���W^FT�t��=06>�1�����3� �i�<�1nfS��
��ꋨ���Q��ڵ?�Y���ah����T�C���@^j���������H�F�jLr%�J,ɓ/&(#t	B�L�:U ��Ä1��nܸ���ۣO�>(..���}ÍMg___�|�m�on�h&���|�9��<����?.,�cǎ�)AN�>�Y��F~�\_�P�'kj����I�XJe���J�E�V������t<�¸��=	�v���1��q:l;y���J���D�m�f���CƐQ�����I�`���x�GD�W��Ç��7�`����a����>����l��KX���b�����e�#����@l��5��!�����21�:_cs������^�j>��C���
���9N�nvѽ����ia�� ��8�>w��xi��l2���?`ɒ��?x"N�?;{���u��:\�6vrJ�dh1�Y��_q��Z影h�":t7oV;�o��V�X!�!�a�8���&�A��j�f���^;����5�[
gΜ�6�"�Oz;w�n�29���
�8V�UĹy���E�q��r�������q�܄��u3Q1�Q�-?�������k�����ǫM�����8�3X�ϟ?�U�ᶒ��ؼy��o��JOKAtt$��y`}-�[�ͣ���݃u���s�f�C�Wػw/��'D�];+���ȡUzh�1=|j4��B����?�p9u���Q"�C�$K��EŴ /c�ʯZo,�(B�估�>�<~��g������� 8���S�A��z�3�S蒲q!";����F`�� �^n��f�R���xU���׹���#���c��defN���G �����x�1\��5V>&�?`[�������^�4$�^��DIaJ
҄7!�,��M�_|B:94j2UK�y����4Su%J��k&k��2�n������,L��Ӊ<��,[h�	��ū5�|r�z}��<ȿ�t/�9�����edm�y�i�X�a?����
�R�t2|�]"LaQA��FPc!q�K�B=��@?1)���V�6֧,�YL���O��A�N�v�Z�|H���PVd��ػ3^�3e�8����ڟLKj�Q{���L&�̶�ab����Z���E%j��Fo[���ۖ��������}��W_����a��A��κ���"�\B�!�����	/����@����3���Å�U{��PNEE9v�.��K�s ���?�mۊ��P���-j� ��Wdd�#19W�ߟ#���<���yr(�*}�1�ڵ���rޤjx�����zk׮��y#�zt�~������#�I��/��j���8��8t�zuÆ�8x�`�o9<�q:�Z�4j	<�'1�H~�{L�'��r�*!)C�y�u21�������x�k�qL7D��� ��:&9s��$2�rx����]�����u�ѻ�k0&��q1�ɀ�DP�p\�p	YY�b^vd��Ù�?H�������Ͽ�տ��WT4��j&�j.�+���tƉ��볤!�j���ʪf%�}���\�V��T�x�ѳ�0�t�ڕ��Ik�r�L񓗛��g �w'���,�E�s�m�y��� G\���Ͼ���<k��:]��m�X&��K��g/�_��E�Y,#tΤ�Q����1uu�h���a0�3!��̡�������5�'�^��7P\�th�%�����t	����@<�d�oײ^���";-#G����?nr\� ���R]"nq�KKKp�d8~�x�����!�_gX٨ �*��l�nݺ������ΌA*5�\�ѣ+�p!~{�M�S�ͽQQ]�d�[���\I�o]#U6���+��K��T�w�����^��o����}��؇���Hۇ �Q�-R�sY<5&6�=�̴��D玞�:y4�_�]���ħ#>1�>?�IC��C!�����%8�����g��P9�ѵ
����21f��IҚ]K�����Q�9���3gz�V���!��B�����.��M��\���tS�(�ܹsEX����qQ^V�����a{^ed�n�q�F������Qi��
]�3մ�Б�T:Xcؠ�1w��&	�����}N��˾�����;t�ŧ������l��'���D���RaŅ�����;�Y�5�D� z�����n�ss,Xdq�VwSP[N��GV�����}��'O4y�!�,6mJ�*�t�v�Y�Z<���?��ы�Uu�����`������>p�W?j�_L\:�<��*��@`��|BC�u�6��dл��?���-��0.΃paV��xV�չD�ʉ^FoҺ(��Ç����:�p`-�Y��f�~1QKKk��uz�u�Oy�K��N`nS���mu֠wR����sM�;�+�~.A�@������k~DvV:���_y>�}ac�F�Q',Ҭ�<|����Ž�ג�c9X�[W�Lv�j��J��%�JX������7� �X��ʜ"EZr$�o��ak�A#����}����k��1�Ѿ�tWqf`�������<5 k�����F��<y8���HV�K�租���+��~~�X�l	.�mB��[ؼ�$<����]�\8��vLj�����2(���ē�n�#H; �A���0,�zz�@���hZ���D�1�V$��j�^蒼�D�&b��_E8!?�N�% �I�35Z�]&")\!�r�R���^����<DFW!##�����:�E�'�̦9c�7�hJ�
"�IL�X����&�2����=���wm°�3��\�4������^Kǂ@=V���gjTgV��"��	bRtR(�hg�-[�3��朜�[
ݻ?D�7
J��j�������tl�����M�;w��E�3�s0����v�S>���갟\aAf�Lp������r���Na��Ld�G��?��ǐ�q������1��oM��XF�ѝ����嬨�ÿ�j\��"�s�2Ro��
ŧ���K�:wKJ�-�g�Oc��`ؾ}�e�$����ni�M�RN�8w�'�}��,Cd͖0��-]�C{�E����}�<��q8�u�WN ���f�q&es�Vl��"<^-z-k.�%�/`��;Cg�n"!�8M�uv����P���H�+"
�����Hi������L�ũ��`������ɞMܚ���z�Rq��,�Ĥ$"f6��o;���8����B?s���[��L?�MNT=���3��j[�bǈ�4.�X���^��Y�"��u� �Ͳ�`j]C�1�Mp&���7bSt�߱��6"���o��߈�� �hO�v-A� ����کK��L�P~�y�h�������
�y��z�w�!�U���8[#??gO�,����r�\����IL,����|�;O7������x��8�߿�j���oQw�ڍ�I[�0�r�?&NiI>����G ,���OvN!r�k�Nᷴ�4n��Ҹ˪�rl f�C��ˆ?���c�y�1 ̻�r� �%T�崜 �o�i�F��5L|F��d�^�t�]6;��� e����5Љ�wM�tv������;�tD#'�Z�F�਴鳝���kG:�!�+3+G�1�4��dt5��~�����g��X����y��r�￣|�t�"�F�� m�PN��}��;``PO\�tQ=��('�\AD9/���YI-��/zxJ�[�>������5����>M�^EV��8p(ףb!����3�)�^!0��1�.����1ަ?Vq�ǈG��b��4"J�A���0�
��xG?�{��l�{��m�`E�e��,),hy(����C��-��<�&7q�1�7��˱1�k�}k����C�6�ڽ{N��7I�5i�M���D
}+�r�[������DjJ�)4�6O�h R�I�aL��D'���\l�+��C�'��M�x��{}`ǰ)���FfL}6�pPy��,��g/!�V����{�"�[w2����D�5r���!��䂢��TT'��t��!#��K՟osb��B�.�p�r�ЭF��	��_�Y�*dex�sw��Y:X��!��P�x��*{��5|h���#TJ[=2�N�!�v"��]������ѓ�����r��9�RR�E�y�7�1!�.\9O�l;�^�s�N
��������DFj"J�3��J��D�x;��C&��r��vj� |��7�-^��۷Ȧ���#~4����+���T�P_4�0YG�4���L��"s���M�����Ů#E\�V�>�(�n�{`�Sc�w����u��w �S�H�-�!���N)�i�c���k,M���	����kK���'���4g��w6������)��� ����BhmX>5���S��b�;�r��S����S��&6"�L�R]���[�
�Z�[1&[���,���L��"�I;�tU")��r��ߥ-8��I	�%��߫��� m
J�Ը�r|��7���SQ��0ş�1�Ԩq3.w�
�@�����OH)�ъ�".!��1��|
y�4�p���Ӹm	-"o>�#XY[Ӕ���
�2��4��]��4y?�P6Z����?G���A��#\�����q��0u�4<��q`'1�J�;#GǴi�`��vN^�719��D��p�B��"a�D�����)C�lǖ!g �s�ZC��=��;	��_}`�K'�}n�_?��G�\\��k�j����!?.Qd#�i�����Gh1k�,��{�XV[�K(�J�DyҌT�Ji02��hK��t��E eӜ���9F���޽����� ��7n��H��T��`8Җ���BB<l,|}�����I����k�t�p�d�����y���;d!)�R�`o�1��Z��-߈C�		��r[��1u�:�Gѯ_?����Z��Ė�O�#�l���9��/gϞ����}$((��O@�/��'�!+�j�V�;��^-1��tvV�wuU)τ�@����͙3�����6J>�����c��ܙ�8�Sk*'��)`��~�9�=������֋#�|�� B�/ylD/�J=q��-�������G7v�"�#��u���|"�gw�܆�T�sg�!5���73��_���B����pY��H��t�DTYi{�G��e ��52A��Z������`�o00ЗĪ<��B3���4����^T���\��dQ�������_��ocqdcg%ȳc��J�Ytp�Vv�Z;N.�&��g�*<M����&\��|�^ః�Τ�0\�&�du`��C�1~L���_W$��{�a�#=��3�@��G�.;�M[�����Μ1��V��Uq�
��6X����"�c��ړ��dxT�R5>�a|��`�陙����Gwc�VJ$Β���$��	ǡc��`�(--���V�@Z��Hׅr������*���8})���Db�PG�����锯�^�2��͕���CJt���i2ǟ�\��SZ����}�����������$��4�o���gG�g}YT\6]��'�6���o$���8�5�����eqqi�Z����3:�{,x�Ѿ�e�	1��G� �ϝ#���'��oee�v���6KV��z-ݻ�`��\�Py��=rx-iA��w�E����-���~�9s�=�����;��`_k�����/
���W�.7��[ύ��E��Q����OsZaj�!�t�]����Zb0��x=6��.rr�8�q��L1��� �^]j�\�����ϒ���iY�M�ׇ���فZ$����Q������C�Q)m��dOr_��L!�>����Z����Llv?�ZMe��}7��e3��
y
o�����*[���<X2��? B��ECʧ�ڙ���wiAXe�E�]���t�\S�cuϿ���>��,j�0�Ң����N#��j���q��D]��!D)W�ћs�C.oRw����4��!�Ƹ�Kq��}��5=)��z���pcQX���Lϔ�k�U��f.#q��N��,�e_�uT�Zs�ː#L���[-[8Վ�7�8��j'�󭬩fDD�8�'1q�I����Ի�{�����\9�KlDI`����1�G&jB:fŘ�ѵuB��	"�t��C��A>z�Z��s�r�˘��'ёk@�Ƨqa9����%��w���@ԭd�e�V�**�\#��D��
��.^�}��܏�S$&��\B����R�sws�8�-������r'��u%��,,��\����q�L�a=8�{-����*+"��yE�2����x��()I����;�
���	7o���fb�rW�����R�%
�f��AX}�p�,3<,�)x`RRN�L۱ee#�6G8�&�P�f^�Ģ�Hfv�O���O`ǯ�Z5)�"1a��m�m�2�ҵ��E9A��터�:xN'kf:�-��5U��F�������^̜�2}S�]��E�-����n��W,k����&�N{Z�p�<|�*�����n��~ǒ�Ǳ���e��a$��'&��/�Y��BG���O6���۷o���Sq�)]�T�Pl#ny�Vrm���b+b�Y�=�3�r`��KXC-���Α]�<�;�`cRrV�p�����֖5�ĝu-6|X5�t�		L��Č���y�������2Dbvk����lXX� ##��`���))�Un��"~���t����X�B��F��%���;8 �����@�՘R_�V�'�\��r޼�e�*.kkmm���]5��eb���%��H�XA�ዢL���o�ތȨ�`�c��)n�&��l5�%�c����Ll�.���B�_��D�XZ��ɜeb�F$a��`�ʕ�)#<.�m�������k֮]C�{8�7�4kR���¬�(�L�/%�@R~~�H̝3�A����,���� `G��2�� ��~.W,�B���q*��y�U�Kc��tf�~����sQ\Hك���#���/
)Ozi�(�\s�fn���M�N�R�ۻw￸N�{���8.5�%J�Ka��Q=�E<hʋ���8#��k11؄��.F"�ﶖ \����Ό����=Z��z����_���s�W��{��S]j����u@qI)��y�P�����5�WpqQ�Mh�?�1����z��[��ҕ4��?O$00Pl���t�|_u�8��ˇ>9�˄fo��l��HnK //�?�H,�޽����SD�oG_��׋2���J1~_�h�?���HH��@�aT��IIQF�O?�$�ɇ,��PJ���AF6*X�qi@F��0qd!��������?[��U�?��oE%B    IEND�B`�PK   �`EX4�Z�ȅ  �  /   images/7751e6dc-0a88-457d-995b-e2164771e840.png ^@���PNG

   IHDR   �  �   ��   	pHYs  %  %IR$�  ��IDATx��g�\�u&��z	9@ ��$R�HQɒ,QVζ��cY�GvO��5�cfyu�{���z��V�gdIv�%9Hv+��%1�9�@"x�����s�{wݺ���l�^ݺ���t�ާZK�T
���?�H�R4������4��H�8�u�ߤ4Mu�1�
U+�z���g�߻�d^� uA�$M���T����vH��]�/ns�9J� �ܤH�X�m9�{�4�F�:�� r���������R��do���}������'4>>.
l�W��;�u�����`�y�9�Q�P�@A���a��F�V�x2��KZV��\�T���D��N�ҩ���z�8(� ��䤼��r��Q= �o���.�L�-[&###�ȹ@U7nZvzx�
��	hdm�:FZ]�!����4��b��V���-Z���A�^Fl(��G��z�j5�ߏ;&{���Çell,Ae`�q�ׯ�M�6�bŊ,��T�:۲3�~t�9&�NS�H�`it Ϊ�#t:&X��ҧ���V�W*�<�z��CCC��N���'Oʑ#G�����~	D@b�Z|��X�����^9�|�jMj�{]�Vӊ�I��¨L#�t��)�`$E�)�t%r�N��@g���k�N��)&����q�'WصkW�I  ���pl��ı'N��8�ڵke�ʕ�t�R�B�,ը�
�ȱ�����
�"P�ܭ����q�H�S�*�TTE����ȱ��V�N&8:r饗��ŋ��1�b�u�������{��^xA����:��v:���� �m j�=::�kd��X��?��vh��~��
���R�t���L����W�T����7	�tb��@h���ؾ}��(�� v0�u� r�@�Ql?~\��+��"�=���޽[��wN`�i�� $ 
���y��8����P�*'�Jv�N�;�R��"K��i�2>6*��=>vJ���O����� @b��@WUҨ��A#�������3Ő�A��RF8�Z9<\ ��桇R��J,���z�9�|��:�
��b��k,_�\��R4�U����쎥ި��ގ]å�/M����9�2>*�d�T݋�㳑v�(�H����&�;����BD�����K��3�(P���p?t(�I��dG���;� l8� �*��,4����e'L�ɤ*�)�Ru�:4(I%�1��=)'&'r�l�ڱ�JÀE����N�L��α܄:B�@��E��O<��:	�u
�:�h>S��V�X��o�j�*Y�f�,Y�dae��GKvC�tpP/KW$p�˘�c�I9՘���)sn_�_w �9S��6��8e��١�q�p��m��݊>�"����(>�f�#�<">��<��Ӫ��kQ��9�.�Al�3������ǃ����|'p�Y ޠ$��\����qA6���%�hى�p|%u�#͍P��S�����r��`���<�#�)�I'��C ���5��t J�D\���,�t zX�p�������&�9�A��� 7ظq���O������q-�,�`�_ �k���QuxhQ�n���Qԗ�:X8�8�T�Jn8 ����'j2�����+* �&
�J#����=�Z%VY����	����Snq��K�Ê�� �������9�����Q�p �5�	��RupxI�N}��p�<�wε���q@I�hL*N89y�@2�q�q�A=���رT6}_��>k��3�A0y��>ݠ�Bd�[�*�"��!H��߰a�~, :���eEPW���@����Iy�'��5�g����So)�:u�ɱ�欠��L��߱E @��E��8���8��4a�'�|Rv��!�?���n�s�z$t���P ��M\J*����ܰ��`����X�')�U_:v�d�c��Zx)�8��57�]�&9:唷���Fө���N8�^�J��v ��d� t<:
�~�;�r�I@+�,N��|*аP�9��$��7����Sq�� ����p�I� ��\E19/�2�jE�n��%�t�5�1ꈫI26*��L��Ny�R�Ǎ*��(�\�i�О:q��<�����߹s��I~���>��c���Dr��9Ȗ-[䢋.RK�,�kx \	��υ`��L�B��~�"P�#U��ٟ-��:9�b�	�Ę�H��;���'�������;dljRj�4V��Vr%��ƱA�$�51��^��G}T^|�E�,;�q���� ����e۶m�4t�[�FB�c`�`(b ��װ�7_�z�/�R��ĤN|(14Z�'\c��W�������Gd�XM}'Z=$2�+{��ֆ&����Q�@/A�P_�\���Q�9(��G6oެ��l�Z������7n��j�Q��|�j�x�d��C��A�������^r���Ծ�q�N�u
\ŋl�ݤ���bMV6"�N�pγ�ąe��s�=r�w��E��(��� �7� W^y��#+64�3��N�+��폍`���T{4�y\Q���N�j}�(���㬡"�8޹�d���R�$a�m��F�Q�m�N���h���ѝ��
�bb�8AY������ٺu��#�"�.vǊ�b���*��0NƬXnD����TMʒ��>���R'�`"k�M�q[����H�AbtL�����I;��le��n�g�}V����T\���$�K �׽�u��@?�BK<;֊	�|t�3$��$8p8=��9h�3��G���{�E��I�.�~8�gb !��
b����T'��܊��E1���ȁ��k@�u�쟳���ҙF�
+B FV�^��_�!�7>qoF�[ˋb��1��}������Q�tm	⦑hВ�$�z�#M;0��M�.S��CpZ ;�Cn�(�j�	Ƥ��@��eGb?�f�n�`h췊+���d��+��j�sA��y
�j]�!�P$WJ�"�(t��A���1!�)J=�H��_Q�,2;�[$48F2@p��
�	�W8cW��	8	@����UK:І+�ok�P�q�@�q"�~�y�Z�n�&��PA(c^چ���D�o���ĸ�"!����vBJ1�:{װ���E� 8	��Pfq�zK=o����� j�0�m�F�^�w��܃�Ƣ�܄\Q9_T�o�-;U'���>cp��֐E��|�r����cO>.�u\��AU#��n��«3�E�9��H��	��	�B���;`$�8>(���؁���E]���I$���F.BNb���J��J�������e�
��S���P\U�4dd ��ԍ�Cr���z���ToR��S�|��Z��D+�!���Cs��_�� g��ux��M�Q�E8�'ҹJAd;��=(���>�b+�P����Zv��@�X)ba'M�'2M$�e�?V��pHJ���\���o:�`�������u�]j ���	���Q�lha�f�k_�Z; M/)<�D�h�F�W���Aִ���{�(	~C�7�u�������vY�5u�z�C��EC�+ ,p���������x��^��a��-Q��G�3���t#�մ���гK���"Ϛ���3˖�b[e�^���� g�K0��L�+S=�9�&��WL��¡��c����W ���_��;�t�u��dT8>q-N)X� ]��_��e�HV��w@A�G��&�)�� r.��60���~b_9Z��vb�@� gD6pr�bxB'b'(��:t(�F�W֊r�k�������*�Ëd�D V˟)�� 6�5B��JE�*��W`��@/�~B��'}���mL.�%��!�_t��O� �A/bz)�*��zJ����*���Ŭu��3���5�+�e��A`4H�%,�f'�z ��%�\��� ��:�!�� �ݠT��pR�܌���� 
��-9��-G)��덤X�	���>\��*�'��`�����  �]w�b���X��v@
]	��@������X�n� �yONX̅�V�\��/��/��P�C���#���o�N="G�ȅ	
��>�u�S)%7��+�5�y�� T�.��9<��A 	,/<6:�l:)E �epwCB_�o���G�J��K�nh����h�;�㌁���l�#r�X������V��v�k�(�'��7��^vn�X{�*�8��V�� ��.�b=E�z;�\��:��3��R�D���OƝb����5���oT�H6਌ze�<��``x%�����Qx�����Y�AW� O���\��?���	��
	����L0>�6S�:����Ԁ�.��)m�����xNXc�ݦB=m���������щ�	't�RA�0�����@W��E}���_��n��@w�����r�D��mS"�� ��UW]���?MfpF��)�Z�¨�(�͚�v�����"P�3�(d�t��#RHs3�t�C?A'�/�������ϔT�>$;�a��P|<3Eh7j>P߁R�
#�,�-��� -��; � pۃ��t���E���M!�����d��w�X߂��c`4La�`�oO�v�LV�fQ�(�qf�.���,'a!��0W�֤�>��&��������0���0�X�?�09=�Ѷ�(i(do�%6�����`�2ByH��ّ39Z�Ѡ� &��r\��4k��9�av�=���J���������`J�U��ԨM��WOHc`��̜&y���#��<�: �Ɩ2>�`����������>t(�ǿ�K6��D<�����T���0�~� lx��lF���)7�P���������IkX�*q5�'446������ˡ�_��)�[:$������_�F�n�8�+��.l8[bz	�$�$�O �l�Z�w��)"�,�t��a$�v.����:�}��
P��?޺S5��5�t�Į�P7�>%'�#{_��ZC�{�lP�T�h(�LJg�c]� �`5�뺵M��� t<�@b���>9Q1�ߙ��n�u�SuJV����ɘĎS�D%h$)���KT�":~�! ;A�jԇ�8J���9]�N@ccD^���7�A�4�����,�ŜN Ys�F���C�	 ����H�u/m�	=�19.��K��j(�ak28�<�I���щ�%�{���>�]�z�Q|��:G%]� ǵ�^�N5��3	���=zVa�0N�����I��#�IL ��d!R5����T+�e b�q�zq��%U_��:� �FUi�X���ַ&�v��f�� c^a� ϔ�loY@�	Cm����w�� (��~�^;ղM8Pː �0pf���JL�4ۢ�I�|������\��
N5ľ��:��$��\�	��F��	lv�9ʂ=��JvG�7��m�I�1��:24����0N�8���-Ԁd�%P< GX���(4K�:3�s��={M�����g�P1+�~��22��v=V���b�,8��DOZwVO"�Ȣ������`�	��:��)U��W� �.�>hp(��"=9 D��g���,aNO�����vY�-ƭ,T���Ҳ�h��P'֍�a5��˖ȱ�dǝ���3�6&n�Í����=��R�%D;=��x_����a�̙Vd������� �������i2㓞W�߃��{0��ₔ�/���J�;ݤ�p�;�@��!zdղ�rh�+�e�|��p�8��������5��ށl��e۳ᘲyB�t�Ǌ�'�9��g`�|��텪�l(�3�$s�Y��q2hJMƊ,�E�Jٳn��D1u��%D���C�'�@����6�N��Zbx&����!��RuI\�v�j8�lh�yM�?&j�ɔ�4no%�a	�P��h��>�N�C����|�u��<��\�b�B@!_�"�T�K�3��] ��#?�W����4j�~�0L �N"�e�:J���E�@��a@1��f�s�c�K��d�dw��/|'��+��a�U�M8y>>�}+����ޖ��E��E�5��"Tl�*�
�h#G�:�MY��� P �ƜY^�T��H�ˋ�Եw2.��[BW�N¸� ��n��uI���Xf��8� [C����`j�GӞ�g���B�J���6��x�j@qb(�בa̒.Rn�!���-VH��s��bl��Į�A��,u���^�z*<g!�c�KvGZ�8����@	�g�����Q���Z���>��Ų�����Vm�:ne���hl��V� 8h�0RT����p�% ˄ٲ��I�r�N�
��Ԣ�(�H�X�'��p���;.��I��":����<_�k 6(�ލ8��	��,�a������)`�>:�@���a�#�{p�$�c�d ��P-������'H&]����|�LN!t`P�'Wʑ#G�著\���bo��C�yj����ӭ�`Mef5Zg�|��DգGw���k&uT�t���Ī�LL�����Z9v�;����xPV=@�X%���:��;w��,q~�W.fCX��
�s�t7�V+���;Y�%W@<�U!Y��%w��	����"ĝ��
�8�%�#k.zݤy�sծ^�B�.1Ċ�6�h!Ru�ֲp�5"�!�XLΡB"b3b���XC������w�J:�NJ����0�.�&뚷��	�t2�BkzW#GY�T]���ĹJ�2)�JM�XV�uve>�!�ˢŎ�,+�I��+��+�*X�*[	d�ҋna��Q�������[Ȇ�5A@O��*���z*�,\�o�"Naq��/�A#�{)v$�f�Z���Z��`�2>ZR0�e���ű��x��d�s;�PC�F�2zj
�&D��5�S�(�ju��u�fUh���̲얝5^�:ʱ��TG��JREh��Vݨ��v�4W��ccnsJn2�DV�X���j9�D]��pB��
�I�6Q4���n�#!v��\��b}(6��}�)Ȃ9�m�F�U���e��S���ɀ��k��l�d��ǥ���b�iD'yP#?�y���j:i��L�z�\KC��̼��b�(HF�u�,Ph	Y3Љ��(�m�e��ה�t���@GV%��R�r\&q#��T&V���R�>�g
����r����T�8�`�Ċ��V��
�>�q��4���mӭa;_��x�%�cI�CNaT˦RAj�>REicT.�R����u�����|�����IE��v@ ���0�������g(,�l9G7��.��ߊ�X(T�JRJ5=���q����B��o�V�������}Z�u�� $(�$���p�RB�2C��M���,<�N��١yӉ!�x�i�k��z�jC���Lտ�X�Ө$>�f���rѶ+��d�c�8JM��1����̚#v�
��`��L6��H�W��z�(TZ��-6�P�q�V��ܜ���R�q��h�2��^���͠0�:ꡠVN���ņG��̀ r�nD�Q���� �J�R$`d*����,��F���Zq
h]h�x�8J]���0t��u��Yl�ֳ��^��@ SG��ɂ�(e;��iZ�JKɀ�Gi�X�ҙ��$q�Xr]YX/��/�t�{�-��֌�l����}!R�����]<�,�j�b� ���5[������II��|�@B`�������T(Dt[G�.[K���mt�!`�I���=�l	u���{,gN3���d.V�����bX1f�
-u,�̾iᦶ�%���2n�P��@�&ْ��gRF�2M��{��J���c9O�"���·��=�	T,�S��H�2M�@Y�!�J�,P8�D�<�7�`���2g[t^G��D��Qԓź�\��v}b��:'(1/�dv,0�y��l%U;��P�J;*:⺑u��;����J�3��-Q,����J�[�E߫~a'�e�����fu�nD=ǚ��9`���@)�&�� ��qq�݅L�PlL+�O$��~r��9���t��$՗r����:
�J�\��y>E@P�a]�b�l�z�|�s
(t��qG�4�+�
��3� m&#�lJ�9B�:�ȱ�����t�
�F����@61�<��9�M��C��}���L�9�j����s��tN��	@B� 
���y���s(T^�=�E ��<���t� D��b9�B�;S�`�²���x��º<�>��<���K�J�H8�5�j��|Ƶ ���8�,Bp(�Y-���(��m�?���ڵKKrq�Zt6K�vA 
RQq-�u�S_��`�R�*`k��7��#G��޽{� ��Ž���7�-<��Z�c˖-ʙ��i� �DS׆�P��g��_|Q9��� K_��p,}���.�2����D�5 )
 R�E��1��Cg[nҫ/b
J�}��x�6˗/W�Ž�s�y@�l�� H�9 �$�M8��� ����5�*���	=�k
b!ʅ�YP���=�:󩧞R� aA��b-�Nd�rXP 	~۶m����h� d����0��~�i���4�U���
W� �xz= ��=pM\�V�>�9L��t"�D�c�=��(S�ֱ��P��F8�˯ \Xj�1�eÆ�i� ���� �b7�Sй9���t��Kk'��B?Cp=l�&|�d�ƍ*�E�g���`�RY��#֊AJv%�b0�J1(ۦz�����e4_cjP8�ϕ2�M(�r�I�u$�ZP@i��<W9sZ0@)�y�1��`�*Fݟ��ӂ�yP�,-(���V�kn�5�ˮ]LG�f���B�;��b�}��嶀��p�T�s�βs��:Pz�gz�^���
L݈K�rr��WƥWY(tVߪ���^t�^Xz/�񢯥,��q���t��%y"�U��%z��u�Q��.r{�t�bŔ��a�H�'-DZ�|���E�O�����Ʊ� �e!Ҝ J/�`&�$ k!u#.��$wZXV-D껎ҋ�ы쟮�RVϭ"�8�L���������:P���^�ԭ^~�tծ�c�<W��9����%�t��"�
���uW!��ŕ�� ��x���2�����kw"t�<{�?"@	��F 4�iKrq�8��M3���`$�~�wA`��a�Bn[V�iGv-�v�6%����ݦ��~�U��
�u�`��� ��κ# B�X�Ye����ظC��u�	�~��P��٣�� �	!� DW@�3�,���#8p��XY�p�\���ȍ�8�vj�&-;�Q*Zkv�}XO�k��	��L�N��Hm��/B s{9�@� :93Hc@)��}hP�F(v�t�.#\`��
��3��'We63�~8璣���> ��Ax'����Q��k�NTV�����vx7rJl���h�bqB���KzI[�XW6G�� o�B\*�E���t:�r�F�5~���,+�lU%�G�s�v4"�5(:y+v�>�T�`�Np���NT��n��'�\��V����s�����X	�k���ȷ�U��ʦ�F�+��"�?��n 8	Fuk6��2�u�vǰ�9Í@�s��F�8�6�\���KRI'�粶��0�>v���U'(�G��T�xe�� ދ@x׮]��<+�1�醎G#�m"8����;wjr�zt��H�������D��Q�ޏ����o8�\�}��6��*�|^��b=Y���(�;q��� ���5�y�0��)����l��������Z�ZQ9P��'?Qq�"��ɓM�̚��N�m�^]ݎ˧bGE�����~4�q�#W��N,}$�6|7vR��"��Y�ɽ�{Y��KV!���p�xWxw��n3���m�bA�Ca4"�\���:!�*���R G<�ի�.6Z�ߩK����B���n�g�1xn[F�*�,,DL����E�1��8�����]�mF�n�y�8%@p��(v��֭*�zK[�;�r��:	��JѲ`v_�XZ�&j�����?�<�y.�ex?�.���7v2Mi��9]6�:��n�[v�{VG�ov���/��:@_�6bu�}P�	�w�}��q����w�
E���� '�X>�zBy�n�֍��tlZ��Y�9�8)�1#d����s�5��]���g)�������Y�\x�
kPe��Ȝy��؉�8�YcB'n�Ei��|+lG�d��n\����^�[/>�^�f"��m[\C���rq�� j����b���ꙵe� xi5X� ��$z\��2�ɸ^��r�^��K�c7�Ý)ZJ���p,�W�W�iJ��K�����(Xgd��ݙ/h��p�S�Vi�uѫ��+��-z����^Di���NT� � Z~���gHX�8\��4��������Y"����	݃ �F�� ���e�m��˙�L��nϙ= ;���� ��;�+,��%�\�\�������h
a�B?��
D�Z7�L�^I�n4��2e#�L����n����'��k�B����Ve�'8>�:�^�@��	�&u5����$H <�A��#;�^
���?�~�6�{y����x���b{�95h��c��M�,�D���]��K@��bA z0� bPŭ8�1�e&�^D�Lܧ�%%?-W���A��K��~;!Jˉ����b��F��7�a������g8z�LL�zu��	͔2k�*ks�U�%P�6���ݘ�]��	��q~��������t�kkKu��3�����Lcg@3e[}ā�k�
��� jCp<�
j^�n�ZA��g5���A��D ��>Sb�<�����E�>��O��⌁BT�[����?*E˳ײ�3��d�6��8Og�����4�Ќ�����y�Y������=�yZ�tF@iT3����tv��_�:�sF@��67�~(��� ��bLM7�
���t��+s��s��N"�ҝ~ՕW��_�Y�r��'��oP�{D��,ZRxaV=
�8M���I8
�'���_�]�	�2`h̊�tT���5��4ϰ+R�]�Qw�l�zM<K�����'=��=�S3���<o��T�OM�g�+�,Ǐ���/�(����5�m��b�V�oc�u
^N3��"p���X�-UUV��.]�L~�K�.7��&m�Z���!�)E��x�*P$ֆl"��H��(8J��L2 �hR���)k�4 *@�ĕ��9+���LO�&j� ��Q�~�6M�v G%�\KexdX�9*���_�:Ӷ�uh�ڹ�mV!ߟ�A}/{�O~ҁ�rĽ���'�� 7�(��hL�!�-���M����
S�����L���B�z��ԍ��A �!\����w^�R����zFڑy�Y{Τ@q/�8.�c4�ħ�V*���B߁r�7Ȟ=������gċ�ꀲo6-GE7�*F�?�3�i�(tr\I$5�S�w�끐T�w�Ԩp��i���K)�)3
��*�R=��}5��C��P{�g7~6��@�|ґ#�e��29QsQul�*9Q��B�<m�N8��S�O9@U�$�f�����Q'�x+��t��{�J8�U�D��ͻ")���Oe���'q��������]]��9���9��	p���tmRQ��H�^nKE��J�t�"q�M@��i3��1�:r3�J���D�UX�I86��)�W��pF�AZ8�ީ�����I�x�g�	P'N�p��(�[�=h�gXq�$a-T���c�Y��<�iIQ\���̎O����R�]���6�T��gT܄W�T� 7���7LT��[*�|#����32C�b��ji�f��Sy�K������M�xR�ڣ�]
e0�GF�=mJ	l=V�P8,�6�Oxv��e�T@�A,���~�1�s(LI��$+���N�q�L����Ư7BӤ��^)3aE2�7
fT�n��#Fm~+�ٯӄx8?I�=�0K�on'd�9y��-�8RܔSm��� ��1�t�qRO
@9�I@۪���]$�)�:JE�Z=\�:��o�c,%�
Jf�,�馊�ߧ\��IZ����ۦ���W�G���m$-. z�U������l���K��m���G*Af�u�4{� ��uf���;�-�is�2������,E=�9[���!M���Ӽ��zG�Y�3��R�DѬtW�(����?Pļl�Z-����<\q�(i�C�����:&.s��RGY1��^SPf������z'�}��r�F~��M��z��3"����.��7���^�3�E���s6���$S��g��դ%�#����V��]O�w�}�a�T��Ȕ�&o/��=Is�z2kU4��JP�S�tL_p���)*γA}J��n��H�$�x�1�����8*��ӆ��Svn��]S��u�4��Jj
�i�*/�����Z��l�DAGh�*��i�S�����}F��}2+�((��lwVOd�*mv�Y[��4�@�4sEs����45��L鮋��)�RR��A��PY.�5OD�<�c�Θ����D�LWayx[|�u�z���Ùh.~/�\3/�o�GDGG�-�"iڈ=+nK���TN��{�ǋ���36�;`kxO�9�<g��P���+S7�*yo<դğ!�g-���s@�p#�b@���e��<|��ƪ	�ii#�-J��7u��n��xڈ��QPT�wÝ�Ld�,����&\'N�,t�ה�R	a�i��*Sf�柚|
�Cs (��F�e�� f' ��/i,�q4J��\;W�_d�q��RQ�����F0i�sd�k���5�V������3�|bfi^�cR�,jhӆ�����w�od�ۂ/�����H2	W���>'��y��XW��T���/�c��󚹘�5��Pl�DVg.M�Op�U������E��c+�y�M�!`#�[�.=��W55�ސzcR�E�jE9Y�P�4�$����(< *=p�٦9 ��®�UҤ$u?ҡ���z��ի����	�A>j�%��VY�ǁ�����Mj�!�U|0KZ���i�OS�4�RI�R����e�䘜8zL�,^�q�SS�r��h��x�,	��d(�J�
(�B����'����a��Eu@m�/�V�^�XV�Z-+׬�)A1�����(:I|:D��i R�?&�>��8pP�,���H^=x�r�����e��M����"	Qs��zgZ$y$��l�2-@�g_���^�\>���ʳ�>+�?���ᦛd��u2� ��� ��+KG�l����zڅ���ڴ���� ��L��v^B\��4��RK��{��/</�֮�%K�j�J�=��m��$�׭1�ű睐z�G}�(�Y����)�y��=&۶^�i^=(���ge��2��>�#����5֊������=��#�ȇd��]�կ��>rDv��[>��OȪի}Y,���ӥ_�7*3u��D\Y�'�#P���2[ �(as��|��)N�sL��r0͚6	ky��>=���ˬ<���r�J����,u��䩓r���ˮw��M�Ej卓ҲQ	���2>�W��G>�������2�Z�w���w�%_��_���,[�Ȥ;!e��ݲc��o��7��z�>�y���+�ӟ���������e�������6i�VQ��6��^V˿/�Gˈz&v��=
�"gX})�A�h_���V��ڀH=�uV�Y��:40�M.��M	ϭ�A�*'��6n���)��+_��zD�juw�5M�#�
-�ȗ�����������[�����_��:|H��������=�Q�:P�C�s�oFf��`���"�]G�d���c9�l�|hcB&��']cE(�_���i=U'�.��r]wxtlT�Tn�<���t��QǪ�u�����Ik����nsf����[u��`�����x�F�;�(.R���C��~D���FF�����R�~�cy���/.� X����)�˞���3�N~��w�(K����nS�%�մRzB}� ��>+d��v4:�sM�$��E#^\e�O��Oc�ܴe�Ҫ&g{\�ŗ^�]/�� 3� �>���+X6�1�i�Tl>+9��^$xb��Yu������A6]p��;��瞓v�w���M ��TCM����&S�����O��9ٶ}
;Sh�A�t~�a�R�(���òw�^]�l钥�h�"�0�O��r�����U�����;�x�E|&w�u��E4>vJV,[���ݿ��r�nq"�2�uJ����Ntz3
y�q�a:,*���N�=rH9���>��#�t�R�w��U�dk ���)k�Qe�Ps(07��Y0�~�zY=��Y�:�Ճ��9�w��\c�U/S��lf��Lz�[�:7�<��s�]�P���j�?����r�?����x�Wɖ-[erl���xd��Sw��İ��^�N��?��$��r�����G�O�˒�Ke��{��M���ˎ��w�jdsCz�Y4��lJ�R���1QZ�@u:��v}�[>zL���#A�)8�t:<�5>�Q�y3��M�e3���}_3������)�p�:|D�,�-[��(�U�L��dr&��7�Vv�����21>!K�8q3&S����$���i�T����2�;P�ల,%��Q�=b}3�֯�j��>��a5T�!�E���E[�(Pt��0/�%f
_��AIEŧ)wp����q�!9~�Ӄ6ʇ>�a]�d,p�l��q0�9���B��!_��ߓ-nr��	�����u��s�<>P�\K���M��Ql5["�E�{�l�7q>��!V#Fa�4���Aa��௉�0�4!mJ֯]#�<�,���Q���Ĳz%�^���7a�L�D�����&���0u˗.����-r�UW�����9�H�_���$��>I�N��d3XF �o�d����/e׮���}X[�b�zz��dtbR�������x�`ԦH�g��bJh�ل}�A�7�/ʖ��q��m!~f�}�Ǐ�2���RW��,;��씏����D����Îs�r�0�vȀ3�O�8!��}E.�~�N�)C
�p�Ŗ���$O>��.��frrB�,rS�͍7�Au�(���i3�4W��56>�f����LM�en�G�EtB��*�I��lϲ8���̘�l���@��& ����yA"�hSXԻ���]���G���i��S5A�C`z:pP^x���X���&,�k�nu����1�ADDm&P��U�/�Z�R�����^_��]��L�tټ 8]1� � ����G��?����:��c��a��lظQ;�-���D�l��,R��8�U�ˉ���V�8��j����q7B��N�<���ױS�WP�ɑ7�˸ ��ZCV;3��)'����G,�=����Օօ\���`��:հ"�׻�Ο��2�b�J�.��[��6g&/Ϧ9�Q3�z�,��%��1$S`s��S#,-�_�F�&7!"pȐvJE�9�1z'����2� 5O���yE����TE�����>ׁ�����b]����IΖWQ.��Q�,�~���x�Ε��0S�a���XgIQ�զ*?!�r����� � �ġd&��=ZZtjB�.^��#M�z@�\s�LNՔ�T��[sJj%L�A�a^#(�0Q�=&�_q���M���ɰ�Vd}��'5� >���E���i��H>�ԃ�%K� �� �S��4�4%S�|�gEL��$���a�2{i��E�`̶I�p���ELǱcGUIL���K8N����'ZG�z�F��ː¤<��	L��,[�TFGOɦ͛u����xy�q	՜�Z�hD��n��O��'�_�U�ٮ��ZY�D��KM�sr.E�K�����y�Ɏ;�\��b9|��sf���x�v��jJ���c,ʢ�*���_�-?���S�g��z}XR5w,���O|RC�Z�W�.380�����?˾}{UQ�:α�u��l}eS]]�$� ���/����Np	�����܂KЋ����>y�jj�f�?p��սzu��0�kxkj�p�.p���B��p�s����Sս[�!q3�b���� ���s�p�1
8�h��mr�1�Q5�����Wd�CAa�C��z�X��G�����V*U5{�J�A��[����r��r���L��;�5�9��6yX��k)V�IS���]&
����R4�� �Nz�$�lY�ov{�/M�D�MC1�"0M+a�,�
�k�s���|�����Ş|
�[��*ڄV~w��Mp����\=2[4NY�/��B��Z3y�ώ�����
�5K�K&4_fOIB��8�<�/+6��M��z��W���u�x�:�y)�KV}Ȱ�)���Vv���_z�K��c�]����F{߭Cc�$!B�!ъƱT�_��Y�GԕH�|Q�Ud���/Y�t*�V)N��(�2��U뫥�*��P��8�2h�ȳj��`��7����	���>�@��By��i]��r�z��<t<���ƥ���)�Sβm��e9�'���/�R�/wSW���ibR��7�$φ����5%rljV8By�2Y�>��u-8S�����4�I6(�1�G��\�������Q�6�US�v�2,�� �nǚH��n�qMoo�K>�چ}��57_���� 7M_�Lt<b��O���	�\�5z^��T�g+�B�.�u!�:�%�C��*,B=��H(S�h1�b �jh�=#dO�)�j������o�\5RE8�,�O�r3��hyɝ�湍4��o5�\o�O�9��"h��Q7v��h�|�Xg����9&m~4����#�)^�;iw ��oլc
Y�(��ح �KN�u�bJ/�b>�O-�豝�XS�h��ȷ�YP��.��V4�i��ƕ1�O��t�ੴw͙HdPe%\���~4}��Fam8k1=�*0��/��Q6���X�mG�?�V��nw������1zK�0�U�̖���[���J��V�a��n���u�U�*N*�uc���L����Q��C:�q�6�����T"W�"���-����;͜��y�j疲&�ւ��#�����wC_/�_��w�s�}X�V�x�+ȑ��n`�9��1cv��6�o0�T#3��q��
�f�)N�sIk�4��W"_�Qga�t�5�}K��Ł���tL�����Ё'C�.���6���m.�MN���������qp������1#A�:��Dp����hGk���,��L(�%�Nb�fRZa0G�r]�Au���>)Iy����|�`�+L�/k�n�&/��)��J�ٟ�
����|���z=~��>C�6����#��9������l��%�nؿ[��|,�r�Qx8���)B(:]��s�@ˠg��L�>�M�O�c��?���y��/��|5���Gm5��ۙ�zi?f�*�J�����(�8�E�P>~�T��(��C��ک)�*�mZ�%�7��U�J�'L>���*w�e%
�l�	Cr�퉑#��L������ν�%}*����|I� ���֔x Q5y���;�E�қ��=�|��J��6������� �x2M�p&�8�>"���T��P�{�M�� ��e�Z\�k��<��6��cu�8�СL]ws1���o�qw���6u�j�u���3�8E���)~v�f�H�;���q֯���w��և /��t�a������i
�=�s[��w�h�e�,���F��F���3O����"�� ��|EOg#����Ԑ"���X��;��S�Pk�%�m�3��Ճ?�ΧSW�n'tBΚ�t�qR�Y�aI���$���ba]��Wj'a���������D�o�	8���R-��
n;�K�7*l+"f�O����<<gS8��)$�k?S���e���;�b��G�F4OHR���P࿯4`�~3AO�j�V�!��*x��-�鰟�6p�VPR��/ߺ%�:�TϒՁ�}I��+��h�fF�����?���/K��/[��故h�?J~t{eo��O�1��V�����W������@�V�m�2��ՕX_aC�iQ��H�U�đ�P&�M�F�vYƳ���5^��]�5"O�^�7LL�E�Yg��V�U�kS�O���Aeԍ�_�攱l~r��z����f��5X��F��S�$���}K^Pϑ�@w���W�}E�<l�a�bvJ��5��g���݈&8���w[w)W�f�[� ��gK+V�b���Q���S��@�٨c�k�M}pf�i���%��So�_v�ڋH`����G������m��o��o�ST��F6�F�:�����7A(��q�j�G�v��U��9|��+��Q|��M��J��t�n���j���>��I&)�Y�]]���e���/B��q�W<�sskLZ�MuI�E�ݾ�\d_��g�}��X�&3�����Z��;�7�m���!�B����X�L2�de��L���"���U gУb�i��UϸsV���{��-��&��4^��r@��j7�/�&�f���	v�W�ߝ���˟u�?Ɩ{?����?�ÿU��U���C Z�.��\C���	`���տM]�ş{]y��}���hc0�)Z7�u�=L0��ufs�_�ч��3,�L*��[�yC���:��yTa�X>uʑJ��1<kh	�ET��;��'�$���_����=x\��E�'�(�EymU������^(�J)4#1��D����OAh�2��1ĉ�)J��Mu����u���<Z*t�����a����w!f��U���Y
i�/Hw}i[z{:/%Z�R�zB�
�4��\���	�`��� �+�����ec�Y5C��:�e(U{�ӱ[�ۉ�`��,��-�f*_�A�����{|�"�4�s�J��)��O��/m�k3�?&��%Hf�+��w=w`��+�f���R�݀@x��oa��7h��G�O�&{��)�zsm��VE*�� ��皮�� �Y�ڼS6�i�n�9<bJ���W\1���3c�U�⩵��m;"�5�Y���0L�[˭	~Ur-y�{_��v�)
�E��-�+��Z;^����n�|��aP Pkp�_ڈ)wؑi��ި�T���DC�g�g��c�5��+t�f�I�����a�8�l<[#r�׫����ݞ�{����р�����]�3:�+�w��ȢvKe���P��#�+��N�Ӕ�eBD�̞R	�x�l{��WU��¢C����R�'�w�+���ꩳ�O��垪��m��`K<\|�w ,M�!�ƿ5KR�d�E�P�j��7����Q�I$O�^�Y�9��?G�Y�X�^�x�e��������T�([����^w��`O�Ir���j{�.ڽg����tB�y�����ZZ�h��|��}��f��}+���xկ�����/d��Q��U�	obH�j$��Hv��~�U��<#�Ҟ�(���v/�,K)� d�x����c#UVF���?hq��00"]"���1���=�w�^��D�]Dď>�)�7	?ʶ�V�s����故)�zw�t���|l���,���WKz�J=�����-���;��귱���*ρ�5������}S��:?�R"�$`x�-��י{d��B Sls5BU�m��Ċ�	~��f'$�m0��ƗniҘ3��Di��CF8�p�k���;�M_�	!�G�E�|���@�g�p���i����]�jEЕm\��#t�A�U�h��k�SF]����g'n�A��sK����{Д���#��!�EƖ�cGP*�����q�B���XK�x��|��ĻA�;�d#1;�O�%�̚�f�FBէH������=�E�����I=��wB�]�<�Ä`��,LB��ڋ� ͕�c���c`L����.��ۡ1'�@[�&�]�`w��&yH�rBW����uι�ꔓE���ʠ��+:��u9�<B��o�j�ֲ�}��X��A�}+�e�����]R��bK�`�+�ciDz3鿗��G�R�� ��6�9X$箠y7�[����<?���^@���,���Z>��Q֩PO�*���w%c3MG����T�ܖ��5�V/�x�I�lIK��#Q!��CF`��S�)��?��&�C@�e�3�p?��7�H��X��Y���X��l0�N�s�����۰��Pn�|G$��MO���s>�����~���\7:�ޫ]�C&�z�?�K=A��]�	��7�gTY�f���=,A=Iu�M0�
5}�5y9G-?ޫ_�#���W����.5�U��Eh���`N� ����/������u{j\Rn�W;���r�w��.)��X�_!Z֩q{u�/Ej�[o�[�Ϋv}��oק�е���RĂ�H��QY�"%����"�U�	��/6������r���([�6R5�))V�u�'u=�����|����O�jٱ#�h�~̆9��[N�bi�G�˕F�?��L�%�]z��ۯ��3�c�,�J�	�bz[w�T��8���c��~ܤ�'N��kS�kW�U��~r�ș�ϑ�vz�a@�7'Nu?�-��F�iSjC����lծ�NA���9�#d�j������7���8��ϯRQ)�(�f��3�U�;m��>fE;H� �Է�&�n�P<�`ұ]������1P߽foDiV�I���dO��
�\�/RW�}�Q�[Z�lE]a��)J��Fo�Ɛ�&9���R��0��$֨��VB{_�*n3�p|,�����׿�G������8���(M�)�0-�51=ZT*ϡ\���N��A��?�mRX�ӳ������&�q��i�8|�>����򫷊��m�����P��Е�I��Q��P<v�rurɗ/e�D�.א	��4� w
�g�|{2��&z&���"��g��BEDXk���z�����U$~W���-\盞[T�i��[/ēt�x�o���s�c��z��[�����i�_r�VF�'(ߺ�;F$��-\{�����n!sL�9���:�-d,����E�-�B�_�#Ɵ�b�^�9O�:dx��(S����'�Y4m\w,h��+,P���Y:�07yKN�+�]@�� +�W���wp�r��6���]��;�io�)G��!C]e¿ -A Ґ�B듪����9���n�z9]��,�E܊f�ۯ�L�� ��
��9��mB
���ޝ��E�ڳ�Y>o�9�ڨ[������j7�f�g��0�dj�1���<a��s������ �s���"",1�mn`+�K�_�he�4= �Viv���o�¬2f]<�fU��U�O9U~�LuA�@1��Af0�_�Uo�̬�h[�RP�+����[ݻ���ufs�?q)R��q�}�>����xh�X�eV����E��ڴ�
�pἳ���E�#F=Z�����b+G+Wn켨	�IT��Q#*}n��
Z�L�\!c�o���kq�����Wg���"��}�,Y@(��;;\}�~���@&'/xq[^��k�G��=΍a��K�/�v�/Ad�- � oC���:t�o���?�惸�K���]y�
�4��A}Tf��^���&O"�|���?Ìg�_H�>{�}�^����k�fG��V_=5Tj"���`����w ��m_k��E�e�J�K��E�A�Z��|��|�p��SX!��7;c�H�=�Qw/�o�������fa(�ջ�ҵ�{���NX�~�YQV�/��-s��A}mgZ�l�%	XѮ�-�^��歘�X�s��W�"9�3�������|�Śߺ��w��2��#�� L��ލW�2݈{@�i�X�U�������+���)@����C��o��qBD5W|~u��L�HR�Xn��$6zw�g�bJwZ6�n��*���!�Eu3D���ơ�J���v���p�g���K�M�)��<u"YP��b�z�a�t�:�$�����u�a3�L�j�U��+��i�7�������p&R?�n�i,��P����N��*�L8��C���x��s�a�%�'�paNffdԲ�mf�v�때)ڔ��ro��B��\�p����-���D���8�U�������<(9u�K���
���)!�i�:����N���R�W�]�u��#�e�M�K$��*}e)|1~�7ŴP|q[�{�t�qK�C�:51�Le���]�R����k�J�
�ܱa�vz���K�V�D�ߴ:E�A������3�}��@DȊ�!�w�5�UFn�E+���`͆S��^�mhseƊ�	���_Lޚ��J�!�!�)�%:�!�B��U}&?���L�J�NO%uh,ݤL�S���-�xAF#Q�@����� NlS�'���e<�.d{
58#���}��3�Jz�oLv��]��C��C��R!K��Y+sᴵ�;�6n	�M/���h��O������ַ���[D�r1)�K���zs�m���-򛏝�~JRi�3��>Od��$��L��l�'�]�ˊ>OT���E�{]~[H��βM���m?3Z�<���,9�{�EL�)�Ж?�j>؊#eY�1Ą~����! λ&̈́�8_�NԆn㗹:;J���^:���E.	I�I����E&[T�+�z<�rҴ1Z����z�Z���.���$��qDÜ%;	���^�5��-yLwب�T"#��ڝ��GbCJ�B��44�qة��Q��!M3z���,M���{�($L�5����<�3#jD�7��Xso����1z��&�R~A��)3�hG|�\�&m�S%��T�ǻ&pD�S��F��e�1���@���KOs��˭"��t�g�5����i,�����$�Qd3ΧU�2p����B����OY>��y�d�ߝ�?�.���*���X�(0�g49!pF�t[���yj���o� � ��[�@�����Җ�ϓ�],��/%x��S���#suQ��^ji��N+�ؾt���'��J3��IDA�%��ess���[Iaу�X�XN��������[��������W~��z�r��0�1D�Iu� ��ď
��ۛ�Y�~a�
����I���p�p�Jy,��R�ʕ`:����a>[Zf ɔ� 5�i��#����*="������X�0���c�h7�7��A�҂m�2r�5��W��������z�痐#�R����
}�8�_���>Z~��L�$qXx��N��JY\>� �'���Qa�M�C�ฺ@�ya�yF[4��N#���uވ�m��
�F��s�'#��B	����J�R���č��׌�#�Q�Q���/}����Uy��q������Igr��o��e���v��Hr���������?[	���?��V�-�<�hZ�X��E~W!�4/���΍�wV"�ե!)N9"u��f�L��0�~�\�4�`jǱ=�	���6�K�ͯ)���n

���	�?�՞���s7��r����|�����i������>���w�O%��y~ց>�[Ԣ�jMe��§M�]	E� "E����{B�,�?Wa��F���m���"|�n
�b�{#L�ֿA�>������0�����=,w?��k�\1��
�e��(��S;�Wߧ��`+��;�s��{������
������s����^B]�h.6�JS����rϹ<z$���<+���q2����g��}�"���F�?-��%����+�,!�܂��i�B���0��6H(W��j�tQ� nX�h�T%t��{�|�_���n�_&�bo۹�7e_��lڗ}��B_�1[䒵� �<c�QS��B���C�9��s�e��=�̅V���?�dkL3��a%άW�E|�qJ�>7\�[���P�O�iL���_�]&9�n~�������ǔ��*}�����4����RH\ꗖE�yRg;h����u�M] ���7Ct�8��齴P�cx6��wS�����x˵��!�`��?J�;�8�Y��ԷBp����^�&�fJ�\�9=\��jޱN3�����.I�t2o�2{Cl&tt�km��wa-� �Ζ������>?H0q�U�mlE���1�wV����Z��VI��dVJ���2��P'ވ��For6��]��S���@��am8 �����S�&���Mp��p��z�K�� Xv�{8N�(��h7�_�p�+���i^�R�REA�IG4���[�	 ��K�QȞ�Q)"�l��3ݼ�1^�wa,p+!`����[3At1�&�O���o	G�'T�@�5X��Tn1����%_;~j�|��]��W6���jm�(W(,��K�+�{�ׅ������>ͣk��#7����ZOw+×���J6��q�>��/E���/5),�mk���GF��F�c�R���<�q�տ����4e:'/��;��0����kU�d�j��8_'Cq�Sv���G~~��tVUvMR�ah��j�*{L�N��?=)�r�l�e�%ǘ��KќK��6��r��v��p��PJjB	K�X�Bٟ�|�#4s�	U9:�-���k�B�,Fl@�2q��|�/J�y��>�j���-�#���4�x����OxxV�$��P��c����hNh�t�<@W�:s��[T,�ύ��[�rM]��~ �P�I��̘|��l��
l�"����s]b ������ȏ=� ��q9E�y������ѣ%JY��⤝�U%�TȦ�i��崠��_;����B�<��`>kP�R�,ݰ+���N[)B��b����s�~A���#��]t�i4�%�Gx�qwp���4����J����,�L���.!����#�<߾ӱ�>��l����#d|��k��$e���/�Cm��%��@�Y�� r趸��-=�>R��[1hU��ٻY��Y�F~��a�������j���G��#5��>���4���^�G�l�,(*� �{j�C7���$�@�F7��;	��^���?[�wzk��r�՞�w�PTo�م)'y�����~U��Q�
%a���C�GU�4pHh=O5�Z����QhXE��.ZԪ��Q-�T�9�:� Ș&�����΀���A�F��Y��<�,R,�b�e3�6�oE$_��j�3&�;��Q�9�Z��{b�ݚ�ڊP�����_�{�A��:��q���Atr�xN�|Mpi��7�_H%#�mm\��q������|{OÿvI)���{�O����f�zZ�ؖ	�L�����������wl5��D�㭋��,�d��6�^�/���	���a6�R�j��{7� L�_xLX�)��uKO�����F��:�O3/<݌���)�N�up��J~���"T��0X�J�V����?i	��&��x��Y�Ǥ�}i.hW��X��k��<c̔y�J�*�Ӏ����-.�Ѕ�U��ca����KYٛm O<�jU�?j��WL����h��M~�F?� ��\j}r��T����st;L����y9��ָ9���0d����%[7�l���xV��4��Wn?���P�U�l+�A+s"V*�L�qttuv�4��(��\v�NA������ԩ���<�����,^*l�%ò-�;�HK�o��zN�@�:���V��OQ�}\<�q�M�DAjأl�1�J����̣v��S���>Wp�A�4�PŀWE^c��b����l6=r��M�㬛Q�]�8��!�uk%n�d���|�ao��qU����ay��c��Y����u���DP!�p��y_�r���x܃��<_��7OF��o��+�PF�xc��^���07���yrh�0���?gHW��:[�ao��6O��9u?�]$
��D)%���T���Rt}��zk����yO>ς�:�p��͎�Hb�=�\*q��F��5���c�1�r(K%"J�iN�0Q��f��9&����(�IKZ5�>�Z�������o0�SXք��QT>�;o_�W"63@����sJq�y���'�:>M��k���i�He���d��������n��tU�G(tC���O��T^��ϊ��#�
v8�&��-b����7UΑr�
rL�l[�B���3xmQ��=�zi����:��_�,��.�oH���m��,���X /k+��x>p��W�i�9;����@�����ONU��s�^7Vq�7f���ċ|4+��2F��M����������	^&�A�bZn��`�M��1�=�oϡ���ib���̂�h@�=�Ð6p��s+Jc��.�i�y��,3{�C^�Z�2<\�a�+�-�y>�}��
�VۏN�.w��r�\Ģ�5A��4��h�$)E����޼�\��	:�OH
W��l����C:x`ɭ��A)�0���I��RbA��5��-� UV��;�C�Hԑpê~�+)3MaD���]�E����1}�_�P�? )�K����w��Lc\����~1fhN}A���j!������ơ��3ՕQ��78A�I��E��bY%����R�d�j��(�Qh���P�&�51]Dx�o8V����:�ǰnZ����`�-��d�O���W��A��Ƴ���3��Z��Î�U�Kqй���p������|z�Y�F�����y��\�g�x���Y=7_���m*�d������I�l���:Қ)�	����w�û\�أ@�TE�%�E�U�a�]
7�~�ņ8l��5�!@��A�KH'N���cŌ��S��Ε>snM��r�<�Ы�C�V��^��R%;+��̻BTLԾD5Q��Ev�:��Vslޔ���'F�j��������c(�[Ōug�B?A�z�� �b�R�v�Ͳ�v���>Nδ?�HS�̯��?�5����}N��	Ez>��-H�ۢ�x?��8J�/��$����/�qv��bEv�I�����j���-X��RXtѭ�%�9�IDU�H��~��8&�+����3�Y�"��L`��_K:W �N��K���[%ʬ��t9qbeLN�J�;[�e�[e(Ej;͡���+/U��?>�*@�J'����Z�֋U�&�t�Q���V��Xj`���[
Ǿa����ڿ�K+.����^X���cԈf=%:��V��IEΜ#��~G{$(��֮\4Ŧ��
IBN�9�R-u�1���V�LK#��0�'hp���T�\@������Oa������s��L��$!��Zq�J�--s�ܾ�`�F-��ڔ ���fs�4�:�����@)$7&������7�E�����n3��,���7=4M���dKs_�&߱����I�����?#�-�\L-��()��S^J�υN�C֎��H���1=���F�s�Je8���Jښ0$�9b����������v��+�^��4�����omu�x��x��ﶱ�n�GC��x�><���-dXU�ܓ7��'�ˌ���L���v�D�k����5�Q*<K
d����0,�jh���'�\�s|���T�2�c��"ߙ��o5�_�K�!�t�L(RpZ��c��r��slĪ�
��
ƢƵ�զ��]���@k�k������%�$QМ�z&9 ~�[�X��׳�!����H��W�9�(Ϥ+�U#�cl�tk��?Q1��UD75}V`\��~�Q�BU̒(.�3���Ho�!JY�6Yų)k<���ۏ����T��C|rˁ���Q��]�����BR��=��6I�"������S��m�5RۧcW�+.7/��dk8�7���݈��0��ˢd��M��U�̈́M�C
�7�$n��9G��u��l|=O�vӯK� ڵ� k.bͨ�G,�*�Sud�S������tG'w�\�r�DC�������Ui/��:S������v��C|+�\��?�9�hi�͛ޫ��>���OH��_� q�����ָk�M����w
��jԽr`�Ź__����C6y����������c��V<P�RWv#U�� o0raǼO����%��\�|�ZE�HH�	|��%����Iף��c�kq<��n��S���:!�{��`�o�'y�Xْw¼����9 ��[�m������n��b��0~��
�&p޴F�x+L
�(�k%i�<F	��*jݪ8~xq�X�{&��Ƿ�T,�mqR�FH@0��Ƨ��6�uy����I0�z���1k�U��9x�^~�S��$"��V�.{�Ɖ��N��i�mr������S�t^D��C-}VY������+��}T<4�^����x�ޮ��cG���ª�A�Ua�Θ9��1-*
��y7��95��<C�򆀒e�ByK���hC~�/���}y�Ap6�^d��D�Mє�9W6���_���U��B�
�o�c��n�tT��r_�e��!��E&��L{�rf��^{q�>���=��L�1S��G�����18�Z&A��&�	(QHEH#P2��L�F�Q�<��g�P�_���9�{��T@�9�ys^P�. ���qqn�Դ�5��~�~�%��)���C	 -ʿ��jE넹~���FP��fo���y��Ǹӣ濿��:lҍ$�,Ǐ�A��!0w%�OI�r���P��4p����#@Lܷ�M��h�b��q�4�����h.��iAX����c>bi}�a�L���s����c���j-��w�u�lO�`f����{�3p�A��P��z��&c�o�^t�J%��I3$�H�#������纳���>	k���c���]��a�)����k�8+�?[g"?ΗA���9��͉��m_�dT;@d��`(�7;`����v��6/���������I��h���;x��nݱי��֙��&�v=��9)�c�df�d����yD�bK��I���]�!Cn��N��tP��y�}�����˻���y$�g������yΐ���5y�ӂ�O�=vao<�`�׶�@��M۷P@ͭ�9_�0��W|�
��۪��ަ�w�D���o�m?�z^�^Nh^nFH2+P�
�_��b�mPv\�J_�0u�	��SkF��]��u�[���F��G���$�9�<���f���[3�����N���ӎ��7���S|���l ԉ#���W�#4ڂ&�
8l"l�?y\	��-s2��L `/Iu������W#�Pɣ9��?{a���LǓw������8""[�vj���2?����'?�����"J�r?4�Z�����%���g�/9�6�İP�=i��t n�3"�G��H�E��	3��~�@3L b�D�*����^-���c�Ԉ8ZIH�,���H��mg������sT}�������;�w�a��s�qoQ������	�����;1+��Ɔ����YL�p��8Y���;;����ϕ&��N���#^}������u�U��z'�)�q��kֻ
�F3�"[�[��>��D�oE�zp3î�Z�4��0�t�Z|�|�cw���$�*ܢ��7�������x
#$%$�/�U���)���*��'�e��2Q��9
߹��%���aJ�є ULY�"@r��*�w�"µ(ʵ�ʾ�t��#�'?L	��o�TA���;%��υ����_^nE�H�=د�N2�I&p�d3�h�̀�>H:#�R�ac�����tՙZ��ḡY[EiB�%�a�Ez�/����k<�'���Ә����U��ӓ�ݾ���x�T��s�d���mbN9��m��CZ�>p��|a_��l��.������8��`�j�Bb��`��aQ2�
N�F��(��Z�za���פ�֔e5
�zLN�-��b��O����'�F��K&}��4�H�G�ɧ���|���L�c�yխ����+�
�jy�N��%+B���w��Wh�&�~�Wb�AETk	M��`q����u��'CĽ{=��'#lތ1:R<hW��4/��-EM�,C����W��ې���#i��3Y�e�ҕ���Q�$�a�n���X]A�a����Q�� ܅�-�E6p�-6�r�Q���a�ܿ/qS9�A4�n �*S�H\`-�e)�9��?Aq},��|B�R�qR�Ӫ��-)K�_�����F��Ո�	��l�c]Q�U.>�m��7�^y�Tu��F
Y�<{*]�/�P�ӿ�LQw~�ۨ��]{�~�HC�:N��bWk��J��2a���תC�!cy�]"'�Ȣ)�@ݪL� !��h���2|�v��y�J��m$g����\�-��p3�z84 �B�|SG�;�x杈�8�#�M���ϼS����+z����sk����?��NKl��j���J]>M�i�\w��k3�]fE+=#&�>��8Px�M�F$T
q!����:�lhT�ê^��'���8����0�h��&��˒{����	�ʦ0#��y̐Ϸ�"�5��|M����\�Hǻh@)��%�-����a1�J.m����j��x�s/��%��E�����=ZJݏY#C����y���~��izC.�萭��O)�È���׸|�N�(��Uq��e�m���U�פWm3��O�B>\ܯ����-W��X׷z����ۼ��s��6���q�?�QPD�,�S&E���x�Eo(׻	*u��D���hp��a_"I��.����>5�!��������y nK�a�|�iD�iH��T��䎪��#�󚗕W�݄��}��P�hB,��ɋ۬�E�*u��&��s����t���H1u��M5?�Y��v~kV�T�c@�ewn�^*i���J'F���^�=�g�ɞg.&1��g���=3�b2y���E>���p�h�����Z�c�d��ޔZ�DR�R]�/��}���I���L"�fg[u��Y�;[��z�[$��2W���B�k��|:� �L�l;���	�.ePQ�3<}J.X���}#��"����<��IX+��iA�% ��#�.������[��_#P�nQ&��wu����J�2�R"�v�/z#�&�"�W:�M}��r��iA�ϔ��Q;���N��� �j�!�O1�����}�	2z���q�tH�B!T�tS���l<`j�36��t�#҅9�$��?YxU�b�;a�OX�X�-�q�v�k\�l�<O���jJ��\�p�@����U>�+/���[۪�?��w�5��e�'y���ڈ��+�@%�_�M`�y�S�*s��������ê}��Կ��LA�wV5��J/�Lu���~|
��D2���&�CuA���;J4��lQT�,�U������
�,�䉈�B'�T�|��31�rF��犮U����{�#�2z{8񏃘B��>�Cx��G��:("2�R,'��R�����5�t뿞?���_�}�i_5�T,Z�E�x�1���`)�����'�Ѽ�w�'F;��Z��&ޯ�'�E�Y���ߺ6�3�瘞�>���9�?<������?jN��n@�bx/x-�-���Jt�qͼk柮44ѻ,���"ΰs�i#\j�9E�
Qlڡ>y,��}F+1�$�U]i*�^Ơ�b�
�a� ��|U�������߄9�!!}d��0oq�^�h���pV-�8��b ��a�{s�'��NP3a����H�)/��HnY�6��ɮ�O5���y.�y¿u����%%0%F�mE�`���mŅ�g�R`��CF����sJM�`�o���j$�z�a�Qnlhe��0��t������I�1B��n��L���ҎZ�&#uCM��`)N��1�Q�R�(Y�da!�C��e�:�X�K�A�ӪC��jnP�x�gѠ�J�Z�xA$El�}���>3�0u�`���I��i�X�.!�4�!�0R�7HQ	���sοclƗ����Z�$'z�����G�yn�I�ӕ�XHW!�$(�}���Յml���.��U-���3�y�$��,� r��?k��Lf%݉M����G����@%��e��jƁh�R�m`~��c�hJ�k���� qK�l�g���Ÿ�b�v�h0�(u��&���Lp�Yt~6t2�?$����on�f��KW	m��M�]X��X�/�M�-7uuu'��<�~�8Ns�V���c_�ЛPcЍX�0JM�Ib�	S��W�ӛ(է"��������c�{!�@"�uW�������J�R�MN�:HvY��h2P��[��I���Z��Ɩ��i)QK��s	N��\������⋤9\�.�AΘ����de6�뫏}<�|a��i�%'��� q�e5�4����ek�M�DYy��"�� =?1iiiq�1���S�a�!-�%Ӄ����ǜ�C��ngG��b��z����
�O��zIP�(��DQ$A��H�E�%�"	���P���b&�bH�a������9�!q���ZQ�J`��r$�\����>�۷���[�� �vqy�+��"�cF���"ބl{�D^Ҫ�m����Wt�xR]Qg|��O|�r���r�-޷�q�	m�����[������-gp��5����RQ,�,6��ʘ 6��C���eA��v{K�f�?���l+�P�D���X�= �5��B�&7�� "��D⵾�ĂB�>q����S)��Zt���1�B�`����$����Dg����,���NNN�����quu��<x��f�{=�D�c�CW(mx�ԥΘ|�g��t����҅���6��rX��fC�����0��<��, Q��k���w�mϫ��U��R
����򽏹�_6�?�х{�M�{�m`Q�釬���s�q@�ٳglQ��n%!	>v���z��lݔ���1v�ޫW5���]�$��D��h�z���!�H��1%�ݰ)@^���sZQ��b���5c^�j�i@���V6��"�����#���AX<�|��@�%E|n�z��_���mwd����:[���w���z��+�VD�ۥ:��	�j�h%�n$.yE*���l�ӏ?�(�$c�����Ưŀ倏�A�4�����_�[fI�D ep��}�R��_���'������p�<�����_��W/�gi������"��}�*�-
�#�b����/R���}&�JO��c����g������I���:���X�=� �xI�Dk���}��D׷�Pga݊��ׯ�9a��jȋy�OJ�B����Y��.6DX}���u��䔞_^ҫW�آH��lGnm륹2ar��r`�A���#˽���#��=��a#`Q�]\й�a��1Y�W}�>oK��r"�) 1@�����(Q�ES�=|M���1@�D�+�u��4h<����'�Uh���}�W���../8L��u4�ޙɛ�1��]��m�c�%��,ʨG {Y���{����9�.U��l8w���Qpј~�P	g�2m?i�#�=�yԿ^���Ϙ0��)L�wnnk̂(�h��,�)n%�����`����O�j����z�&�,��DQ$A��H��Z��9���    IEND�B`�PK   �`EXv�Y�:�  �  /   images/80b57f79-5f7b-47b9-b633-c76636766127.png$[eX[MӦ��P��݋�;-n�݋��݂[�������	�E�k����\!	�왝�ew�����J�
���(�<����yDF��M@j P�<���_�7JZt�ppq�J�R:�sO�}�tJ��(�cc0�O�1#3?TN�)0Ч�྾y��;�����w����P��ĕ_�l�3)�f����0*�c��r�h�ggy!������?��G`��=�kΣ���T���$����E���=>L?0jc�#K���x��^މ}a�$�F�F.+2cݖ�qY=9�qF��au���,޸?� \��KւwR��x�����Zֿ�e2C��c�O�2����|�Ri���e����VdB,p<��Բ����bM�z:��δ��Tw��[�'��֮ѰaŹa�2|�+:��n�I)��Bt�rF�&�?�y��g�yɊ��b(u0�4ιʂi�	�q���yI�R���,Xȷ��f�.����ӹ�����)2�(�**�I���ȓ(?O��1˺�"k)`���O9ڋ�D�`��܈�N9��R�p�Ť�T�ը�;��ft�51�~�����/�R��GBb��~�f�U�w��Y2�����z����@���Jz��P�Q�*������V�����3�.��+�NI�r�g�P���0�!��2K�Azmg���2Ill�j�{��Bu}M�d�\�l��0 |9�7YS��<>ȕjQ'l'�otD0ѓ������?���5�����\���ՐrZ����6�앦��u�� C)k�ܵ6gJULS�88Ꚛ"�#�b��3�@�e���h*+Y���sȄ����H�Ӕ�͔�wBe��x��B��hQQ���@�#�����[�74�|��)�?!�B��W$
sKˢD2hqq���#l��w �:+͸30K`=0�q����U��0��b��S��?{���W��p&))�'�S(��;�v��-�\�'^Y*�0�D�!OF�u�Y�ƻ4���jHa����
�4i	��s���RJ�(S��_��K7�m�D�S�bD�W�j��z�s���|??_/�=�@�'=����*��gOy�l��׷��A�n߉.B.�KS����V�����f>[�� �?I�<w׊j���G3�Җ	��1N�$��
�_EI���y�
;��w۹"���D6�2d�Az	A�kw�d���s��i���̺&..x��S颡��`-YЎ7�n�8��|jff��)a�������~�w,yu�r�(C���O6�J�%�2f7o�F�����y��Ѳ5�_$XgG%`�v���������(G���biO��/1	9Mw���v+͞Y�mRm�ҭ锾i����¤E��JRE��Ԕf�>mj�e� ���s���H�ֻ[���킗�_��J

���SĦG���=�{����G�FX�zd��'�:�;o�$]��L�tJ3�j�	\, i�ω���q����:��ht\�\=�s	pO�`+�

n�u��a!t����GH�E"z����=JJ&ٔV�v�h
�4�,�_�G�:��!0U�7�i3�!c�h�N/<����w�7���}!�˂+�_��� F~ЍA�����.��Z�ai��E+�J�O���7P0���66�V�@����Oz���Ѫ��l���ഊ�\���#���&ר ���Q|�$��!->�2@��8���x��a��jM.lhN�ĂoB�-eFŏ�L�7
C�w�e��b#W�۷�Mӿ���5���J�C�6��9�T*-e $�����3�yED��S�	���P ��g__{���'k�Y<��'�b��ܜr�P﷏��I�I��4r4Q=RS��k�q�<�h E4q�����=ZJ�yXr�7�hx��j�9������{��iȳ��� ;tJ��.�@%EG����	�m�!a������E������7�R���&�f>��1;��<*L�V�g�/��auk�����4��BR����ӿ�*��):+Y&�����GYl>^\N�bһpB\���5Į�^���SC�J����N��F
�B���(�L�����бƱPeri>U�A���T7#����i�pu�����x3U���j�Y��7,�!�&�o���o��a�����0ض���Oe�Ռ����l�y�qW0�:..�kL�.7�:��1�M+?	a9V.����r�K�������Q�r�2(v�@m0"5�2ݿ�$�W�2u2�t�<3�ׄt�r�B�#�?��"R�DG5�<6_Ha�i�c�*d�фY��fa�u��c}`���� {����!]�>���		1�{�`��L�,�9mǗ��+�x�!�t���aB����m��K�gu�쉏X��ʎ���k0��$d:�hn��!�҃=���"��:z�RY���	�ES
��a���ZÎz>&�g76~X�?b�0m
��|	OK��OK�7 I���p4����ǃna��V���w5�͓s��������乬q�"A�~%��f�]S�+v��m �s�J��W5Z@`{��,�������cE��E*wV1z��X\v�0�7�c6�ä����b���b��h�S����
�I�^��ݹE��@�v�`���d�.��xJG�o��~q2�"�q+�@b�g?X�����]w�!~���#�E}'�dK�8N ��a��r�8)��(D��m�@���O��2��m����f�C�I�[2�g>���Z�ow�F���S+��ͻ�۹�~)���!z��T�\Iү��Wm���L�.a(�Y�a�}L���pNb�{#�)�j�l86k柊�gb%cK�W�	�b�(�յ��'�K���&���+ƭ^ќA�*��.��l����\?Ltm��V���N�*��MV�؜*�V��9��q��$k�.�q��`7`�]c����	����㥒h�������V���N�����-5] ��ܳAyuj��C��,�5��h�����"gSN��M���ږ���˅<��oa�4 6�纍2/�6{��z�����&�(f`'S���6o�Y�� ����w�Ψ+�+%��T���>$��R:�S�9\��Pr����u9\��""���m3�=�N�S���y�����r+���XOĊ�����3-2fr�0,@z��`�n��Z�j�����nq~�Ft���G�־S��6��1�D��}�E6Y� �˒��+����0W}�Mg�z����e�BH��o������c��'�W�Y]�]'Y={�rG���_ʌ�:��O;�e�ѻ�;~��Z�z`P�&}���B�������ƍZM:��7>=)�D� �Z���d��iе.%J��6��R���7�'�� ���'���q;4���9��IW�XY��:�x΁:�\�����c!�7Zє�rC���
D����ka�1}?��)�8C9k�����i'=�O��޾^0�/�0�����w���L�{�ŧ��\!�W� 3�!��CT�#�0�ĕ=c�%��̇g�[>�u��7u�4L�XY;BҒ��xb4��pӍעg�b�|}X���?���d ��N���� 4L~���������{���pE���?��H䍡dڠR�ئu�B�>_��!$�6��O�
�Fnֻ�T���E�¤St�>UagE�S0�j���C~��;�,�*��P�P,~������	�=s+�P���N�^ӡ����{�TP#@�Ņ��D?O���ZIB���Y%�d2b@��`3*I�����*�>9�z9{1{����7c��f��aOw@#��A�.f5x}ݪlY,�|��Ì���w<
�.e���� ��a�9@e��.�@:�-����(�9��%��C�2?�x� �Y$���� ��tX�*�h��f��y���;ie�g>7��F�t�ښ�:#�?�̉�MN�Е`"θ� L|����y�Y�ܬѻ$����-��YK����ş6�_���ܟ��������w#���/2�?�������O��G/Ie�J�r��*�i\�8�'߭� }�%�<��C:\66��� q�5Bp�a.�k~�k�C���;��o��7�p��===�$�sqչ n�+�Ys)Q���]	"����&�L�Q�S�~~� kAzvU7Lo����J��z�v���&E/�_�ۯl��?sH#�����l9/z5%�+�(���U��&Z�L�ú?�ӆ ))R{a
gtΚ��aVʡ^$0�9x���c�*	�0n�e�g��Z���Χ]��1��WsmE�D�#Kvl$I�!z/~G�z&R�Δ�����ȃv��.���4(㇞&_6_���.}mZZBLNZ/�p��'�w�� �3*���nV\-!��E_GFn���Lc��7߇dΖk�g��I����]�i�﫫�Yj���CHά,b3�?Wx
�$��M�rv�^E[��5��,@�&/s��t9���~���~��I��J��(�H1���C��=_�o/�h����U��]1���j��z�vh�z��~� �/�˻���nؚs����H=mED�|�2�����4����n�i񒓿��gL��N�J��En
����[(	� b_W���r�\��������Q�8��;3a��=p�=�rأ��@�}V�XNQ��j*s���`F� k���t�W�I&{ܢq��W	8�ڦ��N�0�D��O�Z�j�w�wݯ�I(�Jg�c��}���yjw4#���\�B�B�}�������h� �_9݀ڡ<�z1f�=�{Q���cF� {�����#��lϳ�q5�!��6��J.T�q��Md�`�D?'=�u0��I�U����6�`B� ����gr��@�bO��a��ց'�f��H�;���;��?
p?���Y���!8��������gQ�Gx�.�X�`��Z�g|j���]ր�x��Đ����^ʽ���#A�P{�Iv�O��j�N���=T"#���Py$P(oR�r��}��N���#�%,��WXJ�����@!����
n��>��&��U���/�ҫ܅�������� �p?�0��;�E�x�*�����!#�W��Iyӡ@TP�}�hA|<�����~�>΍��c%���W�hii�4ܯ�
��X��	Me:M�T�)b�|��ӶD� ��_^�Ԗ�û�����ޙ��2��jK��/���;�	0Ʌ�$��m�x�=y2lj�Zc�j�}z�]�,���`�\G�	`��{z���St��ePeH�^�uJ�c�ԉ�o���y�Q�����ݙV��&� �i�9`KT.��(���<{zzz��/��Q��T>��߀|n�0��_�.
��A������}ЁL������,@�]����TX���kS��@ڤ�xw�i)2ж�{�
�MWb�T�%,
6?�"�D���+%H�m]�$�P�)��'k�����9��)~�Jѫ-���`�N�U���v#@U���O�!wj!�����О��=��ճ)-�����g��PI����×�q�mc���;E	�&%�t�q���MT��F.�����u��p�x]vn�_�/�&a���@�_^^w�����3�v�j�� ���2�w�N�������/������c�gM*.f&�Ot��(B�D^��3�G���6�Ej�J=��QE�S�����'1�f�Ӟp�&�B�ܷދ��%�?0���Œ�tAc!<["y� ������Y�#�c���c����Z�^�~�2Η��/�h��$S��~�8tL�Q�o2�>����e㢬�rf�2I�|cjR�_�8x@���x������\~�����d�X�3Uv7F���Sv�mȿ������5լZɄ��41��2r��"��aA�F�B�O�ED�.G5+R�����ܡ��<�<=�=%��w�=���������{Fɮ
�e����<Uu���o�Q��)��.�Ѳl���v��S��{E��h
�z[P�-a(��$��֚d6�S��_�ʻ��wp��Q�gt����?[[E��ަ:��(���A=�����_�"e��wZ�f`e�-��+�F�&Q�O��*{�5���-�!��Ys���R�w�{Y�����[m.o9��7�C��~9÷h��(=܈Fz%V�	��� dO@F��y1�	�gM8w�8�i�ЁL�P<=���%�I�x�T�����z�p?��h�U��@2�ח6ۺVj����]�o5��JČ����٥f�)�eٝ�?R)ezl��a��a�7�o�پB������m'/^����R�}K�B+NQ�L�]Dqb+D�'if�*e�����簃���HQ6E!ᷴ<<��%6Eډ�PI���UxH�s��h��HSR#�9���� ��I!���[�3��ͥ��s���	K5Z���U��ϼ]����Ӡ^�k�W�`��_.=��*_�	�����[��^"(2ʓ�s�: ��}�ՇR�vklL2���%�դ<�O�b�a��H$�*4�s��} �Dq���w��^f�%q�{����y�=�l�@ul�)}d�nG�"������G�6R���w���t3M�0��ްRM��0+����9���M8�z�l&��p���AX�/�s/�T&�a��G���F�-6��;�SB�����.�7�H9�Bc|P���zC�f�Ҙ��a�K�IG� K�����/�C�_����þ���d�$��б>�� ��u�>�4�/.�����.�G�+r���6�2T�p����E�1��ߒc%D�q��1Ժc?(������b?<A�̩�sԙ�N�~�JnW���ߍw�W�f��P���@�½�d%ԣN�%J+j��##즕�n��-��i���E����#h�,�7��=:j��W�F��i�Wߛ~KK3�A�Y+��ZR+���A-�,����u�����a1�E�(a�r�@Fm! ��a夓���Y}�_o�d֍�Q�>mo1��CE���J X̵3�o�8���(<D�Nʰ�9�[��o�K7Ep�N2/J�ؽ�:6�#_܎��o��ϖ��-�z�Sw�0��$���Yԇ�Tv�3�.l��-��n��G���{�&��k{߽�Np��SdT ��7`@�)��AQ�V�d���?kf�,�"���?�G`c�r�ϰҁ���$���?���%م-�+ji[f��J�X�!>���PUZJ_e�"�]�2�4T���6�3&���Ay����M���\Ƒ������jLQ&���U�~niEa�xl��	��X6vӾL�!4W%�'��r�3�L��6�������7VY���Lpy�a��1I!˵���TXG~45���eGg�s@���/v���;͋��I#���MøMk����z�&�Jq��1=.��8LV[��j���Tn�;,
[9�h�2�;��
�H�y��v�<}L�(���y;	��<'#�0jBby���鼄����m&�ЙJ��B�t��%�j2�#H�V�M.��O�8)���A������ 6��%��$��lQ��C�c�&�.L�����Zɩ��2�X���R������.�S���{��Aư�N��	D�O���I���T�1~,Yx;Yχ�,�D"�2�b1`º���� Rxa���Ah^�
x~ )�Ez6������.,1��Uh<>.��C��]�r������d�S��M!��u�4X3�������9P�>��Ő�[�RY~ԁ݁�O�Gj�.��~2�@J��s���)���5JK,W���~�s��w�� :���v���_�T$�|�x��ԇ1�ɓ6(�w����d��?D�x�\R%�8J"�^"_���?}��%ʩ��M>��m���Z9�f4�
= ����\��5(�/e�^�E�9�I:�Y�6R\�t��P-l-��*�:��|�݃it|�D,�$�&��2��EvF?��A��dUVEFd��:X�������=��B�.�ȓ�;�?���U���'qJJ����=e�t����Y�/������%�_�V<�B�m��S� ����ۜmV��\5��T���$�4�-]��	�ܝ\��KJ�Ҕ�F`��߉�4�E8�6>��$;P|�8���ZTB����S�;���;���h���!��y���Z������h�d'���V����"��)yjQ��W$�a�٦�ʫ�8�S�ۼ "���pEː��h�<�?jk>�f�i����0%ǧ�����rE��sj��9g���� 'guYø�Gl��2i~\�v �ͫ}S�A@���Z����l��}?P)���V����޿�q�Ģ� U&&9��ߧ����׉��`n%��U{�C�6����e����F�3��x�_����ԅҍ�x�T\WM?R�[��@?���t�|�N���T�G.]$]GJEF�ܔ���z�n�.���f�H]ػK[4ހ�V�OW�S���>�C�(�yd ��Ɉ�bB7�\q+jS�٤+8/G�5��9M��:�I�i��G۸����^ ������TG��Ǥ,U���w�͌c�#���q��3��ϰ�*������w��x��(.����e��(�L�`�+�~ę�i\���ά��Yo2�q8�e׃րl�8��v$�/�	���hA�����?LU;�5-|��X�B+7��k�(����c���G�����"/�{���<��eT�Ne|��д�,�������P{��t��oxo�����*8�'�(������&W�)��	�u��k�w
hhK����Է��)�O�>׊L���~/�|�i4����D�\�;��[���|t8z��էF��$�38wF�\�o�d�\�򃮟w��x�z�� .7(+�6��I���sݺWM]�F��Ux�ِ��s�_���Y�p�"��t���7<{�]����o1@�ћ�rյN?rPﻻ90.�ׇk2������r]f\�b �����%�3�"������*F��ٿ��VN	�H����G��U��Z�'�*g?!^�Έ?~�h����'4���=��P�W����Y�Zp�GGG�C6�����4e���[u�u,k^�(ژ ������@��i'��EC�RW�ּ�Y��f�K�����q		���:��_7��d�	�w��_m�K�ԯ�knVt�J�#�u�`��sw�uo	��-�Ȗ�} ���T��Dv�^�{�р$�`9�M��!z����Z:O����gF)��i�����ֱY��OO�wz@�FU�L���ch��l��H�����?{xX	�܂Z��؏1L.�&�(����l�gk��1\V��/.x��=�A�X^����^�i&�r���3R�ױ��B�.��s�[<�_C�a�ڐS��~L��
)^E�f�KHe�켣�6��1W�}�*d=o������~������ǽ]�^�d�NLN�f�F�,���p�X�������k��㖜Uѱ�Ra����/�	��r����f̑� �_~@���'���j/a����̂�+�և��Ζ}WՎI�J��E���AAy�Ӯ�赑:DO�y��vB�Y&����Xb)>���_�vթ���`{0q։?(�pe��+e�.�*۝�q����^(��N�E\���&C�9r���)p(�p��������D��uX�������-
�����/�.Be�G󤳜a<�3YE{�ֺz�P��ˮ)VO���9�r�C�,h��u��b͵��]���ÃB�;;^�#<|�20Si>�%�V�$zgm	N�o��r�Wsp��R�ڨ
���L��>0U���α(-]��1���rۛ�����ԋڱ~����f�ΰ��ɶɏ?�n�0�^^�}*w�!$����s��C�ykm��#�p&��*8֓O5�4��nN����`�ǭ��$������N�r��J��[�E4��Kp�8�[6�\]5����-D��1Q���x�`I;y5 zT������ઐ�#�nӋ~v[�]�]3U9��yh��ߦN��8�D��Q{ŭ�/>m'�^圂/�zn��P����P�o��˦���������\���:tޕh9ۻ�YU������^�R�1Ǣ�$gs�s��*&�"Wȸ�-�ˍ�Rt��hV���rsU��QN?�� �vf;�XȷQe�q��~��<��̩(�q㌈���5Ĺ�ņ-��@Mk���hFK�=`�_�����[8z�������g���� 	������=?���B��U\�V� 9�冐v�F��"dë�����N��F�^%�r.�U�w"A���	��ɿ�4V�� 3Ahjv��l���?�T (([�������WH�1z�]V�E$S�t�V	�T3 -3'>�: �P^!{��r���-���C/,���[	������p'>+!��koD�C~�Q=���f�w��J)aʥ[������s-��,�o*��͟����vQX��/4ɋP�-��,���&[�*W[�c����H�;e��TP`�@�r2� ��F&��`lə7�^j�X�퇭�/�o���"��+��v���ɫ��՗Е^i5 ��N�|��dPVV����z^�G��I&(	d�H�I��
K}a��;-e A>�6�m�������BS�t�OlL�jMnW��,��Nt���٩0�����l>�;٭���Nݠ�����S[m..�o�Տa.9��L���:f&&����i;.1��h�A����=�@)t���zӫ�l�"�/^'��e���|���w=��3���k��߭�2�L��=L�����M�m�y	���C�G�C��z��>.K�i��j3���S�ݏ��M�%�Gi5���3�4��p�\��2��J�\A t;�&�G����X���]۬/xf{]����������66>�^q�M9���F�#� ��xR���=}�c���f�0��f��s���ٵ�.P�\�b��L
w�v��G����t�a���� ������������V
@'����e�(J[�^���_��V�_�r^6V��ӿ��="�¢�w��*�U?�s�fR�d$����}%ED�ܨ�ӳ���,����-�}�n��|��F$���l�W?x��MDҞj�J������}� ��������E`�Q44���y���$a�ʕ&�f�=�~wǢp���MD�e~W��g�x�h����,y��4�z?�蓭�4�N�}[K�rp�cg�)�K@a�V>Z��ɸs��:8���-=<<��,S�6���G�����o�^|��XҚ�s�����ԕ�t�y�E��Z'�O��#5CXbo�6ɅT=�V�k&9��C|r��.z�V����D3�0�(��^�
�>�Ȃ�*��3ss�yrG�\����U�Qy� A_ z���� ݏ���N	�ց���?7Gd�u��u�x"����KbzoFeX#�$�G
xk"	��ʵ8�#�N����y�J��z��< ht�F!����F��v�����^l\����^i�Ci������Dl�{��z}42���?�93U]*K8��XF8�y��sA�k���g*�@0--{ް��H���ys�ؓ`�O&(�PWD#�eݘ��\�t��t���7����_Xo	����R# U�)آ�^e���Ã�~���V,�g�S�pKL�R���{��?ZN>�3Xc=��ל7x��*&��F$,�G@��H���Cɴ�!/πx��!��@O��+'u}s��->'$ �w%?�����d�Lz��,杛r+�����eJ��SrcL�F]��EM��!HhO����sx%��{?�|��h�0��+'��}�m>� o\�2*�n�#�Z�}MbR�|��N�ON�@���N�OFD�*ZHI~z��6c�2�rO��)Z����R����Q�x�����9Ř
��n�G�U9�H����i�~ܷ�"/��Gre|[���eX�z]3r�wz�c.{��h��AЗ		m�֋L)9�m&��C~���Δ�^���z�ʬ�9W�$D �%'�"��d-��Җ�8'U���w�A�F
Q.УY�ܕE?�^�<k���-u��ʦ��f��������ޖj��������c
�@�	9�7�7{�&&n���/O;r�8"�5���uX!�:7���<^FB��ok�<)���g��gA\m )������s�hC�]ܶ�T���B2����b6�m�)_�-gl�R�\��</�Ԏ6�v�6�o>݈��h�/� ����=q}⡝1z�g���mM*���fg� �ѻep�q�Y���"����D�������DёA�o�L�/�~_���bQ��ٙ����@���j%:��Y�"�@���&�T7���^K)�� ��}���xd�[=�`՜K��k��J�F����@��a��g�"=<��!��]����.���CH޿�k�����ݐ���Dg��$`T�	60��"�;�8�jtu���|b
������ƛS��ΰ1����^��蠾Ql����"i���fK^�+��$��4$�e��)�#LT��F�dAZI�q����Z�^A�}��;xG��/���|#�U�?YTbU���Us���^+�����}�m� -�>-&�c*��[�on��3�bP��D��ևVA�'}e��C�*E0}�[�F���d+D���]
�I�8���vYJ��j�.I~�(X�*��Ǽ��X�N��D6�4"�ǣ�܍�0��������ޥ�`K�*�N����f�SƷ�቙h������������H�L��l��V�zz %���RW#?�V��W|��$q-d֎�|��d7dT�;�UJ���#�Q��2%"�s���Ǥ�R���su������,� b�5�>�G�॒�L�*G��I�YG�&���:�y�K�J�ځq��%=�/���<��"�����s1�:>�}8߁a��xR���D�Ƀ]DJ+�]�%��S��NW�t�9(�J�h%oJP�`x+�eo����$��Q�K�;���kxؔ�S��{G�q4�"^M	�g�m	� �&���C#�#�Pi[x+�g1�P���!KIŐH��P4��/�B��P:�H����HK���$��2\.�D�����(tv��<��IHJi�j�c����f+�p�!�9�2�b"��S�5��\$���iv1��ڤ�lo���U�9��j�H���?f�������%Ի-r7N����v;.��TE��D��a��x�`bW��P�a	"*���r���KоŊ��)@����0����#ᚺ��(���5!���x�E�>����הf�3����t�&牟��-Lt��߾l�6#�0�JK�4��I�N �Û�ɍc���M-�74�҆���&T�k>[�������ʾ8�yU!�M�;�!�,�����l	?~��U��l9��k����</�h�dܠV:�0H����8}{�׿�uy\
*�D:E���؄"5m�>��� �i�e��[�n+PZ���;�$jd��I��%I]����M�&.�̕�H�U��3���)�O��p����|���A_���e���^���AW�n� {�my�윎�u�,��G�i��`R�JnU�[(o�����SK�7��X���� ���V�:A_g���x�p4��t����vz�z�����k �/y�!Ђ�O�CJ��Us�To-�r-�~�B7�����j���qfʦͅ���5����%EEǉ�hU�9�=���it�<�UnӬ������NYo���b��ndy�d����k�Q�$�q�r�/�p-?�Vd�q[�0�@�z�"���[Bۭ�e�7�<*#��l�Ԯ���̱@��������"������'�L�f>h������~��r����[���y6��
TN�T����'m�b��gyV.�w�g�n�E���_0"O��긼�����4����a�>-i:���}��s��W�҆H{�öB������=�mk�f�[=��[�޽Y�fT9����a�a�´�+̳��o�Р�|�^�÷O,�R�жy���릠9��" �GC����D�=�'��)M�N`� �^j'���hH��v�s^/�ndxD�	v��M��>-ä�V[D��W>��k��.�ȃ�S悘U����$�.���$N�hf� �BB��QH<���ߝ�pR �������3��n;a�b�OR��R�))��]��S�N�-�^֢���lE ��"K��~�C�#D)є�I��&�ny�%s�Z���\�y�z��V˕��L9�����~�}��������	���`H���{Y�ʀ�n5e�,&'�4G��U���Y}��2�ǜ��O6>���*���):8�0̣#�p��?֭S7�%���K-�`�'�GKr��F�����ڊ���Àk��E�v�1S�k���hF�)b�<^$��lqd�Cg``���<��p�������cN��ߐ�`�SX�[�4�4������	>)�T��2m66����]�̜�=��$��ƅϛ������d0�k�,Tԓ��,�p����N�T�����j�M��s*J��%����׮#rɴ�֑���K7OF3�.��R���j[[GH];��'P�ĵv6��Ԗ�� l�Q�r饀��W/�7{D͋���R�����o1�Dˇ�����۫�����BZL�Ad�&#^[����C�@�;���F�,-ܓU���"Cv�lW,�˙7	���rƥ��jK�w���a�K�{�ї&��ڈh^~�tkS©�.z�*?s��w
��0�V�83Ͷ��,��w�w=赑U�i����k3�y�I�w4s�7�Ho��D�F#�a�)��귓y��(�-���uF�2w�%dNӶ^��m���^^͚mv=��+x���+p�k��\�b��i���8�Z��u�oi�%ޱ����� "O��G�L_���3P�ء5��{ z��A;V��n_	M?wO"�y����%4^`q�G"�Z;Eȇ���������yb�9�|J5{��|��=,#�Dz�=>J�\��/�Ĥ���}�~ax��5B��5�>����d�@{{#�cH����LZO{5;�V�}L\=�yt���ɥ�����K��ܥ��r��c(�B�n�c}���b�����Z�%a@�"6��M~�]�B������7�o_6�')_k�&���-���J=�YO��I�K���o�J����/��.?��ܽ�?&RU	\��PH$/����`��ט-��C��=z�������Va�=�T%��X+�?lnU��� �6�:N��Յ����s��mG�E<�X��a�����rzݐ>|����X��t*_nC(ߋ�qE�����g`¿��N�6Ax�.86N��Ϫ���@0�`��f�Q���Q���Q�o0#e������s���,�S����3����F�wQs?�9�D<�}j�ߝڄ&�Q��j����2��� �+�2����w�~3��;|G�{O� �F��N����e2(A�3/������?���x���r:��qO���`���a�q�q�1�!��O{��*����q�����'g2������(%�:(�˱�#E"��Y�3�9��:1+uJ�z�<�1�^��
�e̱���D,��F��9^:7� �ol*����Ǳ���fH�׶�����!ڕj�H!WwǶ���%Fgm��yV(�9���V�>,w=i�d1�H\�����Yz�v�f�_�<��!��V�ͅ~F�2S���g�-�T�K07��9�^E��s93����}@ ˎfU���n>�7��i:�ޝ�ƣ\�`����@?�:8d+7:X��Aǉ�b�M���՞>�B.FXN�r��I����g(C��Qz����i�)D� ��L�W��-�n�ס ��8�I��iQ�qÒFW��9��hh��9[^��h���A��$�*̵&ѻ̈́"hԚ�Y�|l��g4�G��g�U!�l)xC{lll��$:q���+1�O�g�O%$����E?�t��\#�<(��Ky�U��w�}���),�Ѳ�y��x�	�[�^�k�M6�dd��َ�b����gh�Erx����l6ۑ�Δ&enq�������U)c���"p1�����ȥ��Q��Ut$Şe���G!��bL��Cuq��i�,6���Z�F��Љ����m����1~�������r��9S����;��fn0���Bg�ηFX�k�ժ�k�6�뛊��qM.��iĻ�B���XZO�QS.�&���\h1��ʋ�L���@^����1��5#B���*����Jm�?�pu���D������Ez��,ϧ�?�m8�
N�[�d��'�������_��YB(_��α��P#������"�T�TO[)y�A�%�{)9  Q����,(=��_�]�x
�� �34�VZh������]�ڮ_�f̈́ɺ��}���i,�?o��ԢS3���.�������-�ͬ����S��x@���Xz�JK�V�b�0�2_O+όŎ�&&)T|�9��uEG�O�G.'%C�%*��P�c��� s��O����z藕�� O��GYf:��P%���	�sF��_th�.��|B�F��������#s�2�7�=�+�%߱>�O�~}�l�q}�iO�s�:\��/b�QՊ'�7)(�$č}���|�e\�M�-�)V�8�xp(�B��V\�;w(��^��C��������s����-��<�����3���|I��NO�Z<���|{�%u�i�NK�Y�2��g�>��!Be�d+K~���f����j7ژp�ޡ=F&&&��4�E��O���#�.Gk��Ӊ�/����}S��U�I[E T�'�%�@2)X�|o�#8P7 �������o�[d�/<Z�TOZ�r@WV9�y���] �r�>�V�N�{V�u� �T:ìp�;:|���Ρ�p���Ӎ�s3�F�T3��l��]�P|+�~f��n��h�Ͳ]h����2:��4˷o�O3�����k=ڙ���06:��������fn�:\N5[��+�,�F��V���fT��RBhd} ������y'�=����E�A b��y���+~/���ҿ�=�ҏ�3��-�*�>�nt��X�#�*Nϰ���O��X�����n�$��D�˶�o�<�d&�%ӈ���~GKeR�~�@���*CpxA]�a�Q�����"��ا���^y:-����m�����[�_��cY%3�W�R����i'��s\$�*t=2�}����˝n�ޟ	��PO)�2iT�t��� �RJ����3$4��L��>���[�/#�e��y�Y�v��/1��
ڷ~���7H�uĄ���a�b��������*dB�EKb��뵓��u׆�*�NN(?4>��<iXT��J��Ify-�������|B<9ղ.컙YH�mz���E�s�ۅ�G-�Ӗ�[!n�t���}�L�����8?Ϭ����Pc9Y?�|�J���d��i��);B�(}'*ӡ`4��p��.w����G�R=vv� H�:ʚ��������Ob��&�e�00'���L���圾��g�5�!�F�r�b-B]=���],�|��ò�+�s�-Ǚj�.l�" k���Җ��}iF#����u��� �Q�Ȩ�P�ʓ�v)��1f�՘"�����V&��t(�d�jR��R΄�m0�<�mc�|<>к^�|��~V��Ij��4[B�Q��۶'�1<R���T�Z����z֧p)����W�2�k�ّ̌�EԮ;�2�^pN٥�ǜ���q�;��p����%�����M���-�$U���\ن ܖJw�O��d�b�F�b���b=*l��~�W��mdZ| ����k�D��ɪ�����$X@�K��ڬ�L%Qzs�w
����n�s�|��-����r�Ğ�@'����_3V�j�;��'E`���4�-�1���^DhP�]���q���
�Bvs, ��В�鮸<Y ȟ>���7��w�F��§MZ#�vw"�3���r�����1���i������zs�:K�3V���p����$m���{���DֿPk>����&z�
�&/�	V赌�طvNMQٷ]�eǰ�qw�Q<`��UJ�w�0�~N�	��ͫ�ە����-h� w���#��G�S�(΅����|�%֍�u����䘽�b�3K��eԤs�m��\Չ��9/���ΫЩ��k���Y�ɟ�rE�Í��[�|/a�p�{ �=�כ�n1�~O��|!qO��~e������F62����	mAR����ud4�%w�'g �%�+r���O݄�s/�ׂ�*\������=���V8HP*����W�U��C��F����&)�W�7X�tϧ"���Ƨ,��4�߅��(;����9��I�XdZi��z���ZG�6��z�]���9N� q�����|߈�S>F����q?E�|�,�LF6��i��e3s��]�`hEI]S�֛�X�W���V�<��k���d�냆����:��y�ߥF'Q��dN�F��,����#dּA�W���V�h�Mc�R%��]g�0X�_��]u>���C�\�t�%��jUL�tTh#Yg���L�Y��v
�,Q�ܾ�==S������X���%��֒tj�l
��������Y�����j��x��)�&A�A]�E�%�F�K)�i] 3Ğj۝��_�����鵽Ȋ��G���5��5�ʭ���N�a!�Pg*-�P�l1+Us�X��9��d������:��7��[�%���%����
Pͼ���gD�����gK�i#���Jy6'�[�Ԕ�A�4{"���5�K�#���#�.����{����_�|��9k����/��v��"�9O,�����zi+�KH�~�?`�U�Y��<MΧo.3F���P����@���(� t��m��P#�&��(��F���D�$!�m�\{���=w<�K��E�bO�jj0�,�g2��n���^jr����x�����x~-�MО�Բ7�~'`�5L�*�:Q����o�t����˨B5�N�R9<]v&�����|lTA�(�'%%-����I�����&�U���$�I��ו���˒��7��,,U�I��c�+��4�( ��r�HK�vH��ޏ��]���!��_��I8��ɪ�6�UtG�,�|��Lh�����+�Ds��l��o�cY2@T�b\~�c٢;\����N��Z"o�B\<�.FR"������I�o4z3��됡Z2�_eǳ��3~�=���'�&<���k�a������r�`zFF�幓���Zz�7�I0���k}�]Z}�5ڱ,�az��wje.*<��79*Z�ε�MS��7d�i]��S��^���h��Sc|��.���v���X�N�:���x��a��3�Cek1�L��=��Q���c���ֺ�>�D�LU8�fB�������8컣cB��n���Ԥē�
�F]�H2�R/+��#�^k�s��\�������D#�\�z���A�h��Zv�Zz��f$ƿl�:�Ěʄİ�QN��d���l��g�N3!���[��IJ��!L��C�y�Pr��S�P�u!��gg���xjL�S�S���/�����ĝ����#_0�Zq�m@c?�V���ӊ���a��̢�k��b��ܬX��h*3�"��n8����� ���<R�����n�u�ȹ 3+۹���ۛ��\�-�/�Ui��K�QCt�_Ӗ��?���t�=d�����3AIGG�.�g�|u�K;���N�J�O�PD4��v��Y�e������y��*.v��Jmt߅G�U&E����V ��m��oˬ�<!��\�w=�/YĄ�k�7���8�	���b)n�)V׃��ڇ�n��E	�^ ���[�!Ws7�O�Oo�/򰜞<���W��S}�TjV;3��c�W@C����M9� ׮��c��Ů��X·r~q�%���zӁ��M�2C�&m^��ǳ��bP�Ғz�L۹5��7_X�����ɀ=aAF�|3H�ϽO)6O��A�D��>ڤ�Q���ٗ�U��U�����q�`;�ע����1%_s�,j\(�q��F�q�E�d6�l�4k|5�3t�m�r���D�%�E�Z_�.f�)�cA|<#���B��O���\�W�K���/�ғlإ���1�ZQj�v��WH(�G���&}��Ԯ�����2����������T>����[�>O���9��w���sn!rL����$��\�Ȏà�Y��i���umLⒷ��`n>���z�}\R�lCN ̫���d��a6õDod�����A_a�Hח�����`�c���t��Z2z�H�~��K3��e��6���;��1�j��^�wz�z��y�o�u�kS6�E����R���������ˤ}זY
��-��6�rV�~�%�|G2j��^�!��]R8�8,i��֫R���=+�C�!Ð�g�}i�x>-�8���+)T@��=d�紼5黔���G�;]H�Z��u6���X�����fǀD���ó�+�`t�$)ŷ�x��`|�#VԔj��I��Ң4�џ���>����䡎V�$u;�-[�dd��Q�r������V��I��}g-��lО�B��5����J�P^/#�q�F��Ds_�>}պ Ш��\�B���tk�'�.�ǅC�
�OR�T�����T��$p��Qͳ�����}���)e�g�H/W�-*����`z9�x9 ��J�-kʇ�E���7H�O3Öm�W�~�6~ݥ#`�3��u��D8��jE�{��^�.��4U.[�$
R��.bދKN����'BsCCq~V����t~�L�XFPŹ[���\O�3h4.a����󫝼����P��!Qc�E��}��(|^Eӕ�{l%k��K�(�	[��0�{�܀����
Fs���� U���|s�%�e�7'�g���韓u䡜E��\]E#eLh�T"��O:���	gy����8�u�ׇ5�E�i�jn�P	��]����TUN�GS_�&�0
1��y�k��d�-���gP�M��>��B`I7BԀ�'=J+֜�.��ss�������4}7�����0*�/�C$�"nQ��K,fP�?��i���Yj�Dx���Ը������ ::����/����������)��H�-��U��u-U��������2���k���v�M�З$ù>(�O��'�ߊ-��pBQ �Z�Ҩh]\D�*.��#T�6y��x��^ѡ��x}؃�~����$]ts|�Yl^|{i�.ԒlS?��̜/C�b66r�� gg�HG��K/d}��@ܯ#2����`��G`{�����I��K୮&��kå74R
|l�N����̦o�`O����M�'p{�x��V���<���-��H5�C�CM�����v"T�����D��4W�L����^K[;�f�O��)W�^���)�/�>�׆�?[�Ў~*T����ߌ:��~��<�VjÛ'�R]����e�B'�J҇�5��Ö|�A 5�n�j��}���<���d�M�|�i*Z�D���({��s*��哓���������ܛ��U����-���އ�~w5�x�2��Po�9N��<З��/�=��Z�K��"y�d�C0�0{�-��w�0��q �`D/�j���=�����6f�T+����;[�@��OD�MY�wרE�v�Ų���^3�c�q3�|Ռ�ÿ��l�~h*��aXO�"��wT�G�MNۍ�t�ڋݙ�%�݅��#ccSiY&���:�<p��&��g�\�G�w7^�Uת�Ḭ6��i� ����C|� ?!�n�z�w�ݘ@���Hbtx�5�(����k,���y=�Y�{V����6��)�ݡ�d�\�av��W�y�xZV�����C'���X�'���f�mb�S�V����r���6��#V#E@-u�n��F%.-�T,�ݾ��zl�Z���Qx��0!���#��7șxP������YdBX{������2�~��ѻ����,z��:��V3/�+I�=wi1G����>�B.I!����Z�E"��g��\�VS�.�[��D[v��^t�)�}b�����a��U2Z(�8j�:H�G�ǹ@m����A��$�OpTb3k�>_���9I��i��9�m����S��ߪ��d}6��:����rC@�J��
.u0E� ��j�9dhh��y����H�%��q�	�o��/�y���}ξ��U&�
j�Z�;��~�������A�&�D��v�'},2���&^��Y�X�{��n�	�v�����dE���e�`����z�]5<�ᾼy�{���u�_��_[oߵ�'�q#�Ô��F/*T@V`^�M�D<�����֫=k��y�,!���t�h��A�s
���z�������#<Sin�2M�۾�o���;II̬,���z0�ou+9y�I����{V%�O��-3ff���A��`^�;�Ǔ��+�O�U�52�L�	�C|��Hy����a�����M�'|���s
��*�Ӄ�QY���Ս1|�&�!tD�1�;#������f�j�?�;A:��̬g�@���mm�ˁ[�z���� �����ra�0���A��kzV�j�X���YF��7V��R�6x�-������UH��������3vׄwzz����H���cݶ��EF��K�X����#�O)��#$Sw�Zf�A8�y��}��������y{�v-�`�k+~@�C�F��n�����3��M�óD�bx}�y*`�p���[z��x�9Y�8����o>ky����yTp0��=����.���'W�s������"��NGR&;IGU� 7x���oS}�3y�?�ȶe|��s6�	K� ��-���l9�a�g|
E��u+�n�y�{u��;�lڍ_^�6�����1������4�%��d�WԜax��
=�
&�[Y-��sG��z��>�C�~���ǅ�ǽ�,��א�뉹vO]7�Y�	
)��͒���D��RA�}�CFff��������z!��z�ǜ��Ǐ+�T�9~OH��3��0�w`UL�>��pm�v��=E�#��i�A/��i\H*�\N����;��O��g��J���1�c1��;U�i8v��_����6��"س8-y|��TN�i�1� G�c�Ssu�^Wn��	�]`�}��m�����@,�/e3��>�}��DJ�!z�%��Y�vF�ئ:�,��*N�c�����Ҳ�%�z����1��[��mO'�3#njI�A�櫍<{�<ӧC|�+}��ZO�"/����-u��w��i�@��	�s�QY8�,����.�ƈ��@C�2��3����c�I{PS��1��ܯ�3�nOdts��鄬�GF0Ĥ�Y��q���X��S��yl�X=�4Q_J��'���Q�V��c�Kێ��1|��8���
ԛ[�܋���ۙ�Y�#�I@`8�������t����G�C[�K����\IL���g0M���(��1%�q��L�Y��2�WX��9F�κ\�ʎ����}'2�6>t�l����M
&H��9�� �-�$k��x,���>�!Ck��'����A�l�����Y������]y|$
�`R�ӱ�n	ԣ�P��n��]=q�}�p�}5�#������1|c��X�2��u���,��r_^=r��E���?S50X-�屌((zwjM䰎�Z�ߧu����RDUL��i_�3vA�om�B��h�c�MNʳ��x:2����!�xe-���xuu�e��Z�W�l�� �JD~����62�_�����ӂ�-��s=��8Tb���9��[�֦ʪ;��Fuf>�ټ1�N�0�	���n�ۏ��c�?�a}���Q����˵_�$9�*���5ZzRدb6�f�Wo/���o��G]��w{�nq�'��������������R�l8��4��t��*x�T~L	h�~W_y�w!%x��Pz|�?��>Uel,����`eJ�<tX1�uIlw��<��D��^ZZ�;��_�~��#�)�J%s�].je�'�k��V�� *�9|�?�z���,���e��+u��O�yI��$tcNK�6�DҪV\"$&f]�SțK)S/S�����
^p�l� ����	��	3_ʌ��){Iy�Y�w����w;�SΨ�9���ǿl����� ��R�I��N�
������Ѷ����%�Y?7��4�)�ׁ�����Z�z5 �.��,�TL͉J������� \�2]���d���v��M��{1gq	��S�i$�F�a�sb�|�7|�0fϹ��I*|��a���6n;�����OIѥ�Ph���^>ޅ-Kk�~%ˣ='
e��V�����e����J�2&��_�X�����=�O ��Pe�E����g�qi���n r���;�=�<$C���#�>龰�l%��,u��m�>�)'"�,�nJz�7"��n��W��ߧ����d�4�I"]F�@�	a�la��tL����T)t��iR�N�{+��$v�M�&��uf��1��q+8x>jf�ٕ���"�n�B6	���3A����3�Crk��p��-@�Z5����ư�M�]L2�������!����$E߳ć"�Y�������Z�}�2t���v���%r9н��
�q��.��ޞi�Y�b )���b'�P!�(J�&a�R69�b��M4�����3G���O��;�LTL���s�4����`(�n$�)($�-ĝW��y�Z��u*�9��k�<�1Q݁k�;�(/`k+X4h�yo���fmu�O�e8t��XUz�0�H�Mֿ%2j��ZC���Ԑ�R/�+�Xwʽ'�]�ºx���5�6�맿��䫇�� >N�C7ӓt���4�Jja��}�[�?e�bG�����D�~I�Aľ h��#��ºZ�c��2�i"���v,"�kfT�S8?ϭ����V�s��k����0��,�����[��P��2���{^�k\�����QH��@¹C��cp��ʐ��?Cᄖ��S��t��5�?��.5�]G�C&Ct�-�Mj��	�Ň}���E�l�c(�M�������{_��nuS�a'[u����=O%
��l)�|ݦ�ô#��+�����@��_��n1 ��V�4L������G��+oك@�nܒ[�F7�*>��=�>��>/m�����e4:y_{�2����<����}{�:?��̀�1B�����j�к�,۔b��{CT��zZCD �̆ҷm�z��Z}�"�Yy���(���G���a�,��D�Y�׋8��\�8�H�ũ>��Ws햋����z�K;V�׍�؞�T}18�J���[E��q�X��O2�}���u��Ĳo� C5��s�H; %ҵ�7�<G�W��H�Ж^ԲL�v(�@ L'�:՜�E|@oMa9���&�Q.[�����f_Z-������h��@��c�_�v�P�l�M��Z	�̧��/3؅6 ���/S��<T�AN{'^Bf�(�(�V��)���BI}��kE���2��"����c�X����Dy�{��8��2 �s}��T��R��e+�"J	+��c����n�����	��*YU#����Z�����ɕp�w�6.C�1��I^�Oc|*.!m�ٵ}d{R��뙱���%����ߦT��Âȹ��>�(�A!�V�iyA�4�(�����_���] �,p�(<��q���kA[���<��<�s�y`�h��	�e뀭���b��M8^�6KP�`:Ҽ�Ň�bq8T)���F�{���Y���z	\����"��)5����)��û�e�t_/4����^�{J��`�Ck<;���Tq�	囈B����-��<x�EN>Zﳨ�i���Z�_�1�{x �b� (2+��ϻ���-���g�`C�o�����z)�цǃ�%�|ݺ1� �޴v���W��o���^U e�f��^���i���M&�G���̪ѕ���;��R5k�J�E�	h@����%�/���Qtr�È�\ 0O08�r��IG�ۋ4�� \V�c�F�a7������������-w��������U9(]|����C�q�yo�P�6�zoW}/�����^S�hCu���׉7N��0%PPr��Z+w|Mg2٭�ǽ	��|EU8s���Y�1�\�T)~�փ� p�p��uۍ>NC��>�V�`��eXs�09���Y���)��EuۮFuL� Lហ���ᔦ��:jP}Ӵ�l�w�!�5 G�[��/�����S��;������X�z���sV�x����P���Ժ6�l({��8=�Vt�x�<���%s�z���J<���L��yۆ
}�ߠ�F���t�bIxS�dC
y#�{���ߌm�}Z��M�8�'�uy*���n�g��#T��!�H/�w���YVLRf��v]9z��!�J�����I!���ĳ�,�"!~5B7��7��o�$4��0�;�B����T�}��ړbs4t�=℞�#c�M��Q"֦��c�an:�'k(E2fxD���X~��,}|���?�$���%�&�j�n�8�+\��`�d�#�ĠJ��A�x!tH�B<wB����;gyR]��������|kW��W���8+X�>���S��\��
7��]��S��YV9<�ƛ�>Y���|�r��e��%Բ������>�CBk�.=��L��ڍؕ���`m1��r3����]z<�$��L�m��RQ  ��J�ݶ�fj�mK�3嫊�r{�땺�桁 ^�Vh<͍�҅t7��r��*d���9�0�PmK�2x_|�_�_�{y�ADқ��/1�w\��%�RaR�ǿ��� ��_�0���1�(�XWc���9��KZ}��Iv۵�Kݵ���Ί���㋶���?�f��k���u��'f��	f�5�h��sM�hfM���i17_�nz^�~�y^Tx)s�p�)>xFF��Av?(¾R�{g�x[�%����P�O���2��#������n!�Ƶw(��ٸ;��d?�o1�9�~�_�\$*���;���<_�TEϿ H{�Ԫi+��U�щ�G�j�C,r�z��h�vmv�]��E�_�ǻ�������r�x_"��́�+�jZ�ښ�ݼPp�(S���h�9��֦Z�U�V�q�Q!	�KĜ�7�C�r���=3�5FN���3�r�� c��0K�?��uB� �hk��O2�5�Kl�Y�^8̎���8q��jT%Ϟ�]�^xl)�{�|��f�	\iʕ_��o�h҃sٹ�����2o,��-k��1��ӛ:v�ih̕��?=����5��j>��fg��1�=*�g�V�v׉�L�'�y�aH��J��?G'�o��C;�mrL"\�h���;Q/��=s�B׹�c���2�D+���K�쏴b�]@s'�Vd���'[�\B1�� 0��]♰�}�{� �{bh�6�vגд7���iQo�2:�T�Ҏ�Ю8w`�|��]��=xe�(E_�6�~�t�0�Z�I���^����]?�r]��ǭ�_/����|�nno�����J��x�M�ZՐ����[����I�7z@�E{"�ď�GB������#5.Gq%C3?lD��=�`�y������U}E_Ҽ��b����,Tz�C��'�!�����u���4 }σf�>�C�fYp�3b0CXQ�'�f���x��� 
��/��\6��x訶%D�CKvӸr�!@S�m�>\����T��nu�Bsv�,3��e�~�������p��gD��'x�S I7�����5f��ի5��:t7�1v�g�n�0ųD.�;�����Pk����&v�O�����\9;�4�d�r��mc��»��l�ݧA�i�l��Ѽ��
��K����c,Z���G6�݁��畜k;^4��#&��&7�(�cMx���h�w�iS�M3~ăN�s������#P��b[	�{���{��bgE#lC�M�Ϟ��L��8���P��L��m}Tj$ [�G/3���Pi�v�IIa�q��\�+t4����ZS�CS|^`�?X̏�� 7$��=G���M_���5 ���M�t�J�`#D��9#c8�g�7T�3��y����WQ�������V��ݟ=�ɵ��+��+��jh����q�oy<����!7X=ªt��
:	��U�ND�V/+�n>sع*�9�E
�4����^{-�k�*��G�Tf�8����!�4l4��s��yFo[�R�򜃙Z��s2�(k�B͈��Q�(kd�b`5&��.�Γ��Eb)�CI*8�(5�mo�����^.�  
�9^=��1zwm�<�U�O�o�8�G�����f�C����
�@����Ν#�����>�rlf]��R#@m)��/�)#$�b�6��U\N�ve�"I��p�q�b���6�Z��q8�K��H�D���r�*8e"�g��:�[�����l(�s�j�y���M6�&1��$����l^z��b�s�fQFS���ڼ8j>�Ϥp��Lډ����y?X�h�Iρ_�ʹ4��*2FG{�9���_��?��]��^�8��w�$H���n)-
�-7o"fu��nu��>���"��t�P��H"h_���6TN���*x<��_5c$� ��z
�Zن਼���4e�U�z�|}|��}h��;���Q/`�.��p6�YL(6�MUG
F�,w_F�j0�I8&��)9@d�>\��Q���d'��������v:��kz�j�w�#q������6����~w����Dډ��}}_Y(������l^NS���W�c��ȃ�${�|%�:3��,�umq�'?�F@��5��ឤ��h+�|t�����|1n7ge-�����Y��u�4!$�-x�t�q�x�xf�zZo/��*y�C�d��S�;����UUV�\�������^+,���Ή�םc�M��&qX�nѥ3��"�X�q]u\��y��@��U�&��1�e���cHkEj�����Hf�*u	���v�DkPA��������n�!/�����Au��]�3,��Iu>�]ۦ:�(O����:ܰ74��k��W9�8�2����a/�;$���/Hl�iR� 2K�Ma~/��*��[y�ml�3צ56�ד"��*��*��A��n���g	�8mJ�ּ�a�{�i�{U�+4l*��J
������A�~��mnmJ����Ѐ5��>`Z�?K�uܳ�%��I�e�Hb]������q��=L�ˣڹ��q^��H�
�H1Gj:P���"^��.W<�qW<>��Qw���v�xďNi��i��`\ܣ�";R�|ޠx�8���Kk,�i�g��N��R��j֮8���3q{�	�F�|syY�����͢>�%,��2ϙ���>S�4�p�F��2S\j�6�j=y��rW�p���Eu��	Y�P�I��S)�X~���U�#��IGq�?��Gq����D��&�3����,/y�f�K�,��xz[ǁ� ��̬�2a��7�\p�r;!�0I��}�oΑD�ϖFQ�|C>c���>�G�^�$!U�U0��!�n��5ȷ���m���aJn��L�����s���ۯ�IB����oǗ��CYt��~��g�}������w���!8�y�`خ)��4)���8�;�g�K�"<+�{5�!�S�[��*�z`+��Ն��<J�z��0`q�;kjxJr\�M<���d���9�	q4��D.�i�PwC�
����O�?���U�8�����7]�?:rng�R����3����!ngZ)�Ŗ�G=�<�x�Q��3�?I(sqI��������ž��;/�,�1�Je��;�!r�`͑�����|�Е.���W�N�u6�}�b���3����Ko��K��e�e�9BX�˰[�s� ��]hoB��֛�d&��w\[h�/��z�f��iiiD����j|�J1��6R����V�h}m����wW�ѓ�IQ���z�G�K {-kg#.6I���ǝؔ����f�6^���`prrr�D�������_�Z���eLLLp��a>G�{��r�3��1[���pʆ�q%�4��RD��1[!�7Ʋ^�Dk�-`zz���G�ߕ���w��Tt��F����f�l˰�,���ĵf��muv���,����̻LE���4mP_O��{�_����*�o�Tzzm�*��A�t5�C��4��l;���"��dBZX'p4�!�p��.�ك^�iu��)bI��f��z�� {��zHbmm]��PUU}E�D�8O�aZ#Ƥ�ϝ3,�S�t�����ל�fk p�~�Zn?����w6�&++���v�JS�rd�9z0�,S���P��!3̺p�����ڻ䏖G%�F~�Iif֗���h���X�욟D��(�w���5�[����СKNz:�K���!4mk:::^�����[�K)�P�3��%t���h�9�y��v�Ʈ��n$�t����߶���wc�@+P�߿�p����,��a��������1���4�As9�N�;�#��
f��J��-t�
�'<z�*~�a^k'0����p��(f��bd|<є>���MUC�?�&��.����'�`�0�3��e;,�<b	B�!Zq�(M �r��Dm����&��>���L�σ��|.w�NNo[u�+�|�~��7z����$� ����^���&9o�$���~)m+  �_ϳ�]�>��]���s�{ Q�ɻQ�k�0呓C��Ğ5��>��wR��������ko��i������Yl}�\��:=�œ�E' юm	��%�������Վb�;C ?H<�PU�:�]�J͌Ww�v�/�D<l1�#e�O*�,o��2�[˱�F���� ��ʶ��A2��sz��:ڡ���D���e:���9��u�K�l^`y������mqR��oN����>[�RX�:x�ai� ���EX\���Ŧ�ЇF��/�����Ssu�
��䂡;�B���ѱ2��w����;���\�d���M�l���w̓���5����[ �*�\�R9���P�J�4���k���4��jeߎ��z6�#b%�v�{�޼�8
WQQ�HЉ%���c)U*SK��V�Q���s�&�`��,2Z���6��-�"��4��w����s�2I�P�rl��"@|��u�kOXl��U����e"�"�4�4[�Ъ7@enA������e�jK�ϡY{�9�Vs�$��:���Ka���`V�b�|�N8�R���������+e�g{e�򋇔������a���Y}��)#�7) g�&v���	[E��X�hb���0^z�bb
�g�|�\E$��D���|2�� �񃿠<b��W[@$�| UU�]����M�oK�c�(*��/�Hz4l�w�ߔ����$���/��m_�#���JS�3����ܲ�l7�a��j;���1z��[ ��/��3��6��z���
�"��&A�$i�, 1^�F�R9�A䞠�l�%�k��'�=���4��h��3F:��āH7��L�ᙥ�Ȩ�M���miteT�=!߁���!�4QE�u�"�5�ǵ�;�ڇE` �E&)o���m>��x�����/�{y���@��M=6��'��8��R�|]�v�%֓E�b�u��&����!�(iT�B�0a�O�γ��@MⓝV�l#1jhV�NA�I�Dknue�>O@r��H!�8��:�I ���W&)��'��8¯}.9�1��ӧ��:��#���D^�
�K��0�c�����L�bcO����˴c���Fu��X��)��s�ݯ(]����<#������ob�x�C˓���>߭+p�F:�iC�-aZV��S��c|�{PS�e2�EA'QM�hK�a�Q��o�c�ao׹��Wj���i ���Tɯ�)�$Ȋ>*Pa��O#�|��&��U��#��ү4J����(�sB^�NWx����6/,�%{�z�IE:���@ �����{V��%t�Ct���\k��������~Y3���}����@G+�4�Q��X�#4� &h�:}/J�&J�� �����B�@B�cv�S4�lӿn�.�57��$���m�%��4�׫2m��ڹ��4@��g�$�M.T�����n�"�d�+��X����=�ly�N�Q���h~�PUX�~M�'�� e1�4G������K$����EoL��mD�I-�M�8 U%�ZB�tl�#�GƔ��;�ev�\s��S��O�]h�^o�h��W�+���t����&c�-��W�_�¤)#��,s&GUXү��[��IP��X�9<0�$K���9�Q���]c�^�s��+�u��^�RN˄���c�s^�v�Ǫ����JM�z�!�Q�+��������wt�]	S�_1O�x����!)���B*٭��4�k�|�3�`���_�n��C2Ǽ�Vi��մ�~4^��U�ȘrT~�,G߼0jF1�B�B��;xPQ�/��ex0�=E|e<�Q����:�)�c��]��!���������&/�:����A�m#;���{:�6ie�G��qA�.�X�'����XP�\��D�+f���D7��g�-3�Z1w���a��-��Q�So;l*�l�"g�8��^JV	hh�/JzO���Ͽl�"! ��˿��Nk7���<�w=����V�bV�VBs8���K޵Z��/D�X�%	�	�}��C��T�Q%z1��vK���'B-|qV��p�}J[S�]~!� \	�.���k��j�8x��'y@d��j�x�K�8��A����'���01U��a[������HHf�܍�B�w|r��c�vK���#��)��~L�Fc!��dDA�o�E�XD3��?�i�������,n��m�e���j駂���__7�NL��"��rh���
�D�[75Dʜqj� j7�^
���ǃ!1�$G4}�'�F;x�n���Չ�e�C�XU"�R�a�[�3�{�c�r)#�bf��)��N�o���ұ��k'c����ӛ��~(H�B���dө��-���ǌ�KgC?]��}D�@p&��(T�.Tv4��4���G�}F��_}]y4��WK�R��z�6"!�ƾ�A$H[7��r�5B-E�����*3y�(���-S�Z�[D0jtڪ�<�t�������{�=���~����|�9�s��5x���|��f��&kwT/e$�0��Kԗ�qr�p�VR�5��ϐO�,=�S�o�V�5#)���T���f�.�A���'�5-#�q��B�b�p�Ɇ3}��c&ͥ���A��̓�Q�1�6Q��z�&�u�g��) ��}o�=�L��
Z�.E��a�����\ǣy�>�� Ǔ�meB+禇l�~����;���j���o���q]I?\5��io����Ƈ#�۟���d�=��H=g�G������h��r�%	�|+��g�Vp�*�����xKW�F���(2XC�}��uX�v�V|���vfH����2��&=z�Q�n��{��   �Bwa	c+ǌx�2$�PYMs^��T}�Z��Sq�Cwp����Ac�e����!����/����|z�$�FO*��Hz��v-�?�&�0�n�~��*ȧ���:�V�w+c�$�\���ᅬ���Aj�DH1�L�"�T'Wo>?`���_�Bn���2��>1���{�n_���DZ�zXU
M.�y���,�N��Vv�y@8>�7�j�d�E�M;�_���r��Y��
RA�j���Dw���v�TО�[=���&b�_�=,1��+Z�K�_��v��n�t4��G.�UY�Y�n!ihl�q�.@�K��5ɰ�Ξ�&vk���CU���j���Vn�9r�5��o�H�ɚ����@�᧿s��;�_I�rM��g�$	�(�5Ҭ-�q)��:�6�T N�B�:)\�%�
�z�-�}��_%�&?G����0���5hT��ܜr�O |%^1݊�pY/��ܓ����F�B>���6f�R��x�*�x���i@o����5)��Y��;�B�\Z�2p��� C�2��b�i="���:
,%d>�7�!�)�N�V�U��&��k
{]�Y__ ��q�is��)�����,J9��u�}�P��>���p�\(�� �q��o"��v��3`2��J��% ���U� �����C��[R�T59�#G��]�(Ư�Q
MH�߹�T˿�_����?�Q+�q����^�ݣ�EH���ok���G
j�Bʌ�k���rk�
�U"WN�w�4Zu�j�2r�M��EY��� ���v�pUtj��%�ɶy73�G�]�)�|�H����5��
�I��xݐ���0�)�jԺ�[�`es�)קޭQL��|dI��%�?ݫS`)G&��׃08,��X����OF0خw�H���Xn�Ek�
��P�e��آ<�!/Bq���@~��I�4��Z%�ׁ/���Ŝ[�d�=O�ĉ�Ï�Ί)�W��-.���"�'#
��C�o�q�($/(�A%��e4P��z������F�fyR�y���),s����γ�;��X,K�V@�<�1+�g�r� ג���l����}e�KUfC������@����K(�K^���?��S=����2���ò��:6�����of0��Q�f�|�NV�u��P?�J�E��wB�8����rG��s��7���ϼ����{h��ZZ�n��������yB��ć��'�]<��tټ8��	=�)a�����03�3(���QM����)�p,��b�8��� �����Q�_}����"� vG�jܬ��2OYQb)B�zS�R]�����5$��3��2�Y]�U'n^xbg�)�-}�Z��C~^??{�+N����z3}����<Tm#�:2��b��&gb��PK   �EX�ʩ��*  �*  /   images/83339b9e-8b21-457a-a82f-74d48bbc839f.png�*>ՉPNG

   IHDR   d   A   '��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  *NIDATx��}x�U��;%�w �����& *Ui+
(�
.��������R,tE����{!�t�{f�罓��0�	��������[&_��w�i�9�ܫ@���h4N��#�h!�O���6d�#W��rl��\.c�P�Đ���[�o���P�i���>(*.�(�:u
999u�B???>_}��#����!��w��d�g��?���˗;�XN�[ޗcAu���>4��4>}�s���A|\4rs2���D�N���Ǿ}���PRRR�~�70d��ر7n���
��9���	I�V���cʔ)��@�JKAJ�M���5���Æ�,^������収������˪�SCf�1mҤI"͏ bӷ��f!��;��`(3 .�
��C�����5�:u
nݺUc�ƌ�aÆA�բw���3		������v�>��?�t���-FƭTl^��>���t�P���c�#��/��":v��>�l�0#_�Z�]w0D8�OT��Q�F㡇����&pr�Ei�!R�q]<<��C����#HL���%_b�c��H�ӬY3���������8w�F��^�LU���lٲ��F�>}�����L�?]�tARR��D��� 11����ڵ+Ξ=��j۶�j���U=�w�^8;;�^�z�~���͐���U�V�][`ێ��)���E�O�(�zw��((+3��˙������������!�0y����믦��r�X#Cd�g��?��SX�|��l�צ��������Q�-�l�׽ۼi��+�by�"^x�E̙3[�өS'|��((0}x||<���� 6jԈ�QZr��m\�tI�]�����`�СX�p!}�Q������V��'CZ�n��5j�b8��x �����M�6U�\���f����۫�|�._�Gn^a�5��t�2�M��l.--{5�e�+Q1Ɉ��j�����₾=[5���2<6�E�ڵ�b�0t����tUeH��Ə��#���u3_� mnaa��^w�I���<��̅���/O���3�˚�5���~�7%�X�j�w�L��$�W�X�3f��TνH$��k�Νj𢣣�4�_~A߾}�V%$$�{IԀ���C�b$5�G����UZ����M�6a����t��e��)3t��5 �:O��gl^�����?=����[��g�+��ps.�j5EE%�����ۇ7�޻{��8o��z{aFWi�@u�EM��kѵc��i�"��㓧��O��'f��/N.ΪR�2QVj�%64���[�8�.]�b�֟Uc�f�B@@�Bg�`��S�⧟~���#ƍ���O�FiW%���ܹ3�]�����5$<<\i��ŋ�&мyyy)mb��8j۸Wt����������=�TaII�?�]������O��w�s熜܂+%�es=<\g_��B�N��	0Գ&�4���P�՗Q;d�J�Ҕ���-����0������DH���۷sNx���KdAxl���tL�0A܀����+@�ҢE� J��ٳ�e˖��֬Y�$?""B���~�M1����W�\Q퐙d$��IS��xNP�mۆ?�Bڦ�$���E�b�0m��Ksߛ��[���s�kx�����{�hoK��;����������{�X�Y�!��A��1�3R�$�Њ�ɭt�%[�ڋ�����i�N��A,�Ar�t�@Ϟ=q��qN�O����o��6lؠL�%ݼyS�����L{��:0��իW+�\Pc�L���	/��������Y(.)�`��RR3�@��\��^���0Rh�*XU�98:�N:ĠM�^��hN���t㜷&H�6X���v�C�C
���쏘ؤ�{�\"+�(�ڵC����oj?��]��Kt�V�� ;N ��ѕk7��|��D�&K+�#3�za�A$~Ů��Č���;ڼe���#++���2��ɍ�����/>�";Gl�����v�� B����v]�c㦭m��j�J���y��w����A���[�(}��ӧ�o�O�	:�N�:}�%�͎���;yyypwwW�6�Q\���Y��#F����������|�w3^�B1 �v|}�i��*�O��_��JQRf�Ɩ&�*Y�y�DӃq��f�i�?&.�}a����tA��h5HK�U�J"�E�2�Yy�b��e�NV���ٺu����8|��r�DYDk԰aC�9sF�:2�E��~�w�ׯ��:AG���ѹgee!88X1�h�ϤH�&���"���g����^0㨽��8{Oe�=��de��`g;Ⲅ����d�-���=eZ���hР�kI)�	��Rl`�L'��@y�4"�}����130��J��U_�������c�̙�aֈ���!�$��)��^##�7(e�����I�QԠ�/�?A��[o��5+�o��>��6;EP�wl�#K�,H�D�!)����sF����3��Wm.k�̗���e������D�������r��Ek4p+=�.&a��4�ٳ[=K/�L쪣�'��Ʈ}�*ڦ����j5�*,o���5"0��$�Yc����	:y�$~`2�/Æ�KЪ������L�V�Wc�~\���"7�5�>;��o��!���&>��>��y8y|��ٰ��h������?�U��88=�6X��ҕ��b��>��lN����3���L�O2�L˖-EvN6&N�;�ُ�'/I�PJs�-.�o�:�M��+�Jd�W�VG5��ɔqO<��C�`Р��SXT,h��l�uќg��73nVz�������[+�\��[���6�_����7����^̫�d|߾��IU�*YK.*dD���Qll,�H�ƃ6�g�p�)�P(�a�v��p����	��G]����O��  ��1�����ԇ�J�T0{dTJ��z����d&I�0.]�W��"kܸ�u!�'���$)����D�&��;	���jKw0��F�4T�����2���E�7F�	�֭��g;�����䌷��A��#X�v%.
C�^�V|�Y\�9�&�ٹSS�������M�#>(YL�^T܈�����s�7Z����V�`��^��7�|�͘�~�����k�A;
<���S�����$�׺wig{�&���Wga�uzswwCw0��=//G`�	�$'Se`��)�PT\RP��2��]i�|��E˶��wɽ:���'O_D�H{�h�N� ;{�����N�h�K��b꼥�I3j��:}���3���I�C���ʞ>%@�Μ��ҩ]�t^X��ؿ�^f���B������ ��w2����}E���jLy)����=~�t��F";�8����Q�e�L�Y�q;>Z��Ԕd\�xFⅆ�'��/^��D;j0�����X����1/1ԥ[_t�>)h��W�A��#��	�����(4���Y<2�Y8��b��t�\U�@```E�.л��;��_�]�Ǘ_"XN��Qbf��01����psu����k��8�e=J�8qFB�U�B�/�1�c��_?�j�]{D�mx(z���۴a)9i*�ИP�N���SڦE��H�<��k�������6�%HUflæ����兵�) ��냟���T�g-k�y��O�p���9���%ތ��G+��4������c��!9E�vT�	d�4XL�s�#ZTycġ:w�ĉ*MN��y+qQ��s���[�X�ɧ�J�{q�I���pr�8�HI������!�s���E����m�7���-��2?�Af`j�!��,�9�YWz�!oL�����ƻɱ��by#r�j,Ŷ��بY�9x��ء��H}lI~*bN��d������cԜ�2Jr-!1C�)�<sA�-!�����B�kRS"�fi���L��>�w%_Y�x?���q�&@՝�����W�Іɪz�գ��e��1w���U?��������NM3�"KSV5�)++O6QX�`΃Qh���Ei'�3��<=l}���<m96�뚊�w�;���X��G%X������p77ԡcO��uW���d���$��̺�"��r��i9[Vq?�*�S�A�,!5]�D���q��i���`��#�z$�{�},Y�G����h�B���ͫ����\UP̺���[�^AE߫Pk�׋�h�`Ҥ̙S�_�>2���A;C��yJ��-0X��1i���`=�ή�<g��̙�z���qèQ#q;�&���_�,�+N���O�6^�L�¯�Vj'$���:��%�~��&� ��'"�r6o�U�D]ށ�7U�Bԥ툍�"~-�~Y%��;bb8u�Q���F"8�+�<T ۻw?1��x��Y*��ƌ���Ʀ�W�a��>��o��ݻ�o�0aE���0�A!��4�A�_M�jr�T�8An����T:Q\���^cQy������)�w�S����.���8X�b���Rq=�
b��U}		iʄ݈�Dr����W���B1k4sj�NG�+f��D�������
�^k B�2���TP��.�w����Y�b�X2�M��u���ݍ��/rԮ�wb�`���oW���jt�T1Y���CZv����u�pա��\�� גno�;����>@C?�*c��g
�����}�w�`0���ZM��?��Q��歯(�X�a�����}��">�f��J��2e��ଜ�AOu�є!?����A�Ӎ���>d��Y
w���1�����VX�}�*3���8g�GK ��9�̀��������F���ġ;QT�(ݨJWCB���hP����ExSah��r�T|c�����)�S>|2���GTt�z���T�%z,��U狊L"�����9�кec�m�T�����OSS,{�K�2�6;�`�K�Ȑ9�,�f��r�u)�fmԺu?Ht�"\�k�OE��׈�T� &�f<�wU͘���
�~o�E���0sѵ[wU�ǪKrt�Ep#_A��0�H�[$�":&�#��7�dD�@#�#q����OO�V���?�m��/y�<�2]�%�������V*M��H�p"�1ʙ�t*��	�����M��Ŏt��R"%�B
�n#;'�^f�;�d�FANK�� ����@PkR����Uk�c`W:�����6l�3 /#7q2r�fk	��{E��Μ�AT�:��;))g�+*:QM׍�>c�{����@�(��C��}�}n4~�x=z���Ř��}�_���9sZৈ;RPm��=�5'�+�G�����ߟg�@ػ�@ڵi0�G��2���M��W+5;�E�lÑ�WQYF�5����ɂ��WT&"o�������� v�����[�����`�r�  M"�W���ե����w_9RT�#f+���[���n�$���T�!�()HF�`w� ���"?ARf>��j�v� �꬧=�	�9R�66��׿����=*���_�asg�Ȟp�l '�����Qi���_U�Nm�bh+*���d����@^_��/��C��)ӭ]�_��S����!,^hԨ!<ݝ
ar�ێ����@A%-U"QW���-�˭�� O<1����W�fȸ�\<o�֑I!���C`1w��6Ĺ�1w���������P��C���pķ�?�6�կ�o�􌳣ڶB���h*�\�̬|1��T0Y�0��N�~�����s�U�]+�"PA��}�ȑ�$�uC�fM)�L_���p�F�Q*ǝ���zH2ea�Vl�(P��Pj�����b܈M��}>�ݥu�"D^ꤣ.�ˢQ�W���4An9x�q3f���dA)3�ο>8����-
��gJ4��ν�ɩ��j�ў]�jeP�E% 9%�����-���"�:B,�z{���Ѷ���0�v+����ph�Uaa�*������>�l~�%�>�N���CGbȠ�X0�3��i^|�U�S�nJ<���� ��>m1*rJm�g�B�(Δ���y�q��j�:|��G�g l%�/c�w��E̘����J���/Ŕ�Lq׈�ͪ<�<t���ml\\�]_�%b|�h�x��C�PkL�i�pS�}�������F�����K�1q.\�UZ��,�I�D�&m(+V���5���ļ�(R�
�������_W�{,���|�9���^}�m$&&)��<�����d�||:e�vX:s�p4
�/_���)i��e��^��e�$���q� ����X���7��R��4yhѢ��^�xu����-��)M�a!@Yi!l�U�$_ ��t��Lp��H��Q'ƟǩC��Wo<u�{$�������B:��h�*|�f��&?Fb�������DZ#��H��T������)�}u����.g��i�0N�믿�P�����駡�=�(@ki���}s�Sͷ�M����������K�n�\t�X�r~O�sY��DF���|zF���*�MEq7R��~g�$�)	m��VZ���젯�/:u쀃w!&6��3�7��֜5��U_'N��?�����JcSu��i��DSN!�L�����h���}x���|X����;��e�݌��������\B�;�3a+�L�i���g�a�yʟI}z�B���)'��m���pw��a]�a����)��,����N�w]R�&2�ı}��.a&�Զ�Y�X�RU;,���QVn�,�:� h��47�%'���k(.5���	��5����ܜtU4���#���UɆU��%��r����J>qxp^z�e%�bv�/�c�>���?���yU�Ú&T7�X�����Uo'CXm��l��\O:����Ŝ�����л{Kx���hq?V�}�]�TQ�sw��}�=�C��"''��<U���`y������Mp��	���µ��ѤYc���u;A$8k��XX1�K����غu����*.�G�bj���>�����jKL��6i @!q7�,/�!C^�	R�����_z8x86��{��(�R"����,�SL�U�Z�i�k�$���.U�Yeʗ�>�C^�Y(.�f�e�n�A��pt�A��O��p��Q4p�ţß���^����rM���p�,דp}bm��\/��Y���DKn��EA^ܝK/��	.7����Z<uEB�_��A��H�'s��Y3,pt(����th\�[z�{]SU��ұq�^7V�M5�*=c4��T���\2��Ѡ�Q9e����34YL�ԅX\�r��
Pc�P�:�A�1}~/�+���z
T�J���	*_��Ӂ��XAaa����~��6�ɪ�����j�MUHbd���`��x�S�`A2a�QJ�N��/zU��,:ȹ�41G��?�+��E�?��b�q���;�$ �V� ���j��7jJJ�<s�.Z�v��B�bE}բ��<9s7�B �=s)pfV.f�[��|L����BB�In:�<c>�^������ީQغyR����ŕ��Yt��{��;���~������=Y���Ж��m�=EE��&=�@���ΒY#.�{�ı֊Μ9*��ة�rtb�0�� o?pZ��VSޑ�k?
�t*ٲ@M�)�#�Y��5�\�2�vd�.Hd�j�ʊ� )�F�_�E���r�ڊ�TVMǛ�G鿙X���!m۵��>$�|}Ȇ�YbI\%��ǟ�����c{�֫T�\A�dɗ�VPQ3>[��ҔԴ��gr�ws��������Dܘ����-[�T�\N��7�B�lnP`�bNEHH�Z'�~���ps^e��I8zd?���μ�
�T����F�����|w+����p�z�Ih�"PTЇ�,�&��0h�D��{���M��Y�W��V����#��&�8�Yٚ>�j�rC����ue����gJ67+`�&f<��D<���V�|еCCeE`��0��v�-rS�&=;u����U�j��떋B��~+,*��Pf��h5N��zy�O�������_�U��Ν��ݻk�y�L�\S�:�'�8�*Q

�^�K�f����ի�j���GmNP�US|V�sW�nݻ#33K��L.�;yt��*\2"O⩅C��$YZ�&H��Nl�<hHJZ:6�]��>�X��X�G��n�D3E� 3
�?�������8]auڃE�k�lm����40b�*<3e�U��|&48@!���س�MN�EM`P���6��`��;�iGG;�����tUp��l�6��5/��ֹ�@oWdފsh]SYNԶu�B��.�4:�wR[EEG�sǦ��p8�Dm@S�L�>Cm��=ńi��%�����Ԝ�V���NN���s
^�������X�x챱��֊!t�'��Vf����gVTt�����uqqD�@_�tQ����nN�()�Ę'�HO��I�+A�׀�m��/�@Bbz9$,B��!�4n ��Ӥå�����n/�8_��?7u(�[(c�,0�1�Z�]J�	c���z���]�:-X���߫!9�O�}�v�q��N~���Ɓ×�u:a�sS��a}��#)�5>p����Q!�>�>A��:z�Iul���l�����Wa ��"D���Ҥ�������{�v��tss7-��������2c�K�+��������mϙ��u9P�3<.&m۶�`5�_�62�/]�7�Ip�&��7�ޣ�7���c��"�-)i�������}��aݞ�]z���T����$�m�>v�TϮ-��z_�o.\�ՙ�}�&b6ZC4w�H�a�����4bX�&_|i��rqv��Gzp�؏¤�"_����u{A�afy��C�"��o<�w�lԹ.�N�w.�9z�T��m�n�Gÿ�;wۻ!�nb>yob������Avn>�����)H�-��n�Q�!U�o��(tJF����⠸��%���r�zi4;g$u]4<#=K��L4S�&Nm~���J��l���-s1��ʎz���Y58O4$��'�����������dc���~��l�wlJ�B��saM�33$��z������{�hgo{A�Y-�������y�b��g�ۦ��oǱ����� �%�k��lN��`�@|�}ש��BZ��J���,�:���b���Neɧ@��mo49��������!�DZ�O�yN\��`�írQ۴Ƀib��C�h6�z[���^>C_!���������y��mX���0�1*Uo'>`�A��7�-3�9�&�ζ��
�--����}�8����`�G���'��8�Pa�5/7�k��p&-I�y*�G�^��f/���x.��}�A��QX4-5���5��6��r��2����7q�/ry���1��Ix������������8��u��--3VLU�c�ʐ(�Ԑ�R���E:���3��9*��C/L�
�HII��:��÷A8N����&t����u��﹩��tU~~a	�FsWsj�{Iqۼ�{��'�'X��d?����j2�L��9�����<r�g���2أ22s���A�O��WW1y��o�mD�ݵ�lEJ�ol�W����¸t���~ґcW+;i�<T���[�e��{y��E��סc�����#ѭ[D]:/����Oi�`ow��0k���1w�{��TBiYك\ӗW��[6�y�J��*CS Ϟ9�h�\����s� �uK>{���Ξ\�MDQ_zF� ��%d�}� 9r��1����mx��>o��g��s�ڒV��#����C�&Ә��x9"UB4'NG�5#�o������R2�1��f�L47�/������{�U2cߡ��+���9	ʚ�P��Ֆ%9~E�q�i;���ahb�@֟U�5��|�ŗp0�MC`oc�����-���8q��U�\Ѻfb�_�};[m�p-�y��J{�Ve7$ٷr劾˖-7�J���,v4Bl���f�zE47b����)R��6m�C1�j����+�0Z�`������VE�9�J��\C�u�խ�bތU.|۱�l�z{�P���
���Fm���ɸ�nG������ܕt�Ͼ�,��N�îDF%���x�>(߼@\���s�jW�ӹ��D�[
���5ޓ�/��3���v!1�����Z��H���i����|��W�Q����ر��:����tt�ď�M[������-.qX�j5�\�p��5�n<T@��KW�Ծ��>��R���;t��M4�8�o�E,�ھ�\\8gݺ^���ƿ�����F����C%�eAwKKL�G�6��)S�����؜)F��+1���ty�r_������e���cz�ʀм}�S4�yQ��"a暩���u(w��٩ϔ�l�{�ʝ��<]�p^����L�;�ѿLW|_�5e�c���K��C�o��fwv���=S��n������3@m���koTJp��K�f/d�!L"2+\W�p�ivho��,�At���}���!�������r(<2�nw1������)S0l�3���.>����{���ys窝��VJ2���Nͫ)�˝�O��z��	��!\ć�u�(�V]ҍ*ɭ��d%�ZSW2k�#��\7hf��s��g)�0�s�<v$j	��0�QS/Z�˗�}�J���!�u��o�IN����֘A������S"�e�e`G��e����?��s��y�c�꾑��o#%��Ɏs?E*۬K�9'�v��U��9�es���ՕhF<���?��Wν��q    IEND�B`�PK   (YEX}[֤�n  �o  /   images/8a867033-535c-43c3-abf2-d13f5470b1ca.pnglyuTN��ݱt-H��ݰ��t�4R�H,�KH
�KKHKwH��H�O�����;�3��̹s�̭3Q���8�8   _YI^�_  �0��H�0�uhv2j2 @m<�%�?�E��  g��T�f>�G4E("t�\�l��,� ?&k'͏�w&��~L�Lb<L>�` ���x�E�W\�G��Qx�?n��[  8_)���zgu('��ryDQ��� ��X!�\a�F�z���z�6�B|c�IW�]r'vC�:�m��*)3Z=U�W���� ����TJPRс���?���\z�ܱ�!<BiEy_o�浇��c�M��"VE�*S�2h6-���B�d�(���OS�����M|$�0������^�5�me0X3	UN���1܄ҹ���H��\�L�*EѾ#Bfm;�t����]����t��=K�mSBx}�;
�e�YD�i�����?et�#��өI��ͅihh@�NS5g�J5��m�GoB��a02�Ů_=Ð�߆E��B�F�>���ȝ��V�*d��2�;Pz�4>�����AȐY\�rG�l&���uێ���H�6m���Z�^��A2$��)�Q��6�e|R�C��n��t'�C�=�8����ك�Cx�mr$4��k���6E&��4���Wx	�%x���3�^�p��6�)�b�;a˵փ|5����9���CR�JR�X٬���C�5L p-���n������~����ӈ6����T^ff"v��c����F���ɚ���*��%�ٸ�Wp{s�P>�م2�&��(p��f���5G6!���2�v�y#�7��k|ĹEЇ��V"��^w����I�	��(U���֓U.��I  A��Ƃ zm���g��C���L���u���ˢ|�h�FC��Ȱ��@� pW"����֫��2�?D{�h��sV3Es�)/����Y�V��X���6[������m[��t�v�}��8jZ�l�:YR6OU�H��y h����7��ά�.��	T����������)�"�%�Y����䰈|��5��vYg���.��1$� ��J�6'�+$h�F������Cى, 4�����g}����Uo������z������ ����n)7z'���[�A٫[�oM9�qd�9���&��?��-6�s�YkO]]B��B� f��ۏ��0_���঵�����+�UԐ�K&����&�MP��d�s�d�Y��5�<��:���5�Kź�+ǵ��ƙ��t�":l���E$�.�ٽ�x
�ZK��4�i�����S������p4��}�b��[:6g�&�D�*�G�G��y@Gù�E��K�w�9�v��g��?�]�(��ڍ��[�̡G5u���j\xϧ�u2TH�l1ygj��c�#�ߚl�[��B�05�r).X엀2$]��_�Ȕw�&�t��	�a�v�E� �0eu�,3���^	�5Bٯ�°�
pL�/&�)\�9h+H1�\:G���ѷ�c��S�8���fQ�󢌼�jV͹��"aHlI��veʌ"KQU�L�Q����]�&j���ag�d�����Ġ��y�Ȼy�:��N
�`��]����0e����5?��[�R�a��_y_�"z���C v�d�X�8�����9�@;�whbl׿gþ��r&��R*��i9*�����P�m���稩�ѓ�ѭ ��ZC��:s�U��:��&	4�C�g0�� ��'3{�}@E��
#�b�ssso20b�H��ѭc�M���c#�C,^4�d��PN�P����?��KKmq=���8��U�[Z"�e�V#T����G?��D+��|�S@�����x��#<ZѦ�Qz)z��5A�5���O�:�D�5N�<�?E�zn,R��D ��ш�Ӏ�k�;- ����Κ�X�����m�p�*&����EQ}�����wx�7�����S���%Q�JQg�<�����A�w��g�i=��]�9N���L�R�@6��'(��y,�������2џJ%����3E��&ف�v�ghBo�=�NG>��'p��V�8�e�!�HG}@R�H !��L �|��/|P���|6@a�N(�8��h���"ь��f^���W��?\��`��D��v>��p��W�CY��D�!k���M6W���m�/�E:62� �XM�֍�-�Y�WE0MJf/`K�%������I�,��\ ��o<�ݳ�׸u+É��9��;{�EY���}Еj6$/q�?���6I�2!�4&I�P \�eg`�T��h��,�AĒ� F�?�@�/�+͏zr�{U�Y�}�^ʊ�?�9 �,��/ሟu�I�o���p,~����������A#�2�`��m�S4蹽�e#�����5 �;�so���9���5���6��}�\�����cG�B�r��L�>�l(����g��=���.����������F����}F4��
8^��:f�K�3_=�n�q����O��4��E�V��P�'gι!���J�*�^7�����G�f������P��y' ����ԓGnn��Tc<q���ǃA�'���l�ƒ��|��T����7�0�H����NTA�{U>y��;T�,��Aq� 5W���.����.�zc��L�l���-��[�_Г<9�����mއŋ6���������֙��j�J�o���
��	�R�%6L��pGA��������k�Tx��h�a���i?������G�K�H2:�n2�g�j��e����P��iȞ��gv������f�:x��@D>�c����c�Sᑨr/t��D�������F�����:��Y��kx:r�G�@�h@�Y�k{�b�h��uI�F�B�W��.�1�5�����Z_@�ɡ;�ŀ�Vb�WO�o7���D��2j�ġ��G+���E�"��Q٭O���)�o�<2��n�����8�%�#Q��ph�ȥ��_A\)��B�M?;  ��όD1��ҹ��:w�̳�~Iz�����_�wuIg&�� ��Iy`o�1��ytx�.9^���9rʇ7l�<���t��#=���ü���왌�8�T����"	Q�y��շ^�9��X�w󢑶uv��RSr�b3����v�Uc�W���v�R����y��պ�\�~q3/��S11����,w��R���G� �-f�ܘj������dy�R6��eg��{��?���jE�o������>�)�� �:*�L�5X��<5�o�}Q�����0zf��~����]lp(��>v�n�5�>n���Eʺ����jF��w`D7z�v�CT�g"֍�Q?�aG�U���3ZFY�5��RU0[#�D��E��X�|��?��!�h\^�X�)%c��"�!��F8:����_O����U�3Gf�Ip�Y�O�`O>��l �C�I~y:��rUg 7	��s
�dg�E�5g�3_��J���{j۝��Ϣ�0?��
S|evN	�u�IP���ݝ��D: �gc��N�ݢ��GY|��d�����dc�����*�F�F2nzj�ޒɮ���{����A\!�_��HΕlzV�_�7$��!C��6_��\~RW`�h��������(�K9���(%����r��t0`�Jȍ.P��:l��d���%��!�㧙y6@���2~���{����1�I��-��JD�y���I�*i�����J��^Ɨ	3�nFݝ<���o�w��>��a �d+�k}�=u��a�i�{�'�6�R�x���B���>�T�	K�V:���t}�S`�|늧����cǕ��O�K�.��0�w��(�c� �u��;��������5����^NB����_�?~"o��Sq��<b^>�T������?�GIS��+=�w�S;�~�&��ˮ�}�8h3;$��q�|�y,V۟�������f��Z§Sb�����,�G�Eo��q��a���1!xp�3���.
���5�*��u��By��N��pQU68���B�ސ��vhdj����t��̈SeH�	�p�9/]�����wQ�#O5]cߤ&� ��	���$�(�G�4� "����줔�[�p�֩+�
��"Qh��d���L����#�H[�Kt��� YMoT�|��|�M�Ib(�N��ZYd.[���ss	���~�_E5^��7R:��$�|A\
���m��J�X(����D�����j/�9|��RtqԘ�����"$�$ ߷�~_p>��� �lyp��a@ë��>�uU[;' xG8�꣡�>Υ�~\��x��&�a����d=���97_Y�D��G�G���g���U�6����O>7�^�w�|�b����>H��g÷f��dV�%��;tM�E�z�XҲ"ro�������o˿Z���>�
w-
j�� �<嫺�R�y�����@6d
�/��5��Zzv�/~3fs����ٴʫ����x4�f�H��oJ���&'��S�}Ee��f�]^F����҅n���Hw|�� w #(ѭE�bs!A���H�5��E�;��zjꢔ�J�P <W�LG.v�>�#-Ƙ] ��c�
b�`��z�d��E҄zjo��RZU��1���"��4h*ӌ/,��X��?�#������٨$s�=a<��y'���������g�#���?p/P�\˄?�{�a�֭��d,<8��b7�ct1�N#��6�ر�%W�����ݡ�-7Ċ�ʂH/sDd	��&�UE��qp�bI?��gK+X����x�L��3U��"�҄��Gs�8�`ѕ�}Ӊh�k�"A���
�&a�pY�/��fQtD��=�V��_�� ���"��ݶ�����me�6xy�Kxd1jz���l�ln���0�J��6��L�!"��Lg/r�y�0�U�L
1w!��g�*�b��bPM�>޲o
�)�މ�`�ؠ����R巃�oc�ֳ�:��{�Qc J(k�7��G>��u�K*�+IZ� ��Zm�/������qJ��T�RZ�R}N]4���|�8晗!���e�{B ��䳲L\̹q�_�Q�}��-��&�'^*b�r������@�-~N�7����?�p���b�:˗�:δ��]O���5�^S�,���g�!X�Wx��g(6}����đçe僗K�g���:��N��E+bj���ȼ�<��,z��U* c�'%���D|_�d�!��匚��3'��9኎{Nzpz0{g߰�5\A���w���搱�x3�$�4���~'�$�3��	BXmjn��>=�P�{t,�XIc��b|�箬
�PO�������i;�4��}ޫ��ʎ�|gʤ�/���(̲F�G����t����e��W�X��,x3���5־$�{���FC�K0Q8��*.��ɭa�OC^i�߯�|ϷCϫ�_%BI���h�.�*'�8�-�HE����Ԧ�E�+z#�u�)$��&�O"u>��a��z�ⱳ6��y{Db���1)��JV��i������j<�?r�(�kS_�S���\*��a�!�FC�R)Ѱ7�0،?�ĜKټ�^��6�$߫x�����⮄�ǋ�j�=!��ħ�����x�eO+,�ڏr!���ݙ2�J?K�~h��	,���>ޡ-�=a��[�Ȳ�G�z?1gV:������@G�|�-�)�s�
�9�?��`x,/�������A��wx�wk���߅�h6�1 �d���u���	�m��8� u:ʁOi�&��x�F�g�Xg��l�*9y��E�
>��L�w_~�e�z���*)��x�n1���8��	:�U����br$<�V=
P_�/r&�:Fd��R]����r�S����7ݔ͛*�����CC�!�cV��'Q�w�%:���o���{hpH�6~��T}$��\�*l�[C
:a�J��3Z�9��H���SHP�MO6,�3Ǽ��R����A�s��O���b���ݐ&��mUns���/x� ~)0v�wwz�a�n�����_'LW=�������cfp1��#-�D.k�����e��c�ɸ�X���L�b7[Ƌ	�g|�'/�~iAk�$����B�W(NY�J�ÈLb� �5�1�#3p���qɓV�vT[����EM`֖����_|���N�Mf>��U����WǢ�2�~v�ElF]���W�G�>�wߩ_��˚)$�EgY� 0$�)�@��n���Y�g��o����i�X�DGܦ�-����7XT���r\k1|^�B&��@v�>�~���$�J8�Z-���VW�����?E5�X�Tw�ub�,[�E�k)i?lÌ�_��j}� p��t�Q�"��y	WN���u<�/>.d�[4�Au6˕(Le!�Dt'1��h���p�e�"j��N,HS��O����f�-��Y����
-��>�%��Yo�hC�$�H����I��DӅXW<����Pf���v^�����T\�y���␠�
p$fG�P�cL��X�K���K�m��^/�Uo��=9Zԩ�.欰��ט���@��MY�1b�s��)����g�Z�@�R}fy�SVW��B�w�,	��q*	}��?+�-$f_������y�;@�Y*�Vם�g�-G�)_�{I&@DU��V�8���jTtc�F�<l�gEj덲>�N.{��2�D]~�̒�-��F 0~�[�s�n�C��󴥒\|�y�< ��n����;���P���__s·��E"7��	���?���5T����{'d�P:������n�+�0���a�O��$��UX�O�+3*>
7Y{9:��
M��o�`j��5����HU�|�̨�H��9��T���f�U��N=���ANror���uu����zG#ԗ��8^-Sф`9�@�bcڷ`�7TԊ�F$'*rk�Rw���c|�ڻz�*Q}��e��1���n)��z�9����}`Ú������cH�\��D&�7ٳ��Uk�ߞݞM�}o)��m&����h�km�i�-���p�|�n���b4~2_k�D���o�bd"�Qx�S��\#�3a��nMCa��ce�qs;�EQ��	���Sf�)�t�F(�S`n�Ui�Ȝ�s N�v?\ ������1I�c|��`��G���H�����r}�tZ�A'��`}*��M�M�e���Gr��2;WT	W:�k{�S?��BK=�Y�c#��mF,����B�&��~	`��b�Ϥ!������Q��:�)R�tH�k�yXs��yϤGr� ��>U�;��n1j�e���^��$e�1k	ǲ�N!����X	�3�w�w^��h��N�xQݮ"� �C����F1����(Z-r �I���Ç�R��!��:1p�*84��|�,��19\�|B��L�Q��~)޳�EC!�	�*$�=f)��b�O<
����f��<�Q��Qٴ��s8&�����s���p�>����L��Zx�'N$�fY-�k��\'D�T�*vw.|�>��l����.6�+���[�@@J�����݃*^�`j���Y�}v��<��"�I�Vֈ��L?�$�n"ݗw;L��|�{�ſ:֪.�	 ����$:;�7�0Zjf0b���K� O����a
�խ�`�=w���[KD�x��]�^=��R��Wʴf3���`�e{���A�����CO׃�c�>w�׻Zo���������M�+��::�0�Ї��Fbg��1.Z�3]��7f���z�,8bZ�;3���ުC�h	��(�n��	�u��h�"�,�Rzf��7�_��|���0a��`m�.2"��ب�NNC�0p#7���̝U�Ʋ�f,]&��rixYm�Q�X���޴(���X0�GY6��^sH��EV_� ���Y�w�f���#����&]�4�Ԁ�rl�g,��
�V�K ^#��n�A��[bʒRu��F�����&i��L	"�VS}�����I�f�/G�seÚ�r��vP���Q����~-u/�H��(�}C���� �<k�Q���Na���~2]"���^�2�/�"�ì��˷:��K�Ĵ��%䒂��Dt��B9�Nn^&�V'P�h%1=G��Ce�lc�?�|+���|m�z7=O�|����韪�LP��D����������>^>�(fءs�S�}+<�c�	Cm���B��w�bz%Q@�N�����b����T�a�RYsʟ��h?�c�Zܩ2kF7+=P�=��`ŀ����@�Q�|/x�p��C�	��g>�&�C�M��]�L�b�'T���Y��B����*q ��xL�&+隴���;f�/T��Uz�m�{*2�N��J�[�܅DX�-;X�`_�|Mrɯ.��v�os�/�b��_+�x�q��`F�)8u8�iq�A
���^�_gB��5�5�8�� f��Y�a��.���G��lO(t*m/IC�7/��V{��{OBQK�/sR�B�<�#���ZDH^���./B�`�x	��/>��\�$o[-�
��$ ��hk�r]�}��\V��=�8�_hꎟ'�/�s޿��h$�yk�x��^��l��r����Q��G�U<��Lz�d�l���ě=}o	|ju=��pha����a�17N�5�+:S��璀�8P�n��e�<��Y�W�pU�N��*Z�����B�����]�5<�)5��-
 �g�R;^��N��Ǎp���g�������)LhS���؏b�b!�Uw��_�c�{A!�;cX��[�m�����`�� �\�O.��_��s[Q������>E�����h!��y}	�}�
���x����E����H�w!��֐~�5�*I�UZ��w�k�Ǟ4������N��v�2�K���@)�C�B��mb�Ⱖ1af o���}�@�sF�v�0�D��n������Ž���^j&�|r-�0�}�F��r'4�6�ϓ��"{[��i�Ns��z>}i��P��O)��.��B�����!��G-#�e|�a�q���W�M��:1&�KG@�����g��eW�>�S��ŕ�[<����U��.�`#�թ�ks$4X�?�1e�D��hEd�\|�Ծ잜/����Ec��&��:�ͰV��Ӕ(j��7ɖ6&[>�o���l�a������Pz�I.�?a�˵p*�X���f1m�R�U�y.�\��vz27ӣuNVW�9T��@��9�ځb��.��>M��������9N��_؋��B�/wv94�ܲ)&���p�Dp��g=`�-PiF-E���Ub�)a`I�5ط$3*�'w�MVƭ����c�B8mޞx��P@Xwf(	���B�g� ��%dR�\a��R������}�g�m[����R�/^�`�	񓱀2tE�����V���#���X�����>��s��1����v���*q0�1�����o�Aā��#��XvX��4F\ߧ0l-�o�S�X��� ">�vd=5"�QtY	������?���C�,�[_�:θYa{�/~$�3,sii�AԌ�G'ف'�x�����k�0g�<&�fLx0���%�"��d�B�
O�J��S� �ޗ�~���g$�m�|��4�Ta����k,�-W' ��%̍\�q�̦�5x�>\�~�����-0�&�w����G��7� ������sE^x��v(��ޢ���[�1�����&���vF/�T�R$${u�7Ru��}b_�t�r��C����Z��"�E5��ς�Dd�i���g�o��`�S߻s�� ���?T���z�����@�D�E��=��O]�Xg���c_�p��S&yyOק�+�'��G?���qY�=��n$3IT[�^^�,��u3M3�0ʁv���j�m�l)�� �� �uI���c�|h.�$�Si0�3����)���4v�N:��_m_����5X�|�O8�i�Ҋ��7��t���o���~85#��Vd�i7���/iP� K�t�i�?�n�����'�������0�f�OW},��C�T�� W���zr$֤dt���o��Yz��C������ȋ�#���Dû��NGŝ�����V��Q�u���b��d����SH2�ݘʣ ���,"s3U��?���я���j���X��Q�_NK\���0�Χ�s��ɲ��M_kHL����a~[��Y<�{5+[���й�q������.{���ad�=0ȀB���I?0PU]cZT�r��=�y��H����y��6�$�s �Fl\H#i��י����CD-ۑ��9_�>��!�A�>��m&i'�Cw.�@��-���e��Y�y��a`Lܬ��أ�Gc��ہ�PR��~���i8jw ������!�n�c��	���֧a�	�\կ���R	�s5��jdh^�Ɋ��H��ED^�?��fRRlr�;_�����k8����Y���T���D+���(wG��'��$��zm`��X@�4G�>��`M���z�$��e��{��S�k[���bߺxY������vٟ��Ml|��7�TS�p*v�}gPimPs���=��A�B�퀌ez�ܦ��K׏��ݦ@���-�/}G����߱��������S���Fk,�՜�H�F8 R���g��X@`s���͍�C������f�%\g�*��:Zf+!����sk�<F|��MJ2��ws7��Y��Q� ��pV!�F�
F�d�����嚄����$�O"׏�~��S]�8!au��������/w!S�P3&��) ����>����WXi�W�cqh����Hb��ն��n�e��-ĸ'3>��.�t��H)��,Tcuǣ�d�>���ƭ�;y��$ 
��Tﰰ���E��1m���s���p��������;E2�ǎ���a7V�!��9�yH��v� n^ ��@6�<�-1���kg^���ֵl�����ȗF؝湞;Y��׻��z�ps����<][W��(�B/�]G���È�:�Q �n�fu��e}���U�[j�N�TlO�X�F�_��F��HUq�\��� �P���x;[u�~���<��$�I#^b�0�
�Zi"ȟ�S��Ԥ�t���Gi^̖��dKW�4e��:�"j
�T���-j�ߵ;2$�Z��:��~m��<���k%4I��z`�����Թ
J�
8��3��
�}�f{�4F�G�& ��{ߗ��[��ޓ�Kk�Y{������|�\H�������/�#��T�-%>z���¹���ğ����Ô�W�q����UvS���P�$�*L�%ӕ3���v��v�QV�_�ݕu[��K����2�7�s��.��(��7G���8����uAI�����W
��@������.
;x��,Gy���J���x���1�z���xW�`u�n~����l��-]�Kf8�:B���+����m:;��|_/��L��56��c���٬���ֆcB�dY��ׂ�UH��'�ϼ�g��j��+;jj�7�U��G��j�O|Jh��*���++XJ5�TG�k&a�	�	~XB���~ʯ$��6�=B��`nA�ȃ����p7Ne��Ш`�X,�1�M�3���T��;I;�ĉUF2QnB�("&��l.C�����t�>���H��R�,�1���0:�,ʝr�Ce��e��}P�H� �O/���6�U�'&=#���^�U��B�:IJ�Z��Έ��N�9�2����K��'��n��L(5�������:_k{�7�ƚy�]x��Qy���\t��ʷ���PB5�8_�^3��W����� �8��vˉI; ILg�r�HU�uR�����+IF��X��gn_���r
��ꊋ���:�mBW�ǃ��)>����]BX*�VO�N���QB+���)M��z�0��$������HT��O�{�N8���wn�z���vO`,�Շ��i$X��^�I�sgh����i�%�a4�N4zJ�	��}���{P�αn���ձ�欈dΧ�Q_G˴A���_b@����d��P޾�ɩ�՞��}����݃��yi�Y�=x�?Y@a���]���7�qU]`�|�cY��o�r�*�*����u���|�_zg�B|r�ֲ}��a\�~���gAcy8�#��K4��BW0�r4�_�����*:!�
qѥqH��?�C�68��aڥ�ý~g�LTzܶ��O4f{m'x]�Uy��c�M*-��4k�Cx��;V#��QBsF���t�!zkH�IX����S������u(b�v��������L�{��ů[n�;4im�0��������V���a��-�"k�$�7���b܏�F$lqvR�6�m�mt�gut��vN$�ɤr����И��2��}��u��@x<��8�k��\2^;`��N�`�$��T���1���r�sE@<���am}����~)q�L!Y��&:�87v�g-cR��,�[�L�*_���x�d�K�h�2�AS��q0,�3�\Ċˬ��BL��1�C[�F4���5�JD<���-^��D@+��B��&nfn��ù����/��Ay���a4�f��8`�|$ѧ�R�;����M#�젌�V�(
�Í�jxٌ��c�l��V��z��Y�?5�������?]���w=�;j'`%���4��4���Mg8~��2i� �v���r��k������o����M���1���Ny;C��!#f>�W�?� �E��R���0�cSޜPr��T9�����^΢u��-x�xX�T�Z�]����'����4�XmJL$X��l�$����\n�в�k���y^?u*�0�b��UG����Ͷ$�t�=-�~��{���������Fn�~�_kJ�иUa116�_W�� PRj�p���4^H}�����E�`�Cy���/�iW��}ۨkAPO�u�-��/��|i��P�c%� ��G~�+/���"�S귁�煠�~W#7�B����#�r�e&�Pf����5��α8�?w�OA��2ً'���-���E���t��5����.P� ��	dBg��U��l�d������������Y�]*}:Z{�/@=o��n"#鉘��D.B*�J�6��ߴv%g�:]�S�ŵ��=��� ��W��d���&�Eև ���F��Q,�����^�U?q�<� ;�[������γ�]1��"��s�����l-m�U��6d��Z�Ϸivy���R�8�[\6
��C��W�!H��v��Ƈu؊���7��&af�#�<q����&c�%W�\��~�PTIԴ�;����+�����N�}2���=4�9T��lAX�쀍M�z���ߗ<�$���ȄP��If�Ϡ4�D�È�D����J;+(�0�W��a�.h Y����M�r�#��x�qnW��?|~{&kAԍV�yS� t_�������{�l��;��{�Ap��{lr����C��L�Q�u�+�Kz�1皴��Ϥ3����l?=0~��1�,�[���.�}Tq�Ox�ਏ�<}�(^������� �������:v��X�z4���~���I:Xoa�iE�m�	���Af6���iB"�q�3�kM�Q���,��Ҧ�M�:����yz����ar�΍^���#�����b�賈�Q��9ԃf�\^2�^U�qt���n�7y���}�e9��(ia�F�~�V��b�E��6%��Hs)�;�Cf첗�ш������v�W���H���E~�9C_�ޛ $anh�de���)�J�pt'B+�e?I1E�ʼU�I��	&�Dw�Jb�_tt]�c��Y�J���$�	/�/�����_m��it4��m	S��&aE
%�=ȟ�/�Fkb�Iq7G�H}
lV�V;r�0���Lo��y��Dڀ�t�#kH�F�M�Y��iS�92�������l
uI�֌D�}c9��n���=ɪ�Y�`��!�=!��껐@����]e=u�I�ˉO�c{}�����A���hƖ��8im���.�DEvD�w�u'o�6�s	v�O��1�>6��$��s]b���4�g̃���`'�#RL��p��~���P�I�p�+5�����
�>��,!��PAx�8��/����F�r<g���݂e�#�C<ʫ��
�݌��8����Bo�{�{p���v��;�ؤU�8V�K��F����;�%����pB�������V��T�ߔ���f�yZ}&]��+mA洮�+��lC�jk6����?���2;N�l��|����%��F�V'&[Otmr5V�Kv�o_�9��ow����* ]@�Y��R�����>��Yd�ÙJ}u�4���)L�y	2���~��;��>�͠�q�zQ܍Sne�0`�w�K����Z�����i J4�;،�θY��BFc0v��!b�O�Zc�̈́���x��`E{�St�Щ��gZ&�w[���-})���l�l���3�s��7�Uy|�y�Q��&������(Wj�iXW�;�S1� 4N� =��
�Y<t�F%��i�ӈ�#�ۮڲ���SL���%"�\���Ƃ��/����8�2�3q�&�^���S���6#Ѭ��� T��
� z�B��viTos���aZ��Wq�m�6@����CB��~`a��n���F���ϙ�ޤ0 o�g��W7ɫE��avW�&�$��
�'�WA��S��4���:S��(�QG�a�i�[mٮ~�F��$�EO�^{Rb�:N��Ϙ"=�xW��c�*q�g������r��.c?R��vʊy�vq���9��	,ӥ����Pzi�wϏӊ���ذ��	�G��lpf��T�Y�Y�}W����$�*逰a� ʳ�
������WKzZ����4����[�=NCT�Y>UE5�]@�m�y���2��K��ʒ۬u��c�wI&xr�}SÎw��4��
��E���)�kv�ߧ�y�2Jo�0���E��)c�3���{og�rC#�+��T�(��}'�hQ�����}��I�T�Mf�o�v��(��oQ�L~�K��Y�
�7�ʃ��x�� �%i�!YU�������\��5ǫ�(]Bh�0����A���.�+Q�4���'��1>�t��j6��,�*�{1vLZ4����J��5�'c���f�����x���Z
@f��C�FWyż�֜�\G��{��v5�3'[Nb�6�Yn�NV�'M[df�J����a�ՕJj�2c�I�������`~K�V��it��i[��o�.A	����k�Q?g���L�s�&XvR�jo����o��+��������s�T�@�HR���sNZ�c���ks�L}�}�<��ąi�-P_�QQ���*-)���E��-�����ds���sA��+���7�^�����<@��s);��s��?<���GSZ�Ȁ��������������-��/&����x�G�9u +IA7A?q?Y\��5l���f�����[������)a6�pL�^G��55<�9��r��]_ڧ���d�[�o����f��U��3Zw���{�@}��"@�>��NS3���.�^�6�����`�3���4߅)�
�1�R�}���Q�D�)��U� �\f�c|A*- !4�ӫ��_���'9eq�VH���+��qɧ��h�9�]���ƕ+�u�B�s+���#��!�؄���Ã\��aȶCo��N:'�%ٳ�=>�5c#�=��*ϦΑq3t�o��f��]+Q������/p��ͧ��![�o��(�o�j��?ߐ�� �r;�2?i,���a�}���>�X׍4I�~���f��)�}PӞ�'<X�2 ^E�橀j���#�x[�P��~�u<�ÿ���Xx��	�g�
'AP�ng����RB�j���ŋ�ε�ME�Q���_�"��;������S-�,L�,�?'B�xz"=|H���#��
)U��>׫��7����T�2��J�8 Dl�\XR��LT�Ӵ� �/ao�n$�B8���I7t��yI�<�>�Z�/����c6	jO3��2��=G���?XX�����	�����^w4�^�azΟ��vk��|�uݼuu_=Vl�1k�U)-.�<I+��󏗍��J��n3h������"H���^W���+f�5�L�-���<̝��g4����)`���̰<�_�4��W����dcĥo�C{z�$x���I�Ɨ?vq�M*��8L�@�~c�J�� b�_DEs���r�y������:��냻�k���vpw�����%���;ww'8�����o�g.�bfu��]�j��.R���t�����=,}�-,�C���=:�$@�[��s�����y@|^B�ͻSzɣ~Φ��J#�N
Y1�$�gI�؀���2θvD�7w_�K�Z�+�@Ҵɳ�1l��Zm���w���a�L��Z���-�a(��B߂怄�D�!�R-D����(3mD��-��:?7��6����
�,�����<����X��NP����%C��h>7�'�_��w|䖜J
��
f.K!�_�^�>Tr1ѧ��~m*��ig}�� V~��>��a�o��a!Ϊb���-�I�=D�@����O�L '��a"v���|�Bi��y�tno(
?[�U]#�;�2�p����#�]�].@�7\�;0�:��:��2c��A�V��.�|!�����8ā��ǺC�D�P�ϳ��*t$K�Ow����Q�^}�h�5f��Q�u�Ơ/�Y�3�'X �ƱnE+</�^*i�m�7��4C��[h��=��QOZ�)?k;_�F�������)R���9_��6��z{v��+�UL� K��u\Ure;t�@N'�Z��~8r�4��8�q0%%ƻ�Ic�>���Fz$,c���*��ʓ����}Y��?S��]�u~���K�Ƨ2Z.t��ᅪ�,{`�&����k���J�����-����[豀�RP�`w�jTR��!aL1�li���֯:Mu\pK�)-��޼�,�Ʌᥨ���m�=7=-�a���g4�A{���S�yn?�+ۍ�iU��3	�AW�u�� Ǹ�u̿�{������Bt�iJ�P�w�4U�pce�̥f�YT)%�`�(��v�$m+h������܇�^py��*=�+k���%�4���_e��,�ƹ�Yu���2]߂q��qF֎]O,��S�`�wo�
ݩ�~��a�� �����͗)N���H�g!g�7w��Z�-j�hRv���h��D���hif�lO^M��3����+���o�-:������\K��a�E��Q����Ϧj�M+�ޙ|��eR� -W�^z���+8�,�^�}��\�̠1�$6n�կ�	Z�28=��NrSV�o ��;}K$��N���mRC	���Ǫ�g�7���_�z::��M�U�,l�ڵA�Ğ�n`+�B=�~
�"��2M-}N�˭T[�DmN��>`�e9�7aH:����W�|��T0�đ�ӥ�2e����i��p�ep9d1u?�f;Г���u�%�Ww46��J�W���'�Ɩ�!�L~w覹&��Hڭ�+��4Pe�Ozj��sC&u
�S�.���E�2��>l��~�$ `D���t�<�O"�}� �5�?�����{s�9����nht��ӑ�V����\[	a��(��t�[������d�qg���`�tKZ�'��C��eee�q1����h� �&)8PR��[�Ϸ8OW��=�oK�n���OR�(�l���-i��v��@���w���1����$�� �rN@^5.�>"Mҟ�5v� @ϗV�N�����0����e�E�����;N��U/�JV�����i���;*_	��8D鲈=S����,v���^�}.cl^[�d,C�!o��ld�^�A�U侵���m����u�$s�y���T�}���^�ڂo�$Cra+�7�L�yߨw���o��R:�z?U�D�W�wP����K|��$u��h���z�[��=��~�� ¬�O�Ԙ-����l6����+'�����\�H"��Y0 ���(��&�a�ۮ�6���SW�n9f- �w�A*��wb�&�F��#��.��XLV���i��9�W�o�%���Bv,��[��-aGG���@m@c�5���A���%}��x�ǃ�!�� myٿ_9��P{0����l��8 0�>���{〈F�?�V��і�vC�2���/��^�&��RJ=��[Z`ߚ!i��V��8{�J$�4'�v�߃#��2s��[���E3y��G��-ZtJW���+
��	�`��6��Mٔ2��\���P�J&ͅL����$t�-�c�n���H��;*݄���DHD41�,Z9$B!̘�y4�@d�HƌF�.�o�nC�,���a��펛"0͋L"�����f��磬6��n�]J� ;y�>�b���dF�H�H��z�R�mD�/��>*�\���'��IL�j����<�1�ާ��3<��4)(�m�)ȓKB�=[Y�򽱛�6�[:ob�[��S:�߿�Z���wx�O�Q<�{ظ6�����2K���#GUu�a�����-��~��|�T5�Ǉc�Sx�s��c�Og�$K���ލn&7X7mY�ꖘ�r'&C��AJ�}�����q`cf�p?�)��s�wc��\G�{��:�w�i����Jn�Q�BMW����X���}���'����7�ہ�Z��
�X��):Hn<�o�fm_Y'Ħز��K���TD����$����R�1{l�4�\��Yk;8g���m4�L?��G2f<��?�(�~^c]n�u��PrM�B�>&{��-���D��!"� Q�qΡ�!Aa�4)�Yr �?s���cy�
�H�`?Rt��wn]���'Yk�U�;9�f�8nb�߅�\���H�.�}���\�����HCD��/HrS�}��G��Ck{b!�=o�M1!!O�*9�_$
ϸ���v4�{���2\5����#>��v��}P"�S���b����`Q���1�tА���?������ķ�!@u"��Z�%�_�$wh�d�=sH���sࠚU���	b����i�3�����6�0P��j˶�M����ّ���;5A� \���=�5����_gG]�[\L�y\��@�~�!Z���/�������S�o�xAQ}���JG��V.N�H'��~y����������9\�n�PR�_"^�X��S��]�kT��T2���n�<dSi̠�jç߳{V�����6����F �œ�R�3�ڞ�;��2-1�:V�d���'5���'v˦�'~uX�
���n0��f�{��*a�?f�E�Us	�L���Բ���}�SQ�z��������SVÊZ�z�uim��1�Pp�;�����Z��L�Ou��E�W��|�L�2&-��R�*����EW	��(౑�<Mmƕ�,�F�iU j�2��n]H�&� ru�ٶ�C����F4z�����`H��\g�.�z��Q��L�ǅ��p����� *!�u����4���Q��$'L$ťCC�yQ�~�D���<�<�(n�mBW�{����~���R�1�΄ @m�~7��cgM�B�1�_�F=����S%>�Ov⃫]��q���6���K���}�Y;o䬋&&���{�f���=����}�Lܡ��*ZLs#:�P(~h-S̻����f�ۜ�X+uX��f�nط@t=}�Zg��E�'�s	Z,�����b��� �aS��t^�͘��s��s�6���&�ކZ�m�`�V����ށ���\��$1��C����n"��-=�%�0�snI{D$��Tha(�RE2P�亜Xl��X�8v����\7��QI��My�s?����W�p��N(�M��n��V�ɜJ�j����A���z���|Z�T|5�p:߹Bz+z��J�݃Qգ������k��Z���q�.F�r����G�o�YJbf�Χ&��96���AB��|�!Fӌ���1��z>P����<LOB{����W�ed�\m����c��f �J������M�#�F�YL�a��p+��t�M2�� y�0E̘-w)�'�yNN�.ӷ��憢q AO��Ͻ��}f����)��c��� �.I@'���k�ۍרtX���J}XO��L.�*��oNeP�5��]}���ܗY��	re�%����(`KgBQ�ɮm��9������ͻZ���{L""$�,R�����rm�co3� ���T�����c,{���z90�4���3
� � <"^��z� U��ZdC����)��v���ki�5�(@i?\R���?<�8�i�-�}�:�HG)C�Ad���^2������D޴�P�5�K:���? �u��N�Y�5q�E�{6�\�7<31�G��4�����w��-�(YQ�a���-5��1���I5%g����[pfn�d�X���4 *�U���7�i	�"k��ӢϮ��!K�z�J�6C�+{�R�:D3��z�P�j�׋��׫���}��4fXǗ��	�<?����#�t**�~B��;��P���!+��8F$�}r��6�� ��|��|��N�{}���4��b���}"���M�Y/���͋�
�	V?I&�k".g	�.�lh��g��S���8K��{��N�Y�ЏV.���ip���!5��m�|�a��l�'�TQ���U��t��+��K�u�[����ϩ�̍=��j$礆e4af4 K��X���n����M��a٬��������ǉ+&��:ds{�iKIN���%�ɣ��������|��hw6���ƈ�F�\{G�V=BS�B�Iɢ�c��4w+ sk�	�B�f�`I�0dW��ڝ�_�
�w�,�u`�>+Mp�*�3X� C�0��'�Q�&��}fbo@�œa��ɵW�\�]��̀!��Ze,jD�d�=���=N}ޣ(��Ye��ذ�Tǻ��/B�9��_���Q���SM�Fp�P� [O��\�I�׏�
��^a8x>uqj��qҫī��{4�%�MT(JdO������ï�ue�,�Y�$ދ�y��*���b�z���}���_��Z<�Z��KpB���呕�q�#˽�E&�:k��6��Z����.՛ݳY�\��~Ć7���襕�_�4HW��u���$؃:l�!�,L��F*�$l�+��PQ�ֶ���,��`��@� o�u�QΎ����L��:�
�\�uF �M*S̮R1��_S��j
���\�͂"�Юm�\�ة�L�)I/9^�B=v=��R�+��<'��E{��f}�=����N(�&u$F��.w�4�=WE���X�$��W^�õ�@FR�k~V���{ީ3�1ݑ�8]�'O7��2D��t��$K��$Á\Jh�劼�nc}�Z�5��Y`
7����t��֣h �� ko�ި墴�Qm���h)�=K���9�C�R�P��{�	�f=�ޅi۠j,���n5�7��2�m��/���'���F⵬���|H��~��Bl�+-�(r,g��]�Bo�U	��׸��,��/k�<�����Ehԣ�,J�+��}X��t!���~<����Lm���_�=D�t�)ʜ�j˥�`r��Gq^�'�ZEFe�x�#��t�b'�f���Rge�_ٕ�j�^����!2��v&Qe�*���F'�>!?N���,cs��üb�&�$���{����u��E��[k���,�|)k��dק�YR��K�1\�[��a�����@���=��c�2�^=�K�,�a$\�����"  ������Ƃ�b�;&˴�k��mg6�W�`OP�q�X8 ��z���?�?��!x3�"��(\������j�,P9�.����\r���2�#���ʸOm��|j�E<�����j	���Y]�2���kA�K�0&�ԩS��Ȯ���:V������� L#'��LV��&�Ó�U 2f��XY,W�ե��c��s�` �b+�ۻbo��sUL����#.�z(�<�����cjyYL���N���SC�1a�( ^�U�=���C/k����3��s�^I�<����r�C�v���zӕ�PјƘ���]���)��9U��m�L^]�,��&l�(,��6�Ls�<#1W���P}���S�s0��1g�Z�,���������-�ЊM�X��Ge�+�v���S�:�g�]M8������O�p�3Z�>Yg�?L9�*��Lx�v�9�I�)���u��6Nד����ʚ���D �X�s���!���W�z�lx��1�^�*�*
����$U���J�����HI�Ec�[/4�J���V����=M�z�g	We�_�?���V��Ff����^���ǝ�����1��ퟳP���'��yi������4�Ϡ0��2�����N�EN`V[y�A������䬉yq6��-X�Jq$��Ho��~ �W��Դ��>��b��E�tT�&�Pl�-��6�;b�sa���լYc�~H�Ԉ�I���.���M�q�0#�{0)�$���(Fl���g�w-3�������f��m��4���8?H��oNRL��{$��|�:���]�:lG��xx�x�^��:Gc�	ļ�m��L�l�=H�b?�/ds�����i9�t��������ݓ�X�꺆�b���@�xw�[��}�j
T�c�G��˰�:�ѳ.Rw����;�I�E��8��������`��
��������5��Y���&qpC�#s%A6*Xa�ú.~�(�^��B3{⹫�W�`	o{8s�HZ�2A��L-0'L���qrF��y� x<;�lQ�A"|�[�y��'�}�cr;̠Ð���~�̷|�o.{k�^-^(@F������G�J�R�2\�fEd���cd�Y��oE��]J�1X<Q�.�΁��H�`:�6�:R�w�8�OCt;=g�}����<;����vT��!R2�0���Y�(y���ٵ�Ju�}�R^(��-z"2
���\��4�U��9���ڌz8�`2�jϡɹ8�v�����_HY MB�~A�X��������px��`��\�!8'(�ɔf��A`���}��N�_S�'�P��xt]ǒC��ۛ䏰؛��Y�~�K�	4E�cux\�("b��p]ߌ3��CA!�&���'��;G��A���2���YE������_7�U}��R��˹�l���W�x��N��$@i�i�Zw�Z�!���� [�H���;l��r޺R����C�g�<�v	�!��o�[g���� Nh�����l>����%���e}�|d����K���T��B��y�^�%��f����v�����@�}Eմ�cFb8�IH\�Euw���2+��L�-�7�Vڳ��ZT�`χP�$�6�.U��6����վYw>��t��Q9B�~*�OSO/�,��p
�"A��*�Q�5��u6�$��APNq6�2*p��ל$O�9��s��_X��17T���G�� -x��J�_Z��wVR��B��8@܄N�<%
.!���6w�> �%�7"Z5N ��MyCz+Ug|��*�/�$�R�oqE¢#�v��Q�����R�������x��/��8]��G\�Ġ�p,�M�����?DU�zxϯtC�QС�]q��zz7�g\��Q�YO�T<�T/vc��h��g@�d�K��9y��(0n�_FF���6��O��Q�B$��)�<L4�%ϲ$%�B��F	����D<
���P�8s��:�Us���W"����QW�,��@���]n-�:�xy��~9������[��H-��������'����kp*#��r������m��uw�0������xE��T��u���ޅ+E�#�Wk��O)wu�5{Gb��:7�V���:�No��j�+n`c�)sH�#��.'T��D.%K��k����Қ�����b�s��O"ݏ �
h����2�Š�7^Qf�t�x_z���_i��AgR�8�3�:V���#í�Zq�u8���`Q�p1���lPA��+��x< H��J���/���[`Pz��*;�G�=�Y�B��Ԣ�/#Hq=�I�N��y�B�z�V�ы��j������qM�i��qe��2)�`C(�|5'5�x��o��NNW/�<g�-r,��i+aD���/>{H�^d$(�S�b��ͰF��N�v����TT�?o�C OL;�Y�J�^%�`�Sj���/�yUX��ѩ�����z����<�Џ�H����Ӻ*(���A��& k�A����*��)Ƕ�;t�$�D�����Y⛮@��]cDǢ(��T1V��3�������a|��9���WSK�7�9�lE�)3��`�=��~���d��͵��)_�lQ S���(%3���QR�/B:�lD=js�2��b/�6y�̬������y�LO�R^���+�yB���J�ԀSʃ嚢�����c�yxB�p�cF�1�Tm6�,֪Ɏ*�^�އ�JN*_��~Remo���ȀoSߪ�W���7�R�����i����گ0#C���2�剙E6��w�r^5�i��Z΄*��޶)?Z~�V|����R�
"�7~M\!��	ƵJ�%V1���/l^�kp�g�iԌ%6�"��1���)ֲ��~i��;�􌪮�,6��'&�°�5����7	�,:I�[*t��@�"����ԒRf�/��c����hI=��>��lHґ�$ͼ�ω�+��@��;�H�H�J	\��T�;�	7�_�m�	8���Z~c�	��m{`	snR`]>K{"^b\�a]�"i�ὥEr�w�M�'ʲ:��*u��=Q��!����D�4^���%UU�O��OEbJ�[�9��7�ꤝK�\�',VC�ߚ^�z���t�wT�߼|�zB��n��w��ʏ�����.��:ҝ*m/$�h[M =�豟�Ҕ�:K�|ݕ��L�,�پ���V�8|`x l� ���na��z��JB�E��0��!Kc8�B�X��b�4h/����@Q�}4�CᎲ�.FtE���kR��X���'�R��Ȧ�����X�cH1ё��q���!���
�KL=Y^�^d�/��K�e���dj��{�=���ﰝ�^��1���ucҬ�c∥�q�Q �Tl���C����2��y#(��0/���9�|�+�w�|��Y�aM ���JU?Yy�e��҈X1��H�ؕ�R�%��
�xѝ73��n�t��t��Fx�iK�7�	��dp(!Ӑ��-yЧՑy͑RDe��.���@<gA�R�.)�e{fLִ�ڒ�����a �bJdn�4D��?ԧ �_Qh��*iL ʠw�bTc��� #�`���U(c0L���&�۬��:ۧP�jF������Xy�d�TC�����/��wQ��g;�˭$�䏧qR!UWa��~H��?/��j=ZK��Q�*��jc}��J��p/��0,V�O��=��0Hэ]�!%�xr��� J;�x*�A&����vO�A��� ��$di�S���i�����
W��=fq��e��: ��tO\R�ޛ>]������c�SC�4�a�җT��x��C�|��j�MG�Ę��v�Tz��@{9�����IێET@��}�ə��v����Sdq���c�����*�~�bD����^Г$7��W*�$�)��-�Y� ov�����TfV��'�b��'V�|!��g��0���$�V*v�\�Q�@��f��'d����̇��悏�B�}��-�1�<瞘�l�J��S^�\��H�)��g���ـ���R;p�@�^������V�"G!G��3���0fN�\������]�/:�Nx�b\v�1Z�s�߆�a�t�V��(��<�~�P9���SiI#b|��ſ�i�ܠS�q��9�Ez�)�<9ِu$�(�h���_����KCx�w��/pX� ڛô2k;G�[0��a�NS'HXJ ���Z+D�0��F����͔����T	70��Y����}s/3�N�U�Yż㊰db��o�`��⫹��]��g^��+e�[t�:���8���):Q�ۂY���˃�E��2����ϫ�ttRY�������`m�"qY�2ͥ�� Oy����y��8����P8MR!>1�ޱ����Z�snb����[Y��@]�q
��wPfo_Y�#XL8���b���x0*tS��T7��2v*;�jz�o�tae�Oh�6'R[V:�ў��̝Q�4�P.5��<����fzTH�5�bЪ��5P� I�oO]^κ��}H]�	���$p���ꫡ�Z�$�r��Ŝ�_5�(-wf�P�� �/ÓEڣ0T_�`}��;�������t�b��|\�mS�Ż�<�y��/.�@���Y�l�Y fq�\B�1��_NI���(�i{ȴ�y���1���OB���[���]к��)�2�9B���zc���@+��%�y�eEI;{�@��孳Y���#\�nhu,�������rt���D���mp#�/��HS8S�{d�ށtiN�����&�}�ME��A���!>�z�Za�՛��-�e��TʏD�����R�9\�R99��>�.����
��RG8��R���T�HK�Z�d(.i�`�!z~da��3�����z��)��Y�E�IN�^g��3/�MK�H�����Hd�H�Jah�g7PM/�5�[�ң�����W�{ؑ
�������&�+25}!F�j��Φ���X�6��ĺ�/%�:5���nj��3lF
d������R��Fk�41Ǡ�Rs����ޓ(�*�����)H�#��_�8��eK^w�����ܤ'�aA��^��/�T%j�n��SA�ڞd�;Ti���`Č��Ej}q�7��b�U+�i��N�Z�M�m~�@��2�*�8��eJ�!'/�����&$���O�N�}�<��m�����	hv�LD����Ib�f�Ní)sQ�Qr�����So�5B>��l~/11���&C��=xh͎P���_���
t��Nj��õ��w.}�g&j�����H������#hZ�� D���lQ�r�T�4�0̀�sJ�A5U��8�m�#!v��& �1>�R#3�<� $�Y�!�71���@%$XW��׸��(�TƯ+���?�P� �1`lΌ|�D��A�B�`{���]��x�x�{��� ��@������ ��t#�����e�F=������J,U���m���h�-���A�߁���h��*����hB��jo��.=��G� �g��^��"CTҰ�l��T'@��ƷAt3�=�����N+����6����f��7:��d�#���_7�Ih���!�*�[��L_�}��_���g�_o$�q���6����P����?����;�"&qFV������d@�~d��[�T7?��3��t>qDA<��QW�C�_C�#G�w5��,�h�u�n����t���q�D�80W�|��k�&9�?;�@�B�x/(1uk��P�\�����B�p\&�CPP7��p1��D��n��o��a6������B=Y��>(z�^�$��&ô S0[L�nF���$��'ܡ%�^��M!�&�6<@�^o2�+5�'������	�?�
��L�{���Y��%�����������@o|y��9���t{����EU���p	�*�g����"E��1	b9�PtD�/
��j��_���3�U�x�C�4��Ǐ[��F��4�S*o��_�6K��
�����m�W�0�	��W�1�PK   (YEX'�T~|  r}  /   images/8c7873d6-161f-426c-8be5-8f6703290c9a.pngl{eTM.β�;,��k�eq] �� �]�Y��$��w��4'H����{�;���T�LOwuU=]3]Q��
�@
 ��"T뵌F@@| ���ơ{-ݵ 5STG�����B}<�9�+��h���@��ߎ���x��4�����v�uQ��0�4�0G�o�p�u�t�u�p�3������y=p������҂<������h���{��L%�����I�^�B���!v5*"�b�!�f>U}��^�#������{��Qj��ͪą���K���������?e�YN���m�a�~��KL��	�����r��R���%|XJ\���A�M���X���k�r��b�e	C�J�f��U�z�ڏ�)�L���\�ģ��E�6���HS�&$1r�	(�� ����CrVA0�B�G���m��|ZT�""�g0G�V>L��)Օ�L.Ůޥ~��;q��C*R'ksu�+�=�G�^3�ꔭl-m��7cE���E3<"b\ok�'�j<M��� ����_0JK�YșI��p񽕓�jjڤ��d��pڞ-$�lQ����Fl�(uz�m����
4Vϕt\���j1r��x�?���C�wR�K��-V5���v����~����~Z㤄d{��K�J�LFM�����&�6�g"S��K5!w���PVS@�l���H�l��z��]�F����ő�{���J�,������*y�ʝ�S(�I�o|A�[�cPќ���� Xk�E��,���qB�#�؊�e�e,�Ε�>����]�>:[��7�� ���OǠD&Ɉe��i3[�K�2�#)���t01�/ߞ;�{��`��77��:d�Ie�L�f#���M��MMc��O��-�B6f3:Uwn��߮�8�F �]�C���-��G�U�p��n�>��R��	�a�?���vp�)1�H1�K�[��y��&\e�ID�}k��(��T\�Οş��y�D�`��κw�A���L}�'2����4��D�����e_��`�����?]F8����9���Hxiߤu�s�/!M��,ނ�+�V���o&E�B+R����XOBcBH�ym�
�*����:�N_�k��g���?�3��~���9��q%�D���4y��;�N�r�����'�N窋K#nø�����6=*�E¥ /�LE��4��i:��Ҡͭ��k���~/}�$��8��n1Y��rJ'���G���ٴT	��ş�;[^>�����/V�r�f+�S�7��w�s�A�y(��׏N!`;nT�|��e���,��0�y�v��0Εܹ��{:Ww�Gz�����!�+5��c/���hS�ӺX����h����������^�҆�vj@}b��oK6�2�Z�)��iVX8�n����Do́3QK���ӗ�����K���O�g=�)&Q'Q������ö���&B��w�I>��2 e"�0b�n��*\��r�O@(fU]הbhCQ:����.2��Gi��zy0�ҋ��"g� ��5�A��bFU�����\��&%�ן�<��ؔo
y��?P�r�.�%^����tj�y>={V?�8�d��k7BZ��#��w.���@#g�FNN�N�Ȱ�4�4՟�o�}���G}���2i�\iwXhô1��V菗k����F�ވ���*kA�R�	��]����#��Lac�Qn�{2,��8Jt����B܅��u���Uw�K���Ո�8��O�W'�o@��p�rk���Yx� ,ฺ�r�ٱ��@�cp �uq/y���������ۗ4��.��VV��D�4zF��{�X��K'�(�Z"�[�4�p�3�^���*8`m���S5�5y��Q��p΄J��o�X=r��}-��+�O�����m�'�7��x�X�oִtBBd@Ks�Rw[��vu̹7�B��47�.���U�&ƾ�x$��tqØ�t�a�;��0�ӳ�DAiF�+��ju��>�.�����%���DOOb�X������b@ۣ�R��<'��v���"|i2�����.����s{i}�.���&�K�+[3~G]��G�7!�/���I�6���b�v�,��V�{J���s�?zU"��D%Ny�bx*�ͳ��V�(*�_�<b�dT���bF檍����8]60�!HDAY�����������eS?5��]��#�� |n�/au�LJg/I2�_��������ȎB�N9�J\���8���a��|l
��X�v�Ns�'�w�&\��qq읭�d~K��uȻ��S��-��ң\��1�Y� ���)�GnNV�^}A�~�)����
�%T$f$M�CB(g�k��J�k5�p$�
�9]��F�.�Ā���YF 9���˽�ۻ�N**�YCY��7�����w����*�
朊�G�p�*��h���Xq�:�Ь,��`��y�ƻQ,9	馾���T[�(�AN�##J���� ��q���TjI�rw<��tNU�.��  �b���o��a��Z�xZd��$�6�9��h��|����5Q���R�Juy��X�D�������Z|����쵙H�:)���A��X��L>��V�5&�#�}<�FE�l�>Fza�i���;�*s�~i�⎥(Rغh8 Ŏua��A�w��Ջ>��,?M�-c!�f�\� �����iU6E
��/�B��d%V�5���5����/��uxR^s_�[۴����j�yW���HM����U'�2F: �Ϲ5ԂRȁ�/��+a�}[�C��~�e��c_�e`��/��W�=�8�En�<��{��&��: �*��^�f������T�:��,c��G'����r��is<�������,��z�7�B}�Ȕ]���A�9i��	4��!i�QX�}%# LhK��s�'�������$fq���>�	ڗ;�W`s<�.x�����+�X��w�%==>��k���J�<J��co�H21SV!��0`lp	�L�}�
�z�aƖK%A���7��[m��b���,����@�Q�(��� Nt����}8����,�z�{�/L�l�r?��S"���l:5��H��6���dۥu2�4��P~y�We�Z8B/��f��y�U���^�CXO�w�)��.~�/W��-���{(k֟Gb}B/���1�b��5:�`Hɖ���Qi��0�'�i��h7J�$0& �]"3�)�C@J�`��a|\�x��g: :7�r{L��cM9'w���\���9[k�w������V���IK�e���o#N'��ߗ���4�Q�������g��Qӄ{׉R/!A�㲜�Gsf�g����"I�n�̳ՕYл� d,@�Xw!��K���6�vC�Z��l�d�*���@�P� �uO�7�<�l�c'
�z���! {��C4��A�X��D��@��{�x�mI��eS{#y�zF�c�<�.�.&�wg �mTrdߒ��H���A.B˒ɝ=7"�Kr"_����DZt'���i(��kyT��S~� ���-K�1����'�(�w����O�]t�vh3H�&ǯ�� �!��:�W�g�;��~W̇n�A��|1�_94�cB���h!�p�뇿>��j,�HA[0,:~�I X��+���f�r��l��
m�X�'�##B��RwT|�����C}��P����:R3�@DLM�
D���s�Ē�n>䣟�\��w~��M �ω���I��
���'8�����c~ϊ�38�h��J�mP�ǝ���B��>�ʋ���W@f)�%	�3�+uH�Pq�Z����F�c1F�����~�*jq�$�}�r��!Nx�pa ����k����cW��F�5��Bre�2���_�bnlL��S�|�*vR9m����NIF$=%�+[��bLI��N��0�{��1&��\��'�㼣�)���w��c��'�����Qѕڻ즚�|�h�]{h+5F�W[�w�b�.p�_E����]�,�¡�,^y��|�,~����|�F�p���8�ID��k$"���eRQ��B��ʹ��EO��g�ˎ�zl�̂r����O�~�9��E=��WQ����$�`��i�޸�s�d�g� r*�WlE�>&eeL�b�PEv,����k�ϳ��Ĩ"#ݔ�7+����%ҟ�iWF8P���{�N�R��O����$P�l����YՔ6ܓ8E�Qq�H�J�y�๵��a�����tY�9iC�}�������0�3��RF�@��2�QM���F��I�u�I��*#B���`�k�Ikrx#��T��4G�j�O����
Ac(��P�����ϼ���ԛ)/�Y��Ȱ4p�g4�q����jT/������U9��.$i�
�d`F#E�Zi�x�^(xǅj@���Ĕ ��}��yh�����2iQ��Ά�Y��d̓C��o���:���*���4ղ��t�"Iu�	$�##DX��f�|��.���~��	������	�2�UE��x�#��vӏ[�1n��\��Ѩ���Q��Ul3l��v�e|�A�eq�H}
�����_��G�Dt���񌑆��w��H�W{@��n�;.����*��%9��N�Y�"	OO1m%rbfffS۞-,ޣ|��Y����M�"q"�(vkI�(�&��|�4I�?���ت�\7?CC�߭+rz]�c���MKDM�k���ߘGW:�=��6u��{`nM8gY�L��Q���R�|u.�l �n�1�!ߓ0F}��`ⶽ4��6sc&,�m!��uTh�}���|�B�$�c\h�\�O5�\�T( If�SBE��/��r̲�ɢ|Qe�?�,pHwQ�}���,$gan���������j��9����sH%�%�a ��{��)o�[Q�UQ�9U��n��OŁ�'�B������S$E�0S���� 傒��GY���^bUDMB��R��xq4D.�H@86u�u�Z�@U$��h�gp�7NK��<���t��4w��˜��w,�`�k�FQ��:��]�P�3W�]�P]�}�U��%�1Q��zz��C�̢���<�;�ŽL2/�r������ޯ*�L/�жUCf��8?�CHм[[V:4�qy#���c/����_�~�h��R��[)�P��v��M�/7������K���M�ҍ�VE�`F�/	E�=���u�[����Ax�"S�5f�W08'$�Τ<֟� �v�{�{��0,*e ���}��q�B���\=����6��B߶f��Z�
H�9�ā�D���eT��$io���L�����y[�ֲ@Am�w�T�E���^�C��!-��@OD�
����c1��5@�&��>B�&��k�:��/� ?<`��Ę�U�n�=�ʬ�OI� Mi��`⋨�8\�܂�Y�P�x.(� �i��Fi$�6���a�WJj���~y0
7 ���C���;�
g��{�B�2�#	<
�
��ssFPG9��g.���|���nW�\��blEߌ�6����y�6x�|�D��}L���?B�o�y�j�q�c2qX�٣ҍ8e�$\V+eq x����,`�3���G!T�^ �%^ ax���Dz���������M��|����.k���Bk��F��C�k���T��I���I�=�'�J���/K�e�v�,xa�zݗ��G��f~h�m���(���W(�!cʈ B����rͦy3��!����r�w��0󳡍�/G�9�
�����LΟ_�����ǟ_7��b�1(�#7���5��)��붨�NFL��)���O��($B�U��X�o;1ZuD�X[ǘcd��s|��H����= P-C�s�Q�(���\*������/Y/���wl�9C�eWj_�lkU.�na���AX9"\+�K��M�;	�0�G�����
����<���KF�Mm�"3�aM�����G_���z!�x��l~��A3�$�����c9ml�\~]Ƒ�<ZL2�X�!���>Kۆ�c�vX~[(�TKO���f���)�����Ӎ�h/ZH�TI�w��r���bL�3�}����*�sx4����H��n'龥戧@<l+�}>Z��ȳ86���>����7�ǋ�A��a�<	�Iu�2	�SLz�&_6�+��N
H^�(P%�4A���u�啼̏a,�൘�~V��������3�"Dd�-<��)S'�ߣmO9I��[���K;��X���b#�4]�T��Vn��(�󣖵OØ�KbBUrÇ1�kh
��;��M��uQ{��Ͻ٢ �hU�Ǜ�?��#���#C4�W����O;c��
z[iKx^�.l�gcg�m���1�}�0�I^��Vb����(�!�w��i&$�%�n�!�|������g�[+�kr�������򉻨N�J�=��+}zq�xӊ�-�4j�$,*�L���c�P*h�TV%Xd9յ>�A��0Q� ��dR-=���|u�!�a�I�[qOBP��I�r(���
6��.�"V�>����u1�~:�soS�g�*�j�!������ۻ����$�ʀ��N&�.�2A�
>�������2���`t�m������ZtBZ�O;�X1��F��!5�`$�Oo�F��^�+e��`�7��^�d��"}�݀��Lrban }��S�����YDԳ¬�IH�����w�l&�� Ş�l&S`n����,a$�=hg/9��!ɛ��P[�w	��܄qD�p1�����<�@fJ5y�-���i)���6���"���7�����
��I~�b��$F}�
.hA-�/'q�o�_���5y6��!��#����������z�������]_M�4���Ꮎ��S����w�n�cvôkbv��6��M�Z#Ƭe��e�4�tδ��$c?���*��������UXHp �F6���A�(M@�}����P��rA	�os���Df��J@��_�a$�ŵ��u>��GٖL��������o)��#�W��Y�ᑸ�
p�s�{:��`���xSY䖄��TkVү��������}>w]qz�^zz���#D�Orimf���.��Cȹ ������$������:
������(!X�9l�o�Z��ˊ�:K��+z7�	�uA�H"��&%����祒?�6�(�/,�)�B�!"5X�LU�+[�����J��4#�tT���8��K���f�X]����j�([+!�.��@�[��2��D��n�@5�PG���_P�%}=vMO3q�eS�N�S�8���k������Q����f�y~iN�iE1;������!$3	�ˡ��%R� �&Q�&�zDK@�Ai���n�X��Y��f݋�qwW|J,��F5O��RȲ,QZ=m�6U��Vq1�[�d3��V.��<+W7�=;�{>�l�Z#��ɻf�Ώ�"�F�ۢӼ4T4*!.�WT�rE1��Z��;�o�����T�>J_<0IyH��0�ԛ�52�$���BU��`	�-	F*���$EZ�sa&"#��[5O�R�PS���J���)���[�s�"K�T��R�U(d�]���P��g��TG����t������Y�Ӯ%[�I���45���\�
�c��`{SO2�������:v���'���/�/m���;v���%��-�RMp�hĦ��~6��ر��BS,�æ֑R`	C'K��~�+׊P~�~���Mʡ���a����XB����<��*��TԘ�*�T����J�7M>��u���L뮆ӹoHc��~ᅕ�3f�|��`-��;�b��H�a;v7�&Dd��Fr�Q�T��8k~}D��9��0r���=�qg�u���8j]�jV�,���/����'@)��/��*j ]���	��v��)�9�a��w�3'�(s�e�2���Ë�>���YN�u>s)�O�D_���5�/�FU'�ǰ�9������\���]u���'L+�V˚R��KV�t����x������7�[�翶A�L��U�HѪq�JN1�,H.�;Ǖw�\�Z�����Y��{�P�� �0�+�B�o.�����0��0����G��(�V��&V�~Ɣ�0�=�a#��1f�*�����c�|�@:�����}�h��T�*�-.5�!i��-Ϥ��%��aʩ$�9ol��/�$N��e�p�C�⠫�b�Ѝh꥞b�N�{��݌�zY�O~ќ�Ͷg�N�O!�4U�[�dè�T��#�bK�q&a>y1�J�]���&�K�U����~�Nf1.�CH4�ra�f.��^��\ҶPP$�M&���Ab���XE5�a�:��b:%v��TX��Lw�\�3^훔>dY��s6���L+s�g��WT�T6TSd�T~���C�%ꛠ�³�O�M�*�m*�Oܪ㝏�r4tG���l��"�������&���yy�ͭ��7*/G�>�շ{-=ϲ��_V+�n}��đ��d�<�U~bV��������U���m�q�#,j��I�|E�z���.�i[J�ג��)�bߴ��ř�p�O�xg�\��2�W��4{����.�g����k%hHn�D����ET? �@JP��0��u��b���LJ|]4{���̽9H�@>�x���#wݥ��c��"6����*��+˦'&֏��^�ƠEǿ�Iw{�a�!?tr��.���m�JG}d*3r�C!�IC��؄�$�Z0&d���
�}y<hA���)ʧ������?������Pd�hՕcro��&b�h|ߴ��5?%��+����ZV7�%��Pz�"��,��!c����Q��Y���,az��&�F���D�uz[�R��m���F�j�+�-���OڙL��Fj�ų:�x��2j߄~*���U9���T���e��ҌH'?2����I�P��2���=��ny�2m�"L;�C�Z�s��2���Ҵ�}�`n�[X��T�9n�}�f����7��u��d(Q��P�\&he�P�����B˵�$>��Ӹ��v����-*�e�Bcs���z���Õ(���Z���>��jҠ�k_}��TZ�vN����g-��N��|6^&����0�}�P��&��p� �@�
��(=F�	e���;9��g�!�>|��\u�_�������T�Rd'�mS�ƹU3\	ѡ���WҲ�uFٽ��B�F�rdё�;�%��2 �@y���!�n�fG� `T�,�U �mCY�$@��W�2����:h�v����tl�40��8�8�b2S�����;��r��5\��4M������H-���ȁ �t/�k�:I��4�����/p0gt�i����WFQ�_��'��D�I	��ˢb$(��ݞd��~":Z��#@�*)���9+����X+s�&�`�q^Z\sZ���)�f-�mʐ;���fz �ggD^2K��܀��jF 4��������Q���Q�K��s߉�+xG���&�!ZJ��� ?`�#������(
�1tRr�����' 3�}ضx�����B���}'�́��9p��4�K2���y`=]`&)2o����C��W&9&^�g���U_ֽ��"H�?�rO3Hfa[���4�3#�J<Q���}Â���Z��?�<^78oJR�&\�B�q��4���ll��ϔ��&zCf="ԣn��";���4_6������,jҚ,�>F̹���B3W���᪲�迈��0���Ow���qFH����g�;����gn���O�7�lX4g"�Zx��o7��#������t�g����@ĉ�(��t�����7"\ϢҌ�^®���ph�m0d�n_�6q�^xG"^���8W���E���0u#K��9wY=ct��2���1J1 D#(��!oW�-":_���^�=���DbM41��64���V+͎Y�Zjɡr *���!�cM�������Ǒɷ�^�k��=O��\Ցit��?��<�<ּ�|WˀV���;8�[��z�����?�=R�`~j"���)���<�I�g���jq�Y�L�J@��م��U��U�F�<S�.�;�x"uk�s����ӕ4~�$��g�eD�5�qn���.7�}�|��L�Rw�_�8�)��i�bB�Uֆ�!K!�6�1bE�̤�r)�nwgp���4:e&6�䭹�(b��R�X1]=�������/�)l��%G��{W8�ς>֢nz���A�4�,�p �49�Ye�x\ҕ_�o�l��{
aq�K�(��K�X $�H=���@(E
m+#Q#�AN��ٹ�ݐ��K����9/��|́Qw�3�1��	��E� O�H_�o��>����ʎ�a�1;;B3��d}U�~#\�V:޾!T��r�9�6���'��XP4�.g�F^/%S�03�/�ſ:��f�ф�$L�X�]��f�{G ����߻�5듕pM�JmJN�Fq+x�B ��T�S0��3D0)(��sR��Spd��Ɲ�Z�ʎfuXʇ�
��!p��&Sg�;�;Ux�����g��G�i���Q�4���s�e3���'�N�v�[/���j�3��s�o��������u��I֣� �a�p��~:�[e<�3Y-Kh����v�S��"�ND����r��Q��ՉO-�4.k�����@0
bN�!�N3�?�Dx_cO(�*�kB�_�o\��J��DC��֪'�ٻVH��⊏Cy�b��Rſ_�jN��æ�L��ڿ/��JRː�G|�]��id�;^��J��>AwM��z{�1�� D���q�����-�-�#�A����+x7~3�yS�	u���ƨF���#(�����~%7���O��3�j���i<�#��ր��$�� j�B����˽��n�#�n�ZW��v�n�M�l������3�8�f^��m����[�{�����`��4�|H������3H��ꊯ:�Y�dv�ctta�m��ec�)��)t0o'�Y,Z΅|o!c�q]P�cx
�a�@3%"O|N�d�)G����	�y?�
����p#��Q�i�tW��� ؆j:�ZS�8;��܇�����P���塃iR��إ,�p��/@�P�)�1��0�\=�4�ml-/ 32s�Ÿ|"�����"H�
�	�a��o#BB�����OȆHv���G���~�n�D����#���/��m�~WZ���X������il��J,0K#���E��~%�N
o~[f���Z�a3�q�`D@sZ+�5~q��3 X�
���R�}�<)�Ll�D����:ڦ�����$�j̃�\d�ҕ�Z��@�9Ns#OJ�j��ؔU�];�쪺���QW�5�.顪��TøZ�Ϸ=��j�ɲ~jh�  C�qh"<�_�Q�м��H lLb%��G���NE��N\B�-.���B�g)�Dn�ZF�w�v�s�R��v��?˱N_|h ��6n.�谺�2�GB�l�F]�5XN�?�6����w��SPp�Q��;�/(#V��&�5�P�؀����k���y����|�#����Jƀ�G��䀝�s��{YWS�����i��,��7GE���i쵝s�O��.1
*����z����A�]7���)����+���(ɋ�;�z�w�1����D��l4~o��M����m%q�����zH࡛�O:`���^=�pf k0P��zX�;#��{PU����0K�Y���g�w>3L�҂�F����ٷz���$V���\�"�3�*n���~˵�w�ݗC��~:uR�厝�<P������15^Ȧ�x�B� "���1��^��Zt�!ٜ�/�r0��VoTMx�r���~9�[V�=� �Րi�������%4qJ�q��i~��A��D����E�b�t@����-G�1���^xsVG$��Թ��M��1��,��,VҨVǌ�c�?��S�j:NŎ�g)�q���
�m��Z�Mk���ju���7Q(Ix�;j8�P"[U�F�4O��V����l�;��t9�-DBa�m�>.X|���vV��dsD��d�*�/.I!�@w��/r��0�L|g7�x��bH¡2�O'W2�k�b���ܿ
bEp�}9�bM���^��0�!_�s��o�b�}X��3g�Ke������<���F+}����4�r��W�8�����+5C�T��ȭ1��U*�����9}�&�*��+՘���<{ p��{��.�ؙEfw%� ���puuK�����W�2sd�&�<ۅ�U�豚��=S�N��	N�24<4D5�Չe\�� ��$s3�"��"J�j�愈�	(�	d���_�讌rΕZ�%�-NE�!{K�M�ܺ�4�����k��J:��c1�	aʸ��`=&;T�g����ah>��.Cwʇ��H��P�$S�T�ç�n��zh����Ծ���͓0&��7�au��Hu{,S��	�f6F�Eb����
{x��#y��D��m�޵���@mU�L�"��pk��X���f��M�͒�x��2�����q��X�C��P>�w��0�&�M���ù��E��wp޷b�I�@ЯʸXӡ�ﲒ��+IL�^�1��_�F��3[�G��mWv2��5�Z�ϚgVNԖ�܈��E�B?�P N�䒲�-Wj{m� ᐽ���?�O�K�&s�X$�J:��ǀ�V ��'uo�Ѐ`�HP����/��EA�c�=T#��4&����^lȁ1JH�Ɔ�a������섩������o�6~)��k[������w���H�ķ�Q�ď��ުS;�����BS8�8�°*�Co�U��H��+���/�kQn�?,{�5> !��:�V�S���OdF��S�x���Rîqj�Yy��xL2���Iyt�P������#�ۂ�?j��=���J7y�h`�M�-Dh��d�󉯔�{��*v&�b�Pߟ�+<e:�PɩY��t<��f���
L�k��ٖM�pJ���4�Ű�&���������+
:j@��\�)�����g4�~�i��"�����]B�WP�w�9�E�A��0YԴ.����/�m<i��������a��P�O�D�3����9���y݁�TTu��*)[6�9ﳜ�nνL�/+Fuت/n����
�b[ґ�\ǜ(��B�'z,��]��/՘Q�t>�b���Γ(1��۸�1-)]��(;����j-���1;nf��@�h��/VVZ�r	�]a�w�tyX?F�q�|���gTR��2Q�lBN��A�M��w�5C*�Q)>�[�MJ�/b�g�RF�K]��k5�~�w6�=���h��Y�s�8�"y�%���U�r��]�i,���yJ��߿�+�GR�����(`<��>�l��\�
�����S<X�-�M�i~����Ϳ���'�e<�y����H%�;��/ `�{x���j�k[ҧ䞅�Te���m��M�r�ӭ6.&����U�)m����+��o��6��u�r!�{bC�ͻ���`�8��@6ڳ��?��깒V��E���$�ɽ½��₲�؟[)�=uZ�!��:��U大a�L�z�\y�ĵ��í�<�p��_��Kb���q���-Q��`�m6Kxr��aq�`�I�yBl�|��B޻:��t��l��ls�Kwsl�;������ýs_>��5Q]�}6���O�VϏ>sµ�5��d	:V�QV6��&���ŋj�����Z�.nY�
��/&���s�OO�,O�O��/�-�2eP}<6�v��_kfT`��=���<��P*�PI�*:q�;(���+�3_Y"��m8�xv.ܷ�l��HT��B2Wr�tm>�RB0��ʐ�c�b;� &��^����}q�����v���_f�~S�m�/\.�""�.�)I�z��n:#�b��&��Q�R�D��g=B	}��B7ag�Yzv)�E�vm�j��q�t�
&��K��U�@ĭ�؅�`pG��T'�A|+�<ӹ��6����r�:�G�����[�}��I��I/4���F��B�U��1��#e�z%U���{0]���r��Hq���k�������<Ŀ���E��ȼ��㦏����[����Z�#���}�������N�r��@�b���Q�A/M�k,�1�u��t�klQٮ7��~f�|ƒ�n_ՏАZgXmqq�"ޜl�n�3���;�b���)Z�����㷼�{�ONM.X�i�E�X��xVZoWޫ�-��3�"�ps�\��I��-MB0	�įo�;>�#����q~	\y�8�1`���ef(}���5�]�J֎{�����MzZ*��AJ��gڟ#���%vmk�9��(^�\���q%����Tp�O��A=J�M-���xV:+�*�G(0��jkBT��p�v���k�<�tq!1	gI�:��<���E��]+4w��d��,��;;t����*	�*��� Īch��!x��G�{��3�Jw�4;]4��Yȕ�!���w��>�C��m�!��,'��_lM�������m��o�d�����\��q��w1���.g:����s�6�H����JcU��i8;�,�á?#� �H�&�{8t�ʳ]�R�$����юM�}�t$R�J����$�6��,q��9�;'���EۈT�������u\�T���=��_�<wM6�~��u�@$/��}�3����uX���z�ʃ�������88]��6�k|��2�դ�%*IA��������8/����ω9�5��49Cv��&js�h`!
S�o�֘�U^�
�U
"s�sQ�47֩��&�翹�n0��]��V�1�uJD�)�>�\�
��Q9ox"���v�6�w�����v��J����!���D������Vq2�w�9�t���W)a�kF��5��#϶����'[�wN_l��`��v@y�*�Ε\�Y��9����X;�������h���v������S��S"�x�I��Я��r�¸�a4�����J�B��yv�C�1�-�����V�,�����q~����l�K��@6�?�m<m�m��e����k�Z��������f@_��H�mG�6;]s��9t�C>�^	��.��=	O.�x4~���^�����1R��3��i�����O������.�_���?�Op�7��������ǣĤu=ߊ��k����ThnzYE �Z7~�Ӥ�o!��K6����5���/�2q�q��r`������V�\ڈdoDK�D,�"i��n�Oo�0�B0ՄW���s�)~�pt��Řw���8�����i���������V/��T���S�D�EF��
{���&�E`҂"?���1����48�_���E���=
׼V�݆�[V]$V9��b�@BWj��ov�xP���[T�����5XӃ�|�?#��AB��!f}H��U��Jn��%}��eO;w'�,�Ɇ4ZO��<� C\bip�,W.�2�')3�ޭ�����Da]�`���o,]X�˶AѫS?$o����£���s�r�]&�� ���ҊWn�[t~�W�,��<=��*�����̶]\�0����V7�wD��@u����8��;N?Bnr�� /;����(��N�'�#U�ɘ~�E�%�F��>���ȌP��B��Q����wA��>�������V�C]⽌C�����X�N����	��5���c� A�W����2�ru�Y�z�e��4���e�O�z�'������:�xVΏU{��pq��lϠ�"��U�<֖��~*I\�Y��{���
��� �����7�Ђ��j�b�	\��7��~���;|.��h�囊= ��2���"K�C���?��\���(6+�۪S�Ȭj?E���̫��g'��1X\���]��Ox\���j��N]u=�ŋ_F����v��w:�O����oJ�Ѻ���׏ ���ΰ�䕶(�VZ9��{.�߬����^�u�<?��5-��������$'��#��6*58�r�&��;����+���O���-J�X����:�����#.���V�'9~;��M�]�jU���FΛ��;�0�j�i=L+�V�$9yv�T�%z�5��t8\�y��x��'9���I�磗g������1�=��=�]���\Ǉ��� ��kV��~�u���j�ڒ8�q��m��:�Y]5\	�����:{�Hh�6Y״]Az]{UĀ�=��!�|�m*<4�i"��$�NN � ��z��J��K�c�N:�m�N:�m�6:��ضm;�6���/3����瞪}v��^G���߲�ߞp�[eE�?A�v��"&ˮK���v��g����k+���.붱�O��&�nĭ��K��������0�_qlk��b�G���Q��Z�R-�3��1���;dW �^�x@��Lr��l�e��(�C+2x&�8npg��w�:��ˡ➔)��f��y�i��x���ۅ��B�������f1`#��/�4�̐L�%�v<���yP�^���f٦RWuH��Jڶܘ�><r;{%Ywj�>���{�%�]w9�W��M�JqI�!�N�p��Q5�0�r������w+�����K7���QG=�
�3����{d��
��h�PQ^�h &�i^�Bx0\B2�{�Dɟl�p=�voq�^A�}� ��+�ݑ������y'ZS�S��E�Ѱ��p�Ȕ��xӅ]I�khG�M{���YuG�d�u����W��w%9&N�c{�E:T����'"�J'���u�)h���S5�|�0G(�}��]	W�r,�H��w��L�,]��عwB���AB���l�����vE~dO���ؽ���a;�8WQȦ>gn�h���~�+���?�H~	0�n�Jp��6]x��!���eo.��5$�����:��yC�a�tM����!��t{}��w3�����xFz����P�W~��Ol���f�[5t��Qtw!#��bm�S,���Y_uˢnȩdS���!�s�rQ��}�d�3Š�����
��qN��g,��.F�x*]��#���YU�b��h�L������� ��>���_����s�4�>ٚ�>y����t��g˕��,��,�1{���=�D�W.;D��<*C��a����a���ݒ0F)���o:��Y8�5@Q�#�7b8�3h>d�9'�wf{^��lt/�{�[bǶ�"�D�f���lcӦ]��voZ&;��ufc
��c�f�j�+���z=��Hh�{#J��c+�	��x੔;�NXx5&��Ԋş%�.�r0EO������˭��;��i�cc=Y�".@L�qA7#�&�{m�Y<���
C��A!��0&x(����6��P��o·D����4h�B/�|P��;�Y�:zqF7�b��*�D��j����X̻��H�ea�Y��5X���µ�V��0�]�8���wX�(
��s���1��J����\�D����@�5�<>�8<A�S2I�p���ua=�K��##�pm'���ď�\lH���2��h�rI�T��jװ�Z���a����{k��_>��W�e�UM�c�3������t_5U��,93�[�n��ܮ�u���I9˸��jw�9�In�]#w�p�(;30\ea*���@ VTU�YtA鉁����۵���N���Yf�$鵖4ى�Jvz�,�·d�I.�q�J�~��IdV��+F�kR�Ŧh>����������on �Ы\?:O��4�Y#��ܯ�h��#�q�.�j�-ۤ,��F����ײNK���O(���Go2��z�oT��a�	
a?t��&�A]3�S�� %��=GvX��iM2u�{Xi�����B.�<X^8p�5iN�"�5��H鼛j��|��'z	#���lc����0���eߢy��U3V7mN#G_D�bEe���kJ�[�`������cQ`��N����ox���WWm������M#��^^�pl�����5�A�!Wi����`Ž?sT��d-�H'�g�Ğ�,"V�~�O��]��#m��&�ŅAF�(fh�&��m1D�"�	))��:����F�o"m;�54��H��e�i{��)9��1n�@�U�i���gN4��7�i��ӻ_�Dx/�Ø���fO�e�y?�|%�e�k���S�T�[&��d�,�1%�n����-c���b�x,(�(��C2 �f�<�+\白j	��,��W�	���Ei�s�� z`9s���{)���q�^kd�;PL�~esv��vڌ��S#���%���D�����_�P9�!�ĸ�.�2���[��^�М�&t���d`�_�d���;����9�4��'�x�.>o �@� ۼ�/�M�E�閄�b�>*O1��	9h7��������֝���{D�]�aS,��� �ה � <6�j#*éh
��(��I١�+,����+4� � bHH��A�&�,���=�V!6��F�&��^�A�O��'�'o#���J���݁�K�f�,D�*��$�C9���)_v~��a~�/�~���ݷ�2P�ϸ\c�Z+� ���|&�D�d94��[�ED��#y�75X��g�ʹ`w|�q<�i^�F[�����AA��~�39��]t3��N�ė��2n0�K�_��W�u��!�갮׵�ǌ�\�)����4�M�i1=��s���q9ީk1�-�/^�=<��y@���7�io.��?̌���{�ƨ黭��_e�1^\���Grs}��$<~yq��\o�č�>�Jc~����
�xܦ���?�K�����^��Nb�
���8���q��gL�r�<�6�#���㨱�r�l������=��.74�	!�(ez�Dt y�½/��qo��W�]MQ�~��Ƚ��?نc��ۧ=�#z�a����:�b�R.ۤm�?\�"��i��*o�^������}?�^n���=��ޮ��\��4�u<��F��Co���~��1J���d�{g���3&ϋ���G�Ub%�X(9����l[��#x#y���NK��!#��<B2��cz��N�����2B�����A�[�y��>Q�{>x�'�_�Y-U�&��yN�վJ�<���9ܿ�g�b��(�91�(���A��@'����`*"�_vfw���mccT����q��~3�0�U����:S���'?����H ���}��%}�W��*,J����;��/H�4qU��&�oռ@3�y|��ޛ_�?���y�{���oԉXX#�d�5�$�3��6g�H�Z��<2`���-�1Ԍ�}�t;O�=;�+5��Ze]���UO�
�Q���>�m��y���=m�Q�t�|�?f% ��j.[,���M��G{���
��8�,�&������������>=-���tۢe�r����+�z�fa�`a�%X�4'���.�OKؿ�4����}5��uZ�/�u�?����7������2ѫ:������+�b�F|q#���s���)R�,f���X��� ޮ����I��"�:��I�R�Y��D����:���dbZ�W e��Ԅ��t�R����P��v����&?ȋ5h��y\��7w�l�#�;!ȘP��1�P����_�p)�b�)a�	Oi�C I5+�5~��W��bA�~ @k�qWD68.[�u�s`Ztx��8�]>�R�:���N�E ���^r�r����	0���A�#��y)GyK��}����m.oa�ym.��e�Y����Z�R���:��o>��\��~i��k���W[e��8ev���c��O80�q�{f.tʨnswg��]����{� �Ȋ�t��{`h�٭���.\�K�����l���s`ck����G�z���E�����Fl3A*R�y��4Ҳ�b� U�P��f�X*(E��V8#RD����e���l~�*�ޣ�B<98�q�0�]0��� �p!11�#�	��f�n����j��|p!X���l�#M��.Β���8W?TZ�
>�I�oB��Ǉj���,N�@g�tİ��n�ᛟ��M2=�4�w&/�v�u�\vL�O�Vի���[���N�q��������+̕��A�|�w �+F{���pku�B��罞.��6����� ���C��#d&�W?nla�}�y	]��/���rgx�;̦s�c~����V��6�S�MݯC �w�11Y�¶0���f�_�AY����>�̰� U`
����5�A�?{�U�*^�2@%"Ƣ�`��I���<)K)7���t��>� z�?�BR�PZ�����˚���7�8��~�k�D]B���d�I@f�H��l�jH�Ug\�cĠE~��B��;����ɕ���8�z3�Fr��V'��Ra#��F!�$�i�~i��'�|���Ug�z�>�c���J^�t+_�J*�r�R!��c�`�p�f�ak/&��N�x��EDz�1D�����m��i�-!_=�s�yx�\A��m��&�@w�O[�7&�0E��z���Z[�s��QH��j�G�G��P�B�E�u��0�P�<�- إ�*N����:��,?ZK�	��ˊ�A�z������G0.�{���捩�k��������IK5�F1�qq�eflt��Ɍ����mF�@]�T�v#`_�Y���{��� 	���r?ߩul�=,,�j�J���I�:��r�f�OA�4da.����;+��s:�d�*^��#�3�l��}�y��%���H;n�<�����G�Y�*eEO*r_�͓��	J���r��t���AB�p��R_��&���S���d`O��M�j��� �����Gַc�+��;M�)3�M�}�%���[��S ^�l���(ц��>/��Զ�+~����ۻ:xCj�D�7hmf3p�@�I4�"l�<���sMk^)9�k~��Q��0?�1�ݎ��g�]2%7��z]zh�6}^=��xrL�L�<,�[�
ٌ�,�F�`��/�`ӝv��16 �[+Pm�쐖�s/�m�7{�i�O~�'������9��Τ�f�55b��)�`��	���)�)�k��Ft�Z��2"
�$d�<
,��C���!԰1�����+�
`��r�t!7��)&��0i����o�l�>[�ߨ�Ǹ�5��ڮ���u���^&n�Z��|�]��|Պ��L#��\�nm���0�ˤB�a@�����ä4
�y�pX��QB �rh���ID&�HKWm����Ыw%���}�T��

���Nw��L̍��Ѐ�@���
-d~!-���z��R���;M���`�I�哝ԩ�l�6=���K��q^~c��F��yt?��x��S�4f��=~h�x��?:3����i�Ju�f�̢��7�r�ʂE޳�ʜ�>��(���F���T��"���b�O4b��5��/�$ywMk�����R�h��*�������f�^�ym��Ⱦ�Ԭ̍�d��p�e�-{SN^�86d�l��0,���v����~��	=5�@�'e��JS�Բ�^S�L�C:���0��k��7e֚�WB����U�O��M(�Aσ��$�d���z������)��-���;�a�Ԝ��+��i��Eq&���m���knn���M�;Q�/i�%Lj������ ���
ڶ܀c�Q^�7�Qp�F�1�9��>8~�-����(!�y>d�&��y讙��{��J��>�f��v�!�͈�V1����ծ��Pڙ�	.R���7QBL�߼P����� �+�<�X�W6�'*�ߤI�D���:�����Ŀ�f���|�����^��>�nn϶޵|�sG�}?a�w3'D0�>�(�
�Ĭ���ͷ:�b�}��d�$郅�/��=��><��|�)��Ҟ;�����G��(Q���n�e)�8��9@x�toOW���6N�'��{"���2���&��ͅ���ƻ�"�ݾ��"�oǹ�l���a�B�o�Yz��w�}>ݒ&+R��D�\:��c�����_��[���z�vf=ɖ������γ*nx�nN�+�����?�|���BV��?�DΚE_�S��OĐh�lHg��o�����l���c�������n�����1'��؛d(�����|gO.NTC�v9�؄�E"����G�2k�l�8í� �?-����9��������ރ��FQ����ɏ̮�QY��F�������<7�8�sn��H�P;�,E��+�;����f�B5��0�L	C(A&���ǘ�E��of%=�:���u����3��f�5�VS��no<��7^_FO���� �4j�����G��g���S5,"T����t����䱆t�W@��b֕h�7����#>��3��J���k���I�4���r6՞L�3�\��e!èx�v�*W�
#I�P�a��>#?M��撷KLޮY+~����ܦ�-���3�����m�m�`�۶�|�Τ�B�~,7��iw��P��f�y���'�l�!w�PG�����fk��e�&W���jW�䏒��e�s�p\aa����25#��Rj�~ n����Ь��B����I�'�7,�H�c����_>�>5?��.���������S�s���n�! hJwc	,WTM�Q�<���up��'//7>0R`��"�|��Җ�<[~q�.�B	�%`��/�_it�����c�H�5�2P"���Q�������&ڀ�$���͛E0n��G�n
x�:OD!�]���Iݖ>=�2�%��b1�n$��Z���{������%���\)���`#�ܧ�u<{-��D���u��'l���۷��ZI�l�W��'�jI��\O����@�܅����k`�CF�~��$��%5�RFb�>rz稏I�SY�ǖ�SA��6F�����t����paryi�dM�KOʨ4�!e((��;���ϗ�G�`�#��®�!5f�v?�]�;/b�L��fȎ�S�_�i-��'�N>^�m�n��yk���6��]�6�vfgϤ�~P����g��*��;7~�/$�:���j�J]ǥQ���0��&�] �P:ms|�R�fh�bwpci�%B����av~gB1�<1�GZO
�H�N�/(bh��q��$�������q�f6�`��m�;9Cu���h�vT`R�lք輀��=(�p&�x�f}�Lp�!0�oAj�z��O���᫬����+�'���N�[��Բoy���8^oDe2,�rX���(��f��Soy�1����'+{�Ǻ�����w�My�Y��u���u1��z��ȘM��e���iKf�w�OaS��%1��2�
�H������m~Ԇ~�͎�kG�� fX�FFJ�t�-�[1�E�{y9���y�^��g��O��{[w��d_m
z�9 4p\;��c���P_���q�����2h�i��C�XJ7�)bb�71/�C����F|4�������~��_u��Q*��L0�*/&���<,.2Muܭ��綛gP^��Ή����N��B�q��M����;>+�7M�l�k\i�ӷ��'�ᖳP.s�.Sh��k��DQ�0�36v�c2Ek�Bw��f ��م܃���V�qY����īa��#��Ĥ|�]�l^*
��GLŌ�:�/��=�g����� ��8ߛ��z���/ ���:��n�dR��օ�2j>�H��?C�J2�2�+u�����N�
�8�V �G]b>;�9.��4��;���_C�w��3ȁo��%S��&�ATH4�)�K̺]pJ����ͪ�UW��rR����F��M8Қ]V�ڼH�gII;�j�<� ��aM��*;�?CqV���f#�/!KӇx�,XJ9�"%D��N3T�I������7��=z��z��g�(JH���/Ըt27_3��}��89H����u���;�(;^����K�㵴�x8��(������3�7YB�߾�x�ؿ9_?�a^��߇�\4}�G��,N���Iا���aqK���֚�Ta^_�5��J��!+_��EZq��.�p�Sk�7����T>�V��b��g3ݾ�oіJ:�h�����ͷ˔j���ۿW�ꟷ�_s�^#O]�[�����z�u.O:���KX��s��k|�Z`�}B�صR+i2���z�y�Po^���6ު�}i�N����������J5@n���ꛦ:�zY@L[W�r�m���l�x�=������2wR��3cI�2��b�x��a�ӄ�_��L��<��]�λ����!���Y�SB��idi���	Β���>3�w	��-�ss�4;�ǴL�q�J0(k��>"����/�g<���193{~Mh����͏%�	 ��201P������ճ'�%x��f��m����+
Wg��B�SK���
4�����>Я|Ϯ��;M�J� �N� x!ď-(��4�$�%�2��bl�5;3��7�\��oC����(! �pCmxT��d��&�b7ļ�ƅ�$P��j���!���S�0�۠Q�y+R���F۾���{�]SbjOw��U{�N�\�>�^<*)�6dz��^��玼=�����
��٥q��#�*��6pP�Zz���a�j{��k8�
�i�Sh��W��`uA��������S(>Y�^-��JR���nkG��M:[��C��8��=S4�j�tW���,�l�yH~�p�	���t��AkpZwxu��O�K�'"^<M8=a����|�!���\�=�s�	Ȕ�,1R�����2�8�y9T��B�D�BdmX+��,L�<^�w�!����ed��&�]�Ť�+�.qޛQ�tw	k���̌�s#p�F���Z�?Zw)߶�P�!�3�C�\�a��?���章g��b���_�H�%�VRZA��3p����w�K$��b��Ǧ{�-_�Ӱ���@�$Z�B蚃a�ԏ\�j��?�?�x�C���~�)���i�E��Ѥ���E�FH���VV�՛�]�>1�;][C+���c���gf'�N�jt��}�@�̏�l���f��͈�[��_cz��ΒjR�2�$��U��X�������G}W�κ�~������O�M��������e��ے���]@��3*-�H"n�	�*`T#���]���s|D�Ȱ����3�Wn�%��~����I����kl�Y�#���)�S�0:�tT�8���R~9@9h�%X�F$_� �>��3�!�jþkamp��;��t(i�T:U�9�,��@�Lt��r�_�Lp1@;Ƴ沽��k�V;T�0�"��	 ,�$.�-�J
ʥ���b���)�z?�7]0����(��7�~�}�X����*�S���+�Nw[9�Lv��N����%E��/k$?��B-)�ㆄtx�pU�'���~a�ywp �E0�#�11V&��"����u��R�����W�E�� ��zz�iL.�%aO��z��	Z�~�^*�l,�gٖ��@
���T4�"(S$�ж*����o$�t��p��C"	za�bE
22i-�EH���}��Ĝo�L�9j||a�\��$�����M�E��Ĥʦ
EFp���IY\C#�re�x�8ƘTC���d���Z����b�C��E�!���"�F�{Krw 8�h&�LV�׺`v<"�P0<���h�dP8""�����}k�%r���}iƾ�ֺsR�/����Ӑ�q�W�_A��K�4"x2��W�mL�]��'�lO!�;^���y�Xr�eo]"^��.A�sS�`iI� ����XY�$Y��M�ՋF��W�1���� �ղ|�w��|��
���}��Z-���mρ8�o�zD�8�4c�t*�[�jo���@�B��0����@��c��=���q�Z�	./�{$�`,nX��r�_�IGvNj���M��pI�IU�P5�Kpvq�pS/>-�����Y4����
/����?/�Ǹt@<]�KR��N�
>��D�,�)G�(�f�~���?_ vV���-l[t�I�C@�g�W��W̦�ғߠZD�7�%��t�$K�t�#�!kz��A���ǌ��eA)��$��?]�f�c�u�?͐�As��3�}�K'M�-���<�x�����֤�=�/E<�z %�SH �:�:��&�� 7b�dg�.)�rV�	I	�vF%8=�@�� ̑� �n�(�PGW�
`R�^{��?1�+N�0B��Ʊ#,YNy%��M:������*[x��nԊL��v���� ���ς�L�O�z���bV�����urh���)01���'PDr ����)�)�n���+����2p�a.r{�dl���e�����Q�[�M�&��~oS�*}ĞX�^��|����L���ȣ��t�R���EZ�#Bh���P��{P�������o�d������(|9�͖is�;��^MԈ��kU�yc	Ym�G!`j�j~�T��]�� ����h.�KP���=� 6a�����.�`OI���@��]�36���h�B�R9�f�~ͯ�CK�3�����h͔p9�&_���a�w��^�&1		~�/�[��R��(�k��e�IN���)�bX��p���b٦1�@�t!�J�=e��突�Yl�[���c,*}W:��KZ��|D�ՙ���a�k��S#���#;Ď*.���X�yK�OZ0�O%j%�-��B��a�\4�]Rϵ��B�	b��i��[�Kؿ�<x|p!�yd�<e������(`�t;���b���ۦ����"�In[>˛��D�,���SZ4��}ޛ�z�R�2Bm���R-�=4^�V��Â�q���'�
�k3x�h�pUA���"eɉ:ݦ%t*�J��b�]� m��Z����Œ[���tZ�r�p�Y�T�����gFD���1\o(����/k >��~�����
x�j�p�>�g��{1��4��X�|PN
>nB+N/9OO��8c^���6���
���u-�����㮫�vs�|���I�[����i�U*t׾�����p�1�=�1�;��{�c=���fyH��P�J��}׍�?C;Z�١1��.F�R�Ӝ	:����יd�"���]��x
uO��d��f}F����iZ��n�Nvx8�u	�}+��z��E,z�{V/n�HD
�3(�߃�~=��X�ЖYk��*4���FSr�].�R�o��yr�����^v�D$����{��u��BtX��v��Հ�z-.�˹fhCz�
^(�^�������Zf�k��04b��'`/�m1���p|����k���)����l�Y�ZԔ���@�M����\W��"m�qY���B��߈4n;t�TS��h�g�'�s�?�2�������{ڛQ<�'ُ�G~�҅�52��Ci!o>,��5{���{��x�C���sp�@�ݰ��f�C+*��� ���(Vgr�:�����������'f�+J�ާ.�<�W�b]������Ⱥ��WC��g�a�TS8���t2��ِ��M��8Wooͅ����T�!�r\�ڠ�A4�9d�(r�h���m� ��}�$.�0��@�s3L���&�R�� �%ֽFI�?Z	$����EbB��ާ{2���w'�ge:��,�}�k ��G���#0k�υ���i�*�e:}6�Qԕ��TAZ�^]ׄm�~���VҴ����Y�&;\�޽��:�˚|O<*��w�J@�	W���� G���I�� Mn2zX{�I������شIdB���s:�_�ܴD��i�X��ڭI<>�HшEpM�Y�Bo�ȗ��?i[�����
���3R�"��(A5u��P̹���8Gm��ˁʻ�Y�l�
�'P+K%��VN�Q����%L>R7����qf���߰�;}�(!9����|A�`|�z�B]�1pN�+�sX8��eR���0��醕^�U/�D[Ǔ|��mT��&;/�U���t����Y;��L1xL�l���@�a&�\�pF]9�:gÂ���ׁuL܀vM�k�C�Gl'+���הh ��D�~c^��8h�J�ł3�G)2����������?�Mt<}N��1�>���I��ʓR�Or�%c/���XYW*��1]>P�W|֔���"S�7u)�0�!��t��h��z#I08��4�~d�s�O��vb�P�j����(����t��y��~��$�JxR5��i
eY�4��O��e(�q�Z��M�dެ(���C�ȞM,���}�dv��0sk�Ֆ��Pb��<��2�Cl� �"K
t �ӰDP@�r�O��p!2k� �����V�=!�r����O=��0k���0t�������[�Q����ڝ���bkb�������Ҡ9ͺ_Dx��0�:�tĔ���1���[����*5%2s��	��Km�� �Md�ɲ���~d�L"�@�c��������dR� ,tC�&�#�h��d�Lʭ��NA�XqLv�O�;����64Q��R�XCI��R@,��/C�{M�C��3Ɖ�*bI �M���(�@E�(��d%�<�Ÿ�,
f��}��?J`�ةbq̄i���U�[E�d��Q"��%�҈��T_7�}kOm�b�X�G�bd&G�����k�d��P��Đm|=֏��p�d�R��0�,�E�)KI[�2�UўGk@��v��
R�aW�Q؏�q7S����]���gOP; ��3&�ȿ.�T��L���`t��yorR�1X���)�w���4�p&����B���g�����I��5t��;�e�׀Y��'%�ʐ����=�	/�S�6vR��/�k�?p��Q��^�j�L��;�D�2� 2�l�����~�+eg��t6����m�b���ˌ��J�����^�D��8�Yb9o[�
4�a�K���	�`F}�g[Q�D�[���')|K+����wk�E�����H�CL�3\��!�u1��u��ҏe�Np�әV�%�[�[q��D��B�v�l~��
�5]Y3O�d& ���ȇ�����h%�E��9�MHR���Ky$��S��d�2��D��N;�~�+a���O��VJY1�d,h��W�&8l�L<O����h+��f��teI�ݓP7PP1��'���T{H�3	���[z*�
yi#3�i���P5<J��cE�-Y{ku�$�Ĕq��WǬ�f�z7�Y!��``+�*�$���v94�Z�Y�X���I/D�ŷ6Zu~��r7����CUa'&&fk�`o�j�;�;i��*���ָ�>�fQK�ϛ�Cm��Lxޒ��"8���
����Q��/��L��?�R�7vWb5�M	�#�a�HW`�p���-%��m��zMUF���|�342���A��S:�� M�,[�P�(�)dmܿ��EP��x�}�+�PL_,� ��8�T�env��c�|[�J�r;� �ih2�R������Vq��1�P_�J�-!�"~`��H����:r�ո0o��tt*��N�͂n�p�FT$z3� ��=>d^#v,A�τ0���~y	"�qZ�(,�rɠ���@��"&�uo�/�2Rѭ~jIq�0g7Iq6Y�1�r��a?�8�ܑT�V8>//���sq;P�=R�U���iOa�����|S��)^+X���04@���������l�C,�N���6��#Q0��}�M�ۚ(q��b�zԤ���쑌;�A�\/�*ч���0����k��	�$R�p5�؀c=��$v�MV��f��^���I�K�H4'CL(h$퍇a
-G�2�}si4��rpQѪ����Ԃ�#팔a�^�b���a��H�845�g8g�+Yeb�6��q��`��Cg�׷�vϱ�eY���<dTC�a�x�Tgi����j��8mh��P4��ʐo��8̥m\ܞFz��O󴙨
�_	-&���]Ro�BCϱQlR�)��-<��D��c�a6 " XF �^W��k�%Kɿ�A�a��G��/|Qc�w��:�f�gm����o��l���Ё���;��Son�f���W��2ᤧJ����\�I'_xN#+�n�P��V��sw��c�J|�;]@�f�zP�fa�V}Y����xpB���n���(�4+����;ztN���=y�ti�>������2Z����{ܔo1?��&rr���ǁ)(�)tf�\4����F˫*�2D�������fA���X +d����70�)����ي.,��#\	��V{�0��BZ�<�5�i�-5K�a��f�k���t_ߦW����+.�X�3%�S;�I4��������H�3Rf�t���%�Ob+�g5��I�:�$���LJ��b�)���n��L,,��X��L}�|�@ǎ��#�R2K�$T#z!�"*�.~�p'�e}����
��Q������5����Z��i# ��'I4Z�;��B#��>��:	�KX�)r���?�����Kvi4�;4�i�v���e4��ɘN/uƇe��΢�J�8x�3��S����-г�=ǋ1ڎy��Z��#%3���b�����Ī�X�F�P:�&���ϫ	āc�\c��WyB�n�����[VD�_i��^�'n�
{�p=�3���B'[��|�r0#�H�ǝ�*D��H�_�f�Z�<���ګ��[������S
��$v�]4�d[�̐"�AˠO����n�XB���R�-��j�J�\7�U+��`�r��Jg��d)Lgc�Y�ey�o&��79$����R�!Τw������|	��e���m�=�>��( �>�Ӣ�J�ĖW,P	�F�A�^Ws1zq,��0^�%��G�rM�8�-I��u��Y<�b�|����]����F�62W(MKİD׌9bvH�٢���y��.i�|9]��^�a$�V�c <)�K*8�Zщ�1���a�H�e�ɯ�[����h�9�U�С�%~g��e�0��A�oX�VA��fj�V^��l稠�BZ� P�C��*�U��Y�)�;�9�����Y���Y�.ܶn���~t8�z�����Ok�,/��:�:�X$�۬�F�W#D1��_����H��1P�/�w�%4da��@���l���i�"xH�Ax���kNja-�Z� `%�i�^��⇡ b�,�~���4�V���^o�چ�R����I�����)��)������"�$�~���BO���N�K�p��z`�����\q
�ْ���Z	�
O�&`�ʐ�D �-��Bq��W֓}��V.����.�f�ܥ�L�����D���8\������Xx&�
�&؆֩p�'M���F��iq	��.)��P�X��S�B�&��s��Nc��s"���wB�1	�A�.��^�������H��~��PK   �EXN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   LYEX�cX�� 3� /   images/9e507620-50e3-4aa7-a16c-7d7ceba17d8d.png ;@Ŀ�PNG

   IHDR       ��   gAMA  ���a   	pHYs  %  %IR$�   ]tEXtSnipMetadata {"clipPoints":[{"x":0,"y":0},{"x":273,"y":0},{"x":273,"y":790},{"x":0,"y":790}]}&7-  ��IDATx���i�e�u%����!���ER,���nY6�4�0�?��a�À[V��Eq(�*��r�9^�y���Z�ܗ�)u������{�9{X{N+|����WdV����у��گ��޷��o��_}��%�s���nl�����s���k���=c��_��T���;�1���|��~E��-�@m|�Q�~�ijq����{�8���>g�[?�7�����SC%����?���Y��x%�w��\=���Ϗ�<di�kb�v�n_��Y�n�"�L��_F<���dʨ���c��/��}���g�뗄�w��D����P��J*.H�83���7k+�Қ���5��~��L�(�����\0��_U����E_�CQP�w
�*��U���;,D~`�,�$}k"��U����6L?��ϥ����%t�*
B���k8+��>�d��E�0J��� .�n-Ͳo�zx�8�b+�=x�z��Z��lY��Ɩ�n�`-��Z�l��@�$�G��oq���/U����k�b-���<����~�9ֵ&�V;�ǵǸ_s-Xim�fӶyn��׶a?~�ĺݶ-�k��$)�k6XK�k��a[�V�u�m��{�^��BIF���g���Zx��ͼ��V�Ex-����8�|�cMM?�8�5��i?(�J�����C����g�$��H�P���
��{�=���¾�Yd���:ݎ����.+��t�f��A��L�Sݷ�nk-���6ۍe\�A&�O҉�M!�u�9�^��k�Wkk4�h�;� ڈ?c �'E5z��-�@ӻ�ه�K���g^�SF��!z��;��E�/� �g Ĕ;͵7<w�S��v��CA�W��#�?�#pC����p�������#3��؇�-=l�ZT9n埭�"Ȳ(ߊ�����҅�f����s[�� g�������xX �S�v�\X�ղǏ�`����݉ث����ޖ��u:]��=�n��v��j���l�:$h���65�V����.};�s���j��`�u��k"��2�Zxm6'Tr<.��u>���m��u�]0�
ϰ��w��ӿ%$� �ʝ ��}��CtGO��0�=��~n�߿��-��r��Z��:
���{͵�~�`�Φ��Q���p��Oh��KƉ�Er��Lk��L�?}�Ժ�X�*�����IE��������'z����i��Dᾥ�V&�������D!��ᛟw�*% ��n�DG�w�ݒ���vzvj�|�5:�^W��.��Y]�8���������[5Ue�f�/?����m�����.@38�*Nd�IYn�.
�T�H�����=����F��v*���C����Q��W���X�b
�~� -DδUxb\���a���D�D!��	������{0��5CJI��1����!K7�4m�p�p��ڲ��ۑ�N��l6�'�g �5���mi���FS0NcjI�q�a��d^%��liϟ?5��*hu�E���kc�E���C�ŀ)���p���pD����J�	Q���V���Y�g/s������ >+�s~7��9^���~^����U5���C��S<�}Q�JQ~����^����N�:�+�|�B�B//b�1)����㦥RI��}s������g����ԲI�&�֤2��f�[!�#��r4Q�:nH�S8��))s� !3��������D#''����� ��̲�P���=��X,6,Yړ��N\07�\	{N��6[�3�8��G����	�b�����P�r͍m���e�T��Y�Bn�/��FN�$��g��:��,ue�ȱ�>5��5+׊L����w�����ë�5Pz
%V�m�Np�<�����M�`�l�;ɥ�#�����W�	p��+ ��W�pq�Í������{r\i��� b�*�m�y�D�����^������e�Z����\+�� �ժt��dB�L��ڃ��6.@�$�~s��ڦ��٠u`=�G��e��F�N��|h����Ў��5��viGfD�"䄨��
�?M��~�D�A��-P����BQWd(h��G�[�,��Q�e ���=�HYm�v������IA�m�G��Q�N�3{w�����Á�jIm���Ȭ�ܯ!��X�j�M.f�&�l@|	1qS�(6��a�s���3�k��s-�V*���ϖ�|v
B�&j|�kD�k�9��P)��hK K[�C~����-�� �|�{R8lq�|�a��i&�;m�R�c��ӌ�N�i���s�X��g�C�^c�T*�~�\(P߼{o��կ-�p��b�L<˚�/jI!��������<�3�u�9uC�@{�1�O�����f���;�@�/+
G"T�VI/-kv ��̳���''�O*��bo#{tvh�~�i>r�y(T���Q����h����f��X:�!��),[X�\��0�����o>�&h��r7p(��|[	Vf�=�4��݀d�D1��f)A�b���F��@UͰ��v{ Қ�I�DI0������d2lHLI�q/��\,u�|���s�9Eۺ�����g[ ��`~�K^�{vA�a�� 3���xo�Acgv	7"�-�jjJWZ� ��L	����p���6ͧ�"$1J!X^# 7E������
�͚��H3�X�#Z�ĸI��z\�����t!@I��a&��m�M1���|&G�Y5��n׶?ha=<#WU���s�B����j�y+1i���D�JҐ���L(�W)��W����F�u�} F�F2�'�Z'}#e@�|����5 ��_�ZH'��t2ճ�8S��Zo87�'׵�����f[P�
�|�C	�!��%M1��p��P$�@���Z4�&��yy@fb����B�#E�29
�ܜ�� ��+��\���bme�~pڶ��kv�S�c~���9����[{{=�m���W{����P[j���� ���0�Hb���CM�g��U���#�x8$(0��T��	B���)���Z����ԣ��l�P��z�G)�i��t��!��v����GԶ9�(<�.`:	a2��x,��N-P;�� �'���E��������m�Z$S��K�ʿՌ/����|om[�q7B;��%"��.�DI$&^�&����mP����.��A�����F��-��(�(p����nI��s���/�{]{}�m���g5w����b^"��� ,�P�e���7�v7��"���?<~b���@`��=���)J�����0l�� �C���J!�7ؓi�Z����#>�������g�4��'��^�w��u:
�
�-Egý=	��b��s��X�3��t�Z{x/�ω�K����֮��*�R��H���wv�{�����2i�
�������A��S���6Q�����>.=�W���lb��L�K>�W�6q] Z�N���nn�Wo���I_O�C4|��'d�^����b�( 6�9��ۗoo-n�J�����p#
..���W.���1��w���a�4�_���0D
-ˁ�sHZܤ�A����ֈW���kG�`��Y�vྭ��&2k�m�&֚��p
�Ӕ	����������̸^���ПR;��FL5������ԃ�x���W����B�AB��QBx|o������xarp��m�A���=���d�����tt�P#�^ϑ�=j��/
*�M����s �`,bt�Aa�����S�9*�Y�g9�
:����)��OS1���1�{���������r6�F.߿�����߁6����j���4)�{O��g���Xs)$Pɠ��ܳIR �&���}�.Dj�zr6о��|�Z ��e�^�a��Y�;B�\��}�"*"�9;;�ω>*]k7���[@fƣ��π:���P��)��l-���a<���w�E��*���U������_�2��3sg4���s4ʴk���S��s���z���EÎ��t^+����U�Q�5`�be��%�M`��l����n!8��7�_�A)���� 咄<T9���3:Pܹ�f�����#�-\ VU1����{s\o��AÆ����G?�>¬���vx@�*?�T�u���⺰ua�p]	6rt?��l�'��Z�Áx�%�66՚l"���K��`������{ݶm	K�JH�u��!zԩ�Ą�ηi�ʹ�OF"|�����G*
��X>��F'�z����`�ѸʵGܾ9̰	Χ�����N�5o6]P7ҵ�9�����?ٷ�?O�B�A!&i����� �]�5�z@O �&c{���D��gT�Bk<{����)�N��f��Ρ��˦�Bhta�$X����͹��gVv�.�C��]�W�*�m���	ٝ�Лk;9������ۖ/&Vm!4[Xc�:�Z����Tr��c-������O�-�r� ���b[H��t�˕�����9
{�nt0}BـVxo�[�ͧ��7�sJ�S�����ܱ-�&i�Ns�z��'� �BT�g��ޛݽ�G0	g���/�o�r��5P����&�#S�6UkA�&��"r
��`����ڍ�r���m�w%�y#�5k�M6�
����)+�F���x�F���_�~t^n���ڃN��BI�ډ��G&�(����v�..B-J1��U<ס� @"0{��#bhoB�?K���Q3|��|vzf�m�? ڸ!�.�S�-��f���:#�����6��RJ3^j��Khl���ė����Յ �K>>9�?����GO�Ё ;+�G��,����j�9�`{��$�6����b���C�A0�[������o�C����U.�'�L��"��	�v~sm���o.Gv3�@��F	�\9k�,����g����u��;���	؆��0bKu��t{�� lN�H�����;R%��h&r�oI�e%�q�zΆ�YK,X>�,%,�F)����_�_��+;�A �A�x��~�����_��F/l�hW7�]��f���3������>f{�}��Ff ��|��Ԛ��M�҅[���'�̤�����\+zC?M��6֙�2��J�����~e����K{s�g�v[@	P�|���~��Ӂ�Q��uvЍ�~���⭆�G��!�C� ��u9��>VAI����ۗ�s�BHO@��6�"͐�s�<o�?Q�2<_�o���"�㚼�p�����Pt?��6��y�g/ <0��@r��y��5���~����RN]#R�@bz|���K��h#�oB_HD���~�
9!��Z�*CIrG(D�z.h<ν-QXB:U`���8N5:01����>L�0IRɣ-�C�1�84w�1ch
�-��~2�r���D|������T�>�]�	�.F6].�5��/��}���~���R� ���'���;��"4��̿��!�68�5�͐泥-��f����{�-sAfPI۶�݈���)4�L�ϓ�d��V��_�xe����ce�����������]/��5�8����_���K�ͯ.���H�q[jr"'(�-�η�Ղ���;�����-QP�Ӓ	��%�M"M|��	�?oo�%00�ht�f��������O�1���#�L:�#�[�^f�+ �%�b9�X0���__گ��ُ?{jG��z��X�C��>���=0�,��r+aJw�4q��N�[DD|�1 :��h�䵉������VGZz���g�������Bɍn,���Q\J�e���<�iN�Ot�=��Cg����^�zT5��0k��e��w���t��[���#�hƷ#a ���`��)xf�P�pM�`��o
_�^�3᪐=��Wp�5�sJԋS��)�-A�5��'Ǒ?�dX��])a�AT��%�Y�$j�t��%�%�pj�56g[z���$�+C.<�9��Y")��)G[�ζ�(��*)w��8��2F;6
��;w�~Q�N*�f<��=�x���jg�߷��ۻ��)�i��ZSH�)`4Z�d��&+��,�~Y
7�\������PL>_����bS���~��~��7"���}���ݟ�o���7�$� �3��!��+�N!��mV[;l*V���^���2@�?����ɀz�.�������@P@��Ax4���Kh�%��z�g���@���&b�"�ۛ/�����PUL����!e���3-a���4Q�r��3��z~D��ids騣�a.�=���d� ��8+F��`�=�p����؆	�W�B.įF���/����?|��^�|!��b��|�h�*kk��� %��3�p󯎜�A�Ƶ�R��yp�R�0���kW+�
���s��m�W6�9�N�E�:�����G�:0����|%̄	Δ�-~��HҎ�������l��z_�ꅽ�xmy�(��D;l���Y�Z�����?>�qѱ>�W��d�UZȷV��S�o���Uȡa�f�"Ey�cn
V������;�G	ϵ�#!��H�ɓNVjH"�N�h�W�}�� ��HZ���'P�	 亴ï�wB�2Q�1�h��I�N4z�)��D��Q� %���?e`�0B>�i���["�.d�3��ĵ���!�vv��E�?�������Oa��Ʀ@���.�r"eX�L�(�7dP�+9��t�L0�Y5�{�w����1�iN-��ͦ��YAX�����s�P����c(���fХ	��=˶�����Y����n&�TE-�_�:Ki�� �?�e�����2�Lf�C��l=����uh�|n�
�&ϩi�k�}F��A)�zh5�߉^`ʆ�8��̀�ڃL��ROL�g4��pT�&�D#U��~�u�Se� ��|�]%.2Ϩ�qx0ĳ��F����T���V�.��z	!��a-`Vf%+{BL)�&��{m����S�^�rB @IkY�s4*�YX���4F� ��(������&�6cO��k��d�g�'�54�`����0$��#�=�&�)��&/L��#�6-2
���vy�=��K׮��Q����$q4����c;���~"��Wwnk�7`��!�73h0���?Cܛ4TGܚ�yN��(������Vᛨ8��0�Cˀ٩kQ
Z"�P�B4u+K�����35����Z�:QJ�@����#�Pљ�/�2t"�A�ah���Oq�sp��h>%�"�d�SRIj*�{큲c+��K8�	���K{�=���[	��o�o!Hb@����
�
�_m�4#\S�Ҥ��;��\U�9��RLJo|!!�nd��fNb_���W/˅�6�7��Ɂ*l�K��[Ţ	]b+�х$Q��r�z�;i@C�4�ri���
D1�f?h1�!R����lyfh��չ�1�X<cд,�� ����^B"ii����e]��HR����KbAX���r%&b���R˙��$3�c
w�3�B`䴏{����+_��i2� ���Ig/�"�3it�۴>{
�B$��=M�V;�!�:%�/�ƊR(�qN�S�<�s-�BN
c��)5���O�m��#=#�d�)�+����a7��i�Z��$��|w�컭Lʮ4�XjV�e~������Z�L!wօ`d�BF���9���h%��Z1�;�Ğgt���?���f�@k_}��&�mK`FU[��%�
&��:� �+0�#~��ȝ�r�׵k)�ʇ��=w�WR�I��n ! p��-��p�b笭���FB��)��W>W�	$��d}HAj_+�˭��>J�V�KR��
u.̴KB�b���%�<��r&fH�@$%KrW�����N�&>� ������8�Hb��TIV�ȃ�#t$�� o۸f�U������$��us'�}�L�c��{�kz������$@jǬ��1'�� j\���-#�>Lc.#������R�s:mP:И�o�i������;m0a��U�B~D�-&��0��W4*�̭�(ٶG�8'����V���F�6+�EA��ԡ�sP
��� ��gC�N��L�"w��Q*��!�WL4������˫�|�*�V����.�[�=��bϘ#3�{���.S�!P&�D��"Wi��K���"M�O$�h`�����ԁ�za�)�r��! V0E����vh�iTS��Ό��iz:k�ZM�BFٔ������m�lg����<vysg[0��
�L	�D	{4Gh����G��A1���f[.���YP\s�)}5��S�-����nco�����c�d���.(����d�μ��id�\�Pzj��"QKY��*�{��;)�>��c�3uE��v�+�
	����),[�jK� ���{/�P$$�DB��I�U )r���D��&M!U麇���x�v�4�۱��ȋ"�L6��a��Z�l;2�r؉m�o~��M�9w'�j�4�}���PA��3�C��Q[y345f��B��#�M2���O�����qe���oW@8������h��Z��X�
��@5%�a|XB�"r�#13ʸ��I�kkWv%4:#$��~���H��u��lػ���I�3�@l���Y[BRd��x�H=�\O��Q��p�k�������g��
	F@�t,&̮�w?�#h���̇�����c~��V2O��?�1����
��A���a}0$d
�|-��ri��a���a�R��iъ&*#�&�U��h4���DtEm~}~%mKe��ި�7i5֥y&�iKN�d� ��0=C�F`���+��B��`F'���R��AwkW���.���Y2�lHْN�P�AS��a,�a1J@��x�l��AQAh��rV�3/(��Ph�=@_Fr�������Bշ*��\�D |}{x�a����BH�(<dLe�M]��б�r�� D�,�fQ�R*E�	c�#F!T�M	�S���������ipL����9�Ұ���+Gʎ�����%�&%ZC�!rٖ�R�<-�Җ�2�ˤE�%��V��;H��C@��~b��Ď�3��)�ߣS7}��\����c�����bn�zC�kYY�r��Ҷt�r�AgBL9��j$
!���
�DX���_��2U/iߖ�%�k2���ua��~1��?t޵�X9/��!�,�题�ʕ-�[g01M�����@C�ͭ��J�'�2�a��{�?�!�9�x~$�����2�JT�����5��?b�Gdח�f�j�j[�׷��ƺ͙?7���D^�Y�e���}	�Ta���̍��������|�4V��:Yz2\A��h�\F�X�ŞBF�3��*D����T`z��J�p�V{�k�M���)���)e������'�l6�������e��az̧s�ř۳�K;<ڑ3� (�Iހ@�����ژ���9D�re�X�rz����->g�83�iA������gM�9Μ�*	��Cc��<��i��i�P=
irK��cM�T�r����ӏ����L-LvB���L��FM���D
4#��C�Q)�g��~$S���J�,�w�#h.U!}���B����s�-z\������,�Q���駟�����}ϗ��{�4!������>�Q�`�+1K�Ӄ�k��qrx�Eϗk�?8��>���-¼q0q�3����{:����M@������ `���6EȝH�1�#y847{�Yy��'ʂ+�i��c{`�~;� �����ME!��h�<�p�
�§%S�6p�Wb��`hbe����,$kAS7�v�+A�����Q�g͒"�0mXV����?9����-�Mj�b)�ɏ?�?����˯���a�׸/��@� y��YH�O ���5�$d���ck�̛ϗڿ����^LH�+[�I���(�t%̰��5����e����!�܈�b�Q����^� ���'G{@IC<�=��C�*Om�=�Y�HI������t]�6r讶KE��li(��z�qgǇ<[G}\nGc�AO4JS���
���4�&A�v»��m��K(�L)��R�2U�|%-6�@��#�`V����]�O�n	!��=񑊝BT�����K"
�xx
�(T�����dj8�Г����#�4�Y�Pg��	gu�N�ș�tn�n��-Eb1��^{c?��HU�~���]�d�Tjj!S����9KO�03���&�Pk���!M�צ���4U�Q�8� �������RNm��� 6*�?�C���`�W�׵��O�E_Co��	WK�0�ߵ�>�Ď���/�sr�h����fE��0V���2VZқ��`� ���%�Fe�mK5:��7����������ATy�����?�4?׽YG��g3���F57� CzL�fT,�EB*��e$Ȟ(�=$�PU���T�m:F	}{:_� ���J����������������/p�R�6��T#c�/��*�Z�@10���1<��ܻ��5�Zvú�i�&U��_�(4uR��]�A�J�9^�R��VH0i�Ek��Z�L3���l�|�uv��	s�fm�Q�L���1IsJ�'F,YH����"���KU�2,J;�B����O����gٵ��
3�j�6��������� ���
�ɷ�o�ɒ2���J \�q�Jjc8�Z3*
��!2��X��J<6��I�Hd�oQaQݹ#e�P�y`��ɩ��2��������'b����i�u����� ����o�}J�%�$]��}?��,t�r��^��.�]*V��GB*]W-@�n��Çf�n��H��4w��s0>�q�uw�m	�Q��u��vR`p�-��04T�"c߀��&�v���� ?� �F��P�ga�f�p�@�<��ѓ� 8z��׿���+��a;R��{�1�zOr����wt���g�kh?�7b��X�[�`hIA��d9�+��h��s��N�T2����lf]�;9�맪�aT��޼ze7��҃�`E�����V�g�,��=�!x�@$������^q�(͞�����~��ڮ��K�H�J~�)�@�r:��յ|?�}�6�hl��RU�''O��~aǧx�%��罽��U���9�m����d��'���ǹ��F��Q�� 3 �ku�dP���sUH0��e)<�0٘WBӷш��7���]0Q�f��]���l�k�F%�h<��f�vBw5"�'O�@� `��
��zq/�2�1{d�~���?Vj>C��}�޿yi�o_ڄ��ϴ��^C��Q	���嵽y{iǃ'�nKʕ�@�񘚐�^'�Q����BNF7U�e�2we�S��΃t
���S��)�Ks8��.K/�M*��̕h�H�mC���]�Ϗ�3���[@���(�%܆�K�����G�y�[����=��QǇF�q���W��b�]׏����Tz��:�\7�z�}2��m-�To6!��lH_���ޘzo@gc�'�F cg�;�����.\�u5R2%�l�Û�ݵV�b��Ɂ\4&�����@����c��R�+<S�ж!m|V�����z�}�c���y��-�.�F������Z �<9���={��@��ٯ��@�K��*��T�XH��Q������V�gYX������/n�v5�YT��E�yY�|<��~�)e���#r�m6ʬI"6�,�f_hp:Zȱʚ�&���S����_����CUC�!�{��[e�z}{���;R�֞���g={��+�����=��� �a�e@T��謢�C���3�ɮ��k@��ŲaGC
ҭ|,v=�AKq.s�4���'2YX��es��xD~�_/� �c0����}���g?��ͱ߾yc��Pa�ѷ��g��FB�L/�맶�N�
�`�w����������vtrZʥ�٦�F�r���؄��~��}&�U!�� m�jv���������YCiN�n�<�H��!4b�e�}���BՇ_�e�c����b ��H=�G�`i��՗���[��J�V�I�-���k玼Ǽv�If;#����>�9�n�q�1��*m�$�H�����Г� Q܎��;i:��LEg%�����̼&�vqBse�K�"��$ڊ�
����lI�f��|m��FL�MZC{D`�H'J)� c����Lň�������@X-q��MԒ`��o#a���pHO�6۶׆p���OaR�qmr3���d�����G�Y�@��1� �
[{���E�0�!��۳z�=��4��olu7��Ad{�0p"��;����{�� ��8k"
��I �:*�$�B;�Ya�s�0��qH��SoVů���~��[ �B��&�0'mp��gcMh�����ԝv9�i��ߵ�9�X��a�3����l�����H٫�\��dt��R��<[�u&ۭ+U~��zh�6x��>���CQ3�l9y�Ta��r%����2�v�����R���h�߼~��b"ٳ��Pf$@9����I�Ho�\X�e����~aLS�a��?�ܮ��O��aߖ���`�7Y%�'mx�;s'(3��m>>���E|��ʎ�w�yի�c�<Z�(�����Ib!���>d�~h���[Q!�R�2���^JoG�����e�ѓ�ܜ��/�=�2�CRJ��y�0,�"i:Z���E(H�|�*}�Y���5�ڳbL�e؅5��pf�;h1V�aCj%n|����L1������񉗣����L���t����ږ9-�W�1'D�J����[%"������Z�֊���JX�teӐ!�Z��ƎT8hr�.@`��-�V_��`�L�*
���|m؜fa¾~�Z~nX�: Dj�l_�&����}�䱄t�Id��t����>W�t��q�}ݏ��3Z�`���L�@hu�1i�22�����A�>]-t6�~��$���n{@W-��2�v0�����ao߼��k���S�,����nmxp���?:U��=^�2i/Nu�4��G0�:�88ꚩ�gك�M������Y��5jKg�����9�c����>%�9a��Bz=rb�3�N���ό��� ��c��)k=W	�OEs;���[V5�U�78�p�ɖ4��J��I�zC�F����[Z�֣<!������|}�re6�.UY��?Z̥m�_�:��Eʼ&o��
 ��������L���-S����4Hi�'��_��(՚}�7��6lE@�Q�R7;�Ȝ!pb6c�5:U�f�q�+Og�4O�8�|���c�H·�(��P�W��Hu ʨ�=XǢ�CJ+��>z�I2Q��B�)��@�6���;�|���Q�D��W�8��
�.������6���$,�aٶ��G�l�*���ӗi��8���c�L$T�b*g��z�����A��
��� ����(cڷ�U*@x@MFa�p(ɍ�UM�m�)�%�J��������Z_��f\{u>j;���ڬ�1�G#�TA��\^��	M��ݞ�i�m�H,�4u�/&���ܣQ���`V�ٜ��6�w�Zq��@����3
�	�#{�Pf
A"3�${��2�И�YLEp��B�n2�V�k{��=I�!%t�8	U�0[`zR��2�?rK[v������ �]گ~���U�WU�E�޿^��ȭ̃^�s>�x����S(I�Ӟ5�PX�~ !u{s'S��hԨm�Tv=W @�9��kz\6�h��U�\9�j������
��Ě��Ϟ�t5�m'�V@�w�K(?���	h�m�ua_����#kE@�t��>���+������� �gE�f�6 n�1眂�v8Wf
*�C�D�UC3-�DN_x��:>q�7�֠R��)D
���2V�:=,8>=-,��ct�Y!ޢ͋��x��(�4�qeu�*<;��T�`�W���dyv�t٪O�3y�y�����޾{8����!{y�=?�T��� z�X��6w�
����T#g�n�qi2�`./�$���:[1-��F��T|V�b=���o/l2ۀ�3��!��R�9�ؔ~�h�;�	�)(�ݦ��2�X$2��촻�/��q��;>:�k�B���O��x��m	v�g�ݾ���b�����m�zx�L�dg���{��o����:6���!����1|ɔqf��t�wcEv�aMCkb?��Z�>>�JХB���D��ɽ-_/T	Lb�s�QHi���j��Ş�l�D-)s�����^}��߲ϕ�ٓo�/~�sms�+�J�U���Ȓ�_��*���n[���J\��$�qH�]��'w@�3��
�>���h�)�4��#l���x��Bצ>/+<�[�0N��A��=��P��|1-<1-���`�̕lwy}a/�iA��t��Kb0 Q�?�@`U,(B�S/����C6B��A�L�&�As�e[y��+��mo�i�>��TO����C\G�^�,��|"�W�H�<�e��Q�ne���YZ��l%JIť��(�]`p�(T�ҁC��˹�ٔ�h�x/Pw��V���{i�C���{�7����7m_م�=e��|�oڭ��
`� �+�����5��&���}���L��{�6��L�����S/�e߆��Ja�Dٌ��PkiX���ym�|օ����3@vH��d����gz�珰���.�\�i1B�dSc9����BW�UҒ):���9{�0�`o���Y�Ԟ==����v?���������҈�_�v�ll�gBb�1���d>e�@������b�{,6-�`�0����9��7�uI;?��ۻ���-!2�y	ӄ�)���l5Ȝ��2��P�l��vxpbO�<���_��O��j�:��eH�c�]�U���լ� �+/�y(4͊m�3��g�8����J��JE�e�+��Q3M1��JV˩��_A0�a�Oռ%�i�H=	��&+hwV��Y��*l����Յ����@�}�x���aa�w�Ժ�,F���&�Ө/�$�d�ƀ��l��؈�'T���Ҫ���&#2�Aӻ�o�nU��苤�GB�;!R)*R~���D�GU=� 	'us�D�S�5>/#�5���_$� � \�%���oFA@)5�1o���2�B�w��`�\]�!C�}�Tt=}D{3f8�1���|�Pӗ�2��:V3���%�C��E+Yh�f6�#(���˨��۷0����@���Tc����SXEE��0��R�I�j*a�Tv_�&�,g��S\�Ц	skϞ<�(����3�jS	p+�C$:�u:Y�v����#U���nΑ�^�xm/_��`<9=��j�ն�>{b����!~?>:�?��e������J�xL�cv���DgC�%MϸtԔ�"/��`�������Y�BFh��қPS�?�;�O"�����奍afQ�3��e"������r0n�.!h! !��~:���@@ά��'?�c��/~�Rj�#�R��\���VgO
f
�\�� ��Wjx�,}�$<Y/U����g�|�A�if�HP�M��d�"&�8k`��4�e�-a�%��c���O��WWr$�tam�@mwc�' �z%�5ؽ/��^�%�_�LDG�p������C��|7GG�8sUكN5lK�5�ܠ�N��纹��|����k2�zÊ����s4�`u켮��#Q�X��l>�|0�}	.��>3�䬥T�$RhΜxzn�����B��V�?���Rڽ��:Ҿ-�d��+1ʋ��2�@��|��%��6V˵	͙A�#t�6;"p�Z�aBK�>V�{����:��l��3TGbO'@��)�/l�,B�����9X���Y3_�>{E��>�E^q����99|jg��T`�$�n��.n�o�a�݊Ih��8j,�a�l*T�Tl�Ϋ�K���6c_��%�@_�)<y�	������������s{w��2�'sK�(���@��`ː4΅!k6����'��/�͟�//n�C(;��G��O4Wx��ޮ6��7Ú��^w��{|j\ 	@���e��5�5�$YTH��{{{'�����B��?U���W�^��V�?�(BE�d���R9FjԄ��U%L��~2#kt�YV�-�Q�Ʃ<*I
�#��(��K�`�����e�?yd��[����
�v����}?����l�����!����D�Ƴ$�U�6�Y�9���Hӕ	u�jg�=�.XH�j��T3n�Nf�M�|h-$%�U�<T�Ԩ���L�+�޼Wg�P9���;�?�=��,�f���MqHs��~�9���N�z��7ꩽ����;0�_�!ݚ�A�A�iR��1�8ڙK�.�`c��O�&GG�[���>1J�iH�%xb�R�������e�P�Y)uس6��#���X�dM�ӧ������?�hy�_��$��aM��K*Ai��e�[� �V �=��<
E֩t;� �fN=���'2#�`j� ,�l�����
��-�B�N"�5���u]����5G:���Y���mA����5������)d�?��f���4�;[*�e+�@���Ħ�������w������K �od���-=���}5<_jk�9�[.�y|�X���J����Ȟ�X��	�V�2�1!c���J$ۇV/_����u�&�PoV)�m�{`�k�E��j
N��f!�*�x1����AJ<'c�޵J�*t=���M2iz)Q�CڊU��}����>��|���я��?����_�����}��o���)P*���B��B�D���觀��t�U
�ӷ��\���#�ܬ`R���(Hb�^�"y놷��	���1Lأ���$��x����
���J(Mm.�De�o\��D"u�`w�b�`�(K5LA�w��k( ���!a:�+���ê�-4_�r[����&e�3��gl]�e2ܳg�a�?���sQh�d�2�Y=���e^�Qwg�6T�Rmn����s�ӯ5+�Q���>̍S���������J��0XS��l��������*t�bS\vN�BR�ltk�3@�|*�5��|oo߾���B)�P��;	��$�hH���B>��2� ���Z#>�1��j�'-c���:){���߆���l����~U��g��)'��
O=���;]h�'rx���~~�wG�٩�f1���,�KE�I|�''r乵;�))(�"`<h��t0Z�Q�6Ϟ=�����+'
��#�,j���4�P1��C�/a�z�m��Ȓ������@�E���"��8
\ sl��*W*�)�t��ȼ��?�oTF�F�����Wv��wS����p��1)�kY�ޯ6��4��͡5z�v4lE�I��+	��<��mÌຖE��3GyE��9������U6�N|�}il��dE:a���u>�_��ס㏢3��O�U�y�PV�&�'J�C��Q{����<p�� 	����*��ʄ귔�Ϥbߋ�'��߅z�=��)�e6��e��Q)�>c�Y�Y�c#
1.5|3h%
���2��g0+h�Ӕ��_� �}�����B�gO������_	���F1��|�H1*����N��<��;a���º�=��N�k�2ӎI������f���9�p�*?B���m��-�L-�˕�+���/ށ]_�P�=���-L��\}ZY����0�Q22�냘��n䋢 ��g�)� ��`��?�o��
+�`BG�v0?�^���b�xY9�#�z3@�6ܿę�L=�k*���7��<��,8R���V{;���'��̶�ѝP,2c��D�e�C�ʛ�K��
6Xb
�B�s��P�u����4�K#_��<�V;������m�NAK�^sn[��Ǉ8k��o.���Vy-&&�奇d�D��bIx=R?�����nw�>"e*7��<5]�$"z
k��`=��$M�"��&���[��@~!R��J�Ff���Ь
hz����V��ԇ�} T��%���ޚ�w�O�"8��=N��N	�E,\K��2Q����,�R�W:0��n�<�[۲����0�1n+���L��$��]ãT��P�Y��6�LrsK��2q�Vٳ�N�Y.B�����,s� �aQٛ�����I	-�؞<{&m��~�+	:�E�#v[s����э��X��[�`�+v	��?R��b%_��B����B�����^`���@k���.ʳYv��i������u��	�&k��5�sZA������j��
�蕯�9�L�7ou��]4O��Hl��S�b�(8c��x6���>fDs�9n�g��z*IA�"2����KEM�DFj��r#cs�|��ׯ_j��O~�#�=�}�t���Wxj�\�^f�ά}4P4�3�^ҬF>�BJj���&L�<̵���T�����q�*U��*|��~�g"�8���٬z��]^\(���O����Xh�K�^�$P 3�)�fӉ� `�wK��h*M��ʒ���MC;�+��(����,v��^�[�k��E�
l}&��W;�h��XUc[�lA[�����Y���'�S�SI/��/�	;�o��D.�ŗq�+���z�>$Q��.�?(�+CH��0�Jue��/
o�Hoz�M/Sg'14{�2i,jf�]��	���ݹ�b�K�
i���fi�'C��In�0�NS��
��$`��*��S{-���/�c�<�@u-��:&9��恂�5(�WoCs��B�d�BF��}\�@���f"
�U3�k@VIօ �؞X'���E��.^y�<F28l��J��k��2�wb��Jn��i�P i�Y�����a�L�T����5`�����ש��"�&��qh�����Y���2���(��^x�̃a3nV�2�a��1Θ����eh������`�\��X��ђ/��M:��n�l����q?�(SD+g.kh��Â>*�	�Ęlv��(��qJ!�*�^Ǻ</ $6	�����W��+%�)���X�7o�h�{�@�����r�!;>ܷ?����ր~<��%<�!$���10�ܕ\��W���{�F&kb�0���0�����&��>��~:VY±���{��n�sY��U�nP���B���#��y�W1�yq�Q�5؏I�	�Y~�!��
�I�2�~� ,�X��<KM��� 	�DɪE"6Q����Ag1����e߆b��j1��YQ��2C���d:�a��R-m	AD⸾�Pa.�F;�5�l�i��<���nw}!"~�����z���P��B�� 7�ƚd�w��j�0;�?����6^_^JS\��z�&��T�aD�f����Q�Ȃy���]�iv��tS���Y\��|��=��}��\
:��/n��Q�ڠ�gw7�#���O}��r%���z���&��Ԧ�Œ�ϧ��@//�"���̮��]�%�^�N���DudjFb�{]�}���7���!i��~T�CYT*�cs!��v���|�yf��`���;�b%9���Pж�O��5���fl]�2 ��3�J7����y���X!���sܯ����˽�����c�a\Ȕ�ҡ aǸg���珬������"����TcQ%��^Q��r^�b�vF�Wc*(?&J�|
��|��;����~>�9��p��/�ǳ9\�n7nҧՉ�w��_�����[t��E7q�J��r1d��V)d�>�[�Ӡ���>,�]�#8�@U'<s�Xλ�f�+�pg��Z٣[H�u�Z��i�Q��%�E�\�C��If��a+���-4�po=�&@Qx2W�Iдg�	��U���*�/� �����N�:gx?C����/�F�U��a���ݱ��Ȱ�'g�ɳ'J���U�EQ�NVn2O@��`<fY�҄ax������0a�Tm������[tI�1������y��>�i���4ϙ�����)��PĮo���`0��T�TUvY�tT0�C�\!ɷ�h�Zo�C��/��Y���
&�+�;���F�T^�^��A&ޱ�#�}&Yh����4G����4�d4�>�U0}��o�� �3Җ��Y3�pS�B����×�
����&�`j�W�h^��߅��'�����&��-�,��=�|�j�i���zfW��z���ę�mK�ͯpn��	Nt��&s��u6K��DU���"��{�MR� Kϖ�B��L󆐻z�ԂD�"ME���&[�~��%����҆��B��<����>��sU�&��$���-2��IY��S6Y�y ������)���͔v:p��v��f���\�8���d�f$#m�޺��<Ӕ���.�J���`n2�gOu?z��X+����,���C��o�f��@�̴�ڑ���n�X�A�*��/�P��w�dc�e -��r�Ki+�A$�Ю󛑄$�����Nd
ƻ���.zd1�J$��A���k�9�i��/���	��a�D�KG�h���ɯL�ʋ'���R"��>�E$�uPX{?\7W�
e��$�;���`+x
D�*܍$��J�n�U����*El�{=h�=�������4��ڍ���a��f�(T8�apϘ>NS���T�a*%E��1�̿��UoYs��ْ�A�E��9:��]N����e����f�����X�1���O��O���ŗ_��s(ʦm��f-ۅ�\����5�U�j(��|�:����44��Li��"ݥѫB̭Vp��T�D$�e�*��̙�M����B�vʱP ���x�D~+c�nZ�c�S�r'��IT>_��D��n��W�z�W]GIbA�$av&���8[}WCX�ғ��L˥/$�`��fɓ������I�+��ܤXY��2S�-�Q��q;�T,���щ��Ԇ�v���l!�ﵮ��}90�d��6��	E�A���5U���GbqR��˵7�.UT�r���&&\��M��	��O�N�ɳG��w���2��kil���p=6-�7m��ݭm�.�U杺_$��Ԝ2�u��hΜ+;��'���.o`��fj�D/���c:��F�p�e��B'74��兽~��T~�h��O��7f��|[��F�1�H�S�V�4C�����P;���X3��L5�fx��?���z��_��/�W?�����n�SIAзq�W/�Vѣ��G(�)�`��d��T~@f�ĥC����9q^����g��A?�i�#U��ʦLS>C��#&�A��j#�h⺃�P��w�;��[�$]��1̙= ���"<O�r�BS��X&M�-�!��v�4�D�v��o
r	s��O�X�,�|�9�eh�r���R'4#��%Be�P�TܥT�j�ժv���̙��5��a`������dd�P�x�����*��H�qȬ��o"���'SzKB��k�h�C��It<��	{����slL]�G�ys4����5o������l���-����x��&��x���	�R"�5P�L�k��r�д�"*ᬗGϟ� 6����V�ثoc��K9�<���""��㏭���O)���fМ�&�񞯾y�rx��o�_XoO���Ǐ���#9�.�߫�����؃����w7��jb~����|v
[�O�Y��T�*�9eD������9i�,+u�!$��}�EH>N��\�Aಂ���Fa��ѩ�[�o�g4��s�v���Fd���Ŏt�zį��O+<G�3��4mB��n�Ī��0�������ŵ��oj�����}�A"�jb�Bk+)S������d��M��l�~�&±�bU9]�ģp�G{��U�Ek��l>ݳ��F��T=f�q�{~���շ�p�����XC�( �aa̓��~ֶ/��3;ythó{q�3~�KW���:��92h%�D�>�+
Bų�)5p�N���A_R:��L�o1l=� CeJ�W���j�)	�HT�S�Vut5��>�3Q,�XW��^�nF^ԣ~ �g�ճ?����3<��yT���z!�&����O�]>��T���D�*���sOg%�6�l�V吧/����/�F�����}���٣G�3��Z�Y�ݖ
�F�+31�*�[ǔ��L����xƞ��0�0������(]01'����|M9�SOy!����&G��V��C�U(�J��B�S���v�Z-����k|��GO?�O>��}��l�8Ӷ��z�J��8�F�Y%��x��f�F�>R�z�̝oq�"CNY;������vs�9.�N;�ai5�Y����պ�F�g�������=}|�F=��Lզ�v*��X�uc�ν�}�_�zz� ��=�����TsUZ�*��2m�Ǐ��t]�v����W��`j�q��r�-Ǽ6H�nvg���SP(9�W>,����ԯR�����n<يm��nOt����+�Xְf�
B�cLK*��s3T�j�ڬ^���S�i1���m���&��!�t�2߄󎆽�u�/�w,[>d�
���^=�fE��QȪ5@셦�e4}�����(G�����և��TB�5
�(M�]^�b�X��25E޼���U�Q4�zU!�!5���k`��ZWi����r���~/O�51��R�ע�.��E��9z���D�k9�����Ql���ퟩ��i[ϐe�9����\Ia#j�dzro�ío��b��������>z跐Л9�z�iT��,�X^l�1O@�M����܉��Q�%���v۞��ս;:ush����l2a�>���=���)��1������3L�D/�d��m�)K��:��_�A"f���	;�5�&����_��/�
y�sE�N���C����ӧr�uC�חb<����o�ݎ�= ���L�D�z��)Y�������o���Y> �x7*�����lzo��W
�z�w(�C	�c�����K	�V�g{D�tzo���2�e1=pNM�#U<{�H���LTTV�xFm��qp��k�m���:WS u�Z/5-ke�w�g�6�{@�,}t|��J�3��G�T���[T���/�C�Iv��"���d��ʄB?⮇*�O��wB�k�j~N�b���T�&�*hu��)��#IuT�j�]������Ј�d҇��[zw)
�"�kN.!_��áh�M	dV���z����3c�O�j"o�[痔!�)��*ԁ"�a��t]��8vS������J�nc@�c���������f3J��M�KM۬�*��*��S���2&�lp��8������'w�q�&�MTN�y�rL�a�f&���v�M	\�Q�ֈa��o�'r��?6�����땴�>���Ǟ?�ru=V8�]ю�*��B'4�$�OdS�5 ��p��ta㻱��b���g�ӟ�t��@t�����y�ZwfSx�<���@���c�����/�R��������xY<������Sb����$��/�5؋����o^���K+7�"%��h�(�������k �;�?<ճ����eA[��*��yD\����4Ֆ����?�8�UƪS�l���28� r�lj/^}c�7�Rj���ʔ��nj��R/Գ�g��g?�珟X�ݱ�~�Ҧ��|d�A݌�qo�!T�a�8�U6��@~H}IUwEcç�"�A�����?�;�`�^*۷��q�k���A�/����OVKw��x�����C~���+��;C�a0Y���Ar�j���յ��Ը^,0v%a|���2�9ޒ�祺���CG;�R׶�!4\/P�?WA�k5C)�����oՕ���3jp��ʻ`�;���˅�3�~���J�la��E�µԘ�;��������x
tp�ۭB�M�����[Ԫ�q�l�T�n���7�h?��Z�@R���ςH�0�Q F-H���o���S5&�88���c���rrz�u@l:]q �R��E��Y'~�ͷ6�L`4���v~m� �� خ���f�u6}e�n�&�_}�&g.s?�<��7��������{��T��s��D6,U�����x�r1�ٱ��U^iʒ�mޔ���j��e0T[K/�먧�?}��^}��������Z(bj<a��B�YD)L�V��
	���� ��O#g�?��a&%��]�`>�4������!���JJ��F�|rcK(��x��̎��4����G�����ݷ?�7��u�OT&�{QNd>�{�P�B�s�#U&�J8�kL|lk���);!bB�U]�Z�f�Z�T.���:Q+R'��J(���*�5s����|$x�����v�#$�H{ƛ&�U}�uZ9"!'��:�Y�p(�A���@/�����+Ȳ�������Ko*�T�<��	6���F��QĴ�З�����W�P̄"3���t�iM���M6�$<|�
U(_���>�7�^��9��,T�l�#���̽����k�8<a��%a=e@��0&�C.�9#<�h��AY1��@ܮ$��VHd����u�>��z�7'j�X�CBܪ�S5�`�)��|�zP?+8]���U�� ;����O�!BGV4�Xֿ�x�Ŧ0�[�%�z����&=�^/ ����iFd�1���C5�ĺQ�/�,�׵�ݠ�RG�7;;��/�:[�E^ aH�'V������Y_�`Hp��"A\`Moջ�D
d�
��A�T4^��8����I��16�:B��KK���5��78�-�p��u.D��. �M�P��9E��6������j�T�;vo�,��-���y���07�W�XG"58�8�P��ha��v� L�~qzκ���Y@,�L�Z�Ԍ5��9�#��%@�Q-½��F�2?7ǜ6$��[m��3��ڻ�um�#�[���.�@oפEр	~�M��K!�:���aP��?���x؄/9s�9�D��@�Eӈ��/���3l�S�
{4��E�;Yh�$��ǧ8���hn$É � �uH���%VfD;4um���vH��ǈ�&GC+��b�#��
����$uއ7$���@������,���;	�b� Ac�z:5e|k�d�¼NxM��s�g���p#K�*2!����a���=�����j�V.C� #=���7Vԛ  ��M�>� ��Ձ#5GA]=�t=�0n��0Q]��H��ic X�����$AҶCO
�)z��������M���f��]��Ģ�A3��f�X�,ͮ��Z�`��n����zM`L����C'���[Xe��Yo	��~�9���U&�!�mzU��r�h�8^t%\TB&�)Z������{��{��0^t��b�Fc��~\�RE.\�*�����j��D����hS� ]��8#�O8�����8�"����:�������.e� *.X��
ɥ���(�&�y��ճw�>�D�,]([���@>!0��^����K���U���];1� �Q���3���� f���=���v�\�����:X�w��<����8�	��A�D�r����]#�Ҙln�px��6�1;|���-0z@$����q@$\��DJ�"�VYOͦ��e�  6;��� 3	��J r�z%�����JtbD΁s��ҳ�BT�}<�'o���HV(���AA��Id��Z�X!�x&��N���z��LVl4�<aŨ���t�t�nm#��F3%@)kM���i�"YL�+��k���F'{M���4VVY�ʗ՛�G T/���#�тf!"�e��-uu�I���T��[اDCGC�FK��
N��w l��Cj˒�V�G�tS��[��u��.�ui�)�D��z���U= ��3VV�-�F��	��$�Ǣ�C�C�);�Փj �%sS5��mn���?2Hz���ɑ���Ao`�H�ɕ�'j���l/����_���,�m�<W���������2ѐ�@"�o�o���7�P�1o,���7���#�0'��f5.�� rީoуix:	Сbj� �B���1�M@�NM �5��a�Y�����uy��Gr������[1���nf�uU��������S-��N�Z������ۼ��!k�;�����h��F�r�+�!��e�6vP�^ �#�V�I#s�=)��	�'*��̢X"&$�d����ӐL�L�TjXd���)ˏA�m`�0m�� � ��MA�\�q0�$M���$K�JMl�+�v(��� ����yz̹��6��턱�����2���
��TO�N��v@�ke\X`��8��Ɩ4!��7򠞎Ɇ��נ�۶���m �
=lv ������iâT^���
02��4��Q��N�������5=Ԝ}�d��<��#J��B����0=���lU�w�<J���4V���R,Z�J�ۚ��Z-=���«�@�\�N��b�$Go���X�4�����֖����R��b�X�p�c�0�MMA���X�!��+��p4�ܒ��������:9X@Y����:�M4����B@z��ߥ2���z����B��>WT�k���p(���5����"�s�bX 8lt���:�^�֛D�B����޾T_S��+rmqU���e��D��^� -��	x�*��7�*D}V@J���j]��dJN�E$�,���f�wΏ�	zO!��Ǜ�a�>0� 6D�`5�O�c���Z��H5*"�d��rKu��Mmk
dqLWtf�"k[u=�<�q"�?�Q{Jh�p�ɭڤ^�QZC\�0o��1N��p&��\Ȱ��?��%W]����s��M�|T���!\��6�)���%[���d��{�����.���>b�̪���4AR	Ş�i�sm��4�E�'��Zc�/�g�5�F��K��LO�)�+����'�4���7�mĮt�d��!;D�]� �����ˣ�,��� Y�.H2�1�E2�Dl�X7���'��&�Xy��l�B�$_`ٓ!�zb��kR�qAZ?F�
-}IOxz����&!0=h�m��/D��^%��4�B��#��%��<��eP������ֽ��.W�����а����IC��ٽ��Q��[���9$F�4��W�P�E�=�u��C�+`���РlIJt$����q��*��}T���4�Ǝ�(H��-Y��r���r��t��6%��z2�rE���i�wZ�Ht!�]�z�H�SF%�F��/xj��ivf!�X�r�x�sL�F<�;H��<�A��`$V�5f?�>�1V;p"�?%G������0r�l�����nerr�h��7�� ܝ��6uEp:@/��VRo-<7ɼ�YM��Nh\s���¼���!�9O;t�����I���n��a�W'����ܚ�&1�h�qL\�Y��X��d�P����
YQ$�����K#�)S1�yM-�N��M�wvV�YP�._�(+�+�6����~�h�J*��Hx6��us@��Jxu�`�� �� B3bO�zO3!	��ƍ�P��k�<�o�\e���d�1B/�� ��2�c�ռ��]ڱ�g;圔u�!?bյ��~g߹���v; .���ܴ飨��D]�H���J}�8e�m�
K�z�� ����v{b7�{Ya�h+@o<]�B���p�_�n���RS�h���Bm�cA����Z�}�/��!Jj�j�\������Atl�j�Iɑ +�a��S�a� o�l���yBZr8�r$Im*���b�Q��>Q�2�0��@IF��T�5���?�3Od��M gbT�� ʎ-ۃ�-��ɂ�#��dSwv�Q�7�a̭�NOD\[L`Mw�BH�@�[݁��u!	i;=�:p�`[�S5���%Z�n��6�=/T��oH��te�,8������k�s�_���wf��1��s�"g=b? ����*�.ue�Zbh��z��Hz�t�I�ۀ	T�7>���m<��aB�:95!�s3�<�=߻wC�˵��z�肄 ���P�I��P�]�$�������`��z2@��UW�b���N$��U������Ⱦ�0Zf�	���o�Ȫz"@�rS���l�/��72�XrDưI��8b��\��Ce��O�p<�'�r��n���< ��T�@w"�%+V��c�����bǸs),�%���z��B$�iDt�ɸ_`"��0ȗ9�:�8>���`�+�:�����U��n����/�ۂ�R@z�Dz�dޏۛ���<1QҰ��F�.�mj����p5e��R1��3:��vа��ajZI�� 'j�j��=���`�E���:��;3.������@Ų��� fC�`�S3��7���v��>�;V<0��EO�"V��fΨ,�� �Z������I�n��pẍdF�4j�
��V$�0��r��hQZ/b��'qڻH�"����rZ/�6e�q�գ�Z��2������q��no�8¤d�����w�*k`8W�
ҝ>a�։��$�6�s9�F ��w5��)�V�2��������a|B��ع1�(�b��!i{��1���=]�x�|�qC�{�����*�58�/�лAEr�7@B�������T�� �hu�@j���&f#-��0ms\�<�1�a�o,�Mݰ]w��͇�0]b��tQ����J�ȋ���̢�7��E_'�m�|�@�|~@C���������gU)��H���y���|��Z�������%y#B�"spE�J%g͝���)h�N�G�CV�����K	,,��)���⯕J��4�m`M",M;�D9"�������JڙPoe U� ��J�#��i���U���Pt�U'�u�m6�1 �I���	�[*���z׸��|�$s���ecM=���Ьr���g�xHf�,9ț�y���j\����a5�{�d�h�z��a�X6�~M�:��v���yÌ�fD���|"4"�w`��+�"�ނ�83�� 	��0�&Ȑ��6�S����mO��N|�c4�/����$�NU
8@EԴ�X]���� �)3;*g ð�?��c�жeuc]7}M����iN�?,M���{i4a����S���EN%9�I)3q��X`�֌q���`-� �&G&~f�����D��غ�a�ѽ	!k�����継1MY�aW*���<CPD^m���m����"4l�62�j�Z�*�m��e�m	�RVjx��&�:�N,L��\�+� �X ���	y� o�l�"�@`��P%9T��B�4P�£S &6�+����|����Ѯ���^y���HՈ�l�Ĥ'I�8fy���T��Z�H5@4�!d Ӻ�oD.	pA3��㠴�D6xD�)���	bB;��A�lFC&Y���ζAm���St���Ր��^��3��'�`��d~շ�Ua�	��֊�&�?9�[)���� ���=�/ru�x#⋰�G����W2ٻn�t�{f���?�QYR��7r��獡(dU!���� �u�K�V��7��bg��S֦�O�9u�L����+1	�tT��d�GD���/��������/`�kØ���8=���B�1B*c�K�#�/ 8��Nf;A�0O�0��_y��Y��hC�u�Ќ�x2�E��X��r=�#��(� �2���(#��Q�4ei�ۥ04��*te{�tqK�{�q#�&t�M ���갗0w��p:���m}NΠԩ�L��Cǀ'e`Ֆ�)`f���~]�9�X���Y��4iΰ)0��ẃ�h,�$z
	*��w�4�Y�Ȅr�X	��W11Xw�:de��ķ�d�pX8fiz�OMN�ߦ���/>-�w��Q��6>G\6Z1��&=JU��f��`����]!�a@9Ğk��y�=,�Z� �ޗ8�Z����"�g��G��e��Ę�V�����A���8��2=&S��[�T����[���KZFD;��@_EI�]�Ў)��_��|j�S�xva8���|v2d����QLMh
"�0V��x����1pǄ���� u��[��F<�f��t0�1D8d �Nb�%%�dga���<�@X��s��W��M��Xx��1���		]KO �L�X���q��ȋ��)KC�$��V1��v�=% \f�$3Y�tV21���
�ݖIG8y	vp�.e�*u�<���|����H(�U�4���1���eI��Yұ
��6yv�&NG�?��A�R�H�L��\Ț>,3�[�K
<A�{��tOpR ��3b�ĐL�����l��2��D��E����<bM`�өI�b<H@��7��FN����@�4�g®بd���S@r��#W��Ÿ/b&?��10��~�N7����:��2�d���i���9~`�ǽ�������R�MKV3?��N	�8�q�h҈jV���8J�lǁ�&:#��QP� �7�U��]ݷr0�s�B#T?�������։U�&���4���Zv��;�Emhŀg׾�g�]�tNޒ�:��<1��.���XX2���%Y^��+�aݦ,�vHG�į��֑���/>,J�Tn`�E�/�����KN�8m�(p�.����e4-�Q�����Y(�$س�I�/:~V1Q+X=���i�B� �q��e�����JL��#�?i�z��ݡh,��Y�KwlMv��3uC��u���Ra�^8�@P��$���C T� ��D�J��ml3�EN�(C�I�q:Ƞ���A#	غ'�ƥ��H�|���8�;8�Dεb�h	� ����r+e�{Ag�c%��T��ds$��ш�)��m��}@����{,pt��*BC�B��v���t�g��>Jl)��ꁾc�B�{Ln������?ajkj{{�&�B��Q����M-��R�
Kz�������V-V���&W:0��<`�xqHy��)
��:g;(P�8��znn�)��d
�w&O!��o��8���)S�rej�rc�!eS��ś��"M�1+U�t"m6�	yH���ŚBy�0H���n��$��|cU�DD�=��q����>Lr��4�ĵ��+��.�k&-g����������gd��x�ɛ->�S;��5%���`���*�7$��D���1��腪Cx9pݼ�!/�z
*�rp~RJQbݫ���[�ݠ�c{��У\	��C|QB�Z�X�o�QQ]���v�d�� Y��Bq�$7:�P�CR�۳S�6?�D��n2��_
�
=�� nuH1��������00P	Y�1+�(|\�<�ʌ=?Ţ��=5�� o�ѥ]�ߘp��E��P;�s�c�H�^��x�s�
ʤ��f����uV�����Zޭ�<p����BkGN�׳P�����J�:�S�0�QM��97X� gM`�CB>rqjt��8x)L�^^���U5xRH��u�=D��]�k�L )�GJ��s�`��ni(��]��Emʦ����V����C�}���]�#w�����������s|smS���R����z����j�De��p�VC�fK�G/���"���?�������+@��51�lh� ����;��]�l�ITҏ���D&�b����L&"�6W� .��M�œ"F̙xs;�0a��5���{�&\T85��
����WN�!jϤ��ҧ���!����b�ʕ��զe/�)jB�#��z"�k7ڬT�2��ܒ��'%>��z8q@L����qQ�ajBr�K����-Ag7'�5����~mIU�f_7C��T-Ju�H͎/\��e���۳���豀�������~�SlN��"��m=�Q�D0Nwp��m�� 2�ȯ�R���Bv8Ŀ���@��I��*ʙ.���x�&����ř�l�Q��I���dK5�`�+��+����l�6�f!��� �gH13� 1�z�Y����̀u��d�%OH!��E���C�TKH�I���Uz9X������Z�z�We�ch׷H,�Il���t��P��ytXø�Q��be��C#=5���i�3! [e�M�S!�D8 �A��ĵ#����ZO$���#��cs�B/�F�M��� @��2�X�'�k�Vg�c�&va(<w�B�d�~�A>gl��	b�%�c���ՖS�	,��\���Kh�l.��.��$�%��3�k�i���o�Ѩ�סS���2��r��5�6��p�씬�rס�2=Y�r~J�u}�]�N�}:�s��Չ[�x}SO����Pz2� ��|�$C�O'�����M_������E�5���JI=��W�B�)�6`�۲��Ɓ�U@��&*8�P�$\���zOńI9@���4U����������X�&�<��>yS^3�t�	�3�������5��6��0��(���?��,�1Ï���X0Y��u��X�.��ȍ��G1Bޞ���(]����7�yv �B�E	�0��Dֿ�)�8���$qL��[������Q"��я�l5t�:A�u�����o�E�7�jP��s�qce.��-����1aֹ�����8D�r 95ԕ�i `,s��`�7\�=�C�C���i��s����/�Z��eșXN��M�UbǷ���N��1�u���^p��^��p��*6l��o�,����ʑYp(�G�,W"t��X�S���M���D(��{����FF"k��)3��[�yVd&'���BI��A�Q�B��5�c6Y[ߢ�����
���Ƴk7de�.WW��9z���L�/�_�1L���ˍ��[�X����e� �� #��H���)��&����,��:��N��TS�}��)�q[[�!�o��ln����U@#�.�ѐ��\J����^X�4��W� b,?w(e�R�X:�䵪�L�Q`��7�^��~��8vI��Գ�f�ZaũC}'	�0	�'6=��i���lM�k�ĢQ�"�u�88a�I*E/2������>yG�P\gjH�W(��b���0��4�d5?���S�OY�j����\4F d1nOY��2t�J?+2�@�!|.i��ԍ��P��e��,"Eu��C"9r`I� =�+�ȁl��������eA�=V���r>��j�y�q���c��Ձ�A��!�GG_C�A��ji�Iw����2A'����������|$^�����b����|�dX%{�����t��eݭ�gT�0<h�&.����I����$-�i�쐯�Ğ'��tBς��yQꂆ*��Tcb+橇�I��z=�t[��-�$�Z��5lщ��'Flf��l_����\Y����?c�����u�E���-77u�k!),�m� ���B.'Fv��qU��^ߖ��	�q���	9V��wT@V�uB��,�wz�U����	c2��Ԭ�ݎ#b(`8A()�"·"tMZ��^�]G��@k5�B0��L2bS�\Y��gޗ���(�s�� ��Y�$%\�6x�/X�@����T��>��H��wL�9#�Pb*� &� �A�Pi�z�(A@��գ�<'�vC
�?�1rpnL��#a��۲���P1�)5T�]�+���VcpmiE64�D)k�:Q�'B�1yf,QO�.�y� �<�����Y����>�A����	���@-Q�fz�"�f���������h��˱�I���H76="���C��d���4h�w2���}*'�9&O<t��t6o.����,�n�Ko�/\����+=��H4(C�譏�^�����HdHǑ�C"3���a�f�;��ıň���dBS�1�
����1q�(��&�艈<d]\ӎ���|f��C�X���8��C��ʂ�T��Gܺ����IY7��T�Q�~��90w�{vZ�;���'U����i�:Q8���U}��4�T+��IԌ2Nl�c���J����
I�rk6�I�����F�e)�5�Lh ��]#�+��{_��"�-� ,	9"���� 1�$��e^Y�\���q9�\Lr�!�,q�v{�!�27[�yh��xJΩ�N�25r$q`=KH��\H�8��8H5�?C��r�0�0�rE���*#0�0����1��7GL��p��\�R���G���;LJ���*����xM��O���!�=n�@jz�\�~��	s�r��A�u�*n�G���MįH¤oI^�[�7-���Q��N�< ��(�c4g�pdaN�x�^y��t.Ճl���3g��,nl�O����ޙ��cH�ٔ_��\����5P�@�8�O���s\��!��f�+�{V�y�55b_�fM���{X��?�N�&H��M�f��s!� ��$��G�~&yu��� ��d��������%�2Pix�h���a;�t���p�2T�,���43&��u:�Cc^��H��L�)zj����J^]�=`W�o���BÛ���I
�'k�1nG�
4?�a
�J�z�������ZG>7�_Uݘ[�Izd��4m��V�7SCz���0��C��:���$�9� �QO�S!��x`1+���	8 �G� CBcM%m�_B%����ӳs��_y��um�,�鸲і�����w���>�n��.\P�3wӃa�c[�}I������AnCI^�q|�ѐ�)�aʒ2�� J�������)��#�J�e�
�L�x)'%��G����c��{�,�pGNH?-�{�ˌ�fiyY���e�Rd+C
j��Y�|@c	H{�gLz��q���1HM���D[	:��9P���գ��?/O>p�L��B�V�óO�����N(?~��$.���LO�S���|�$�`{�Mi�͢/s���W>'�߽_^}�Y�˟Ȕ��]��i�� үvK�V�Ը��~DC�]W!?|�M饨�H�IDR�಑G`n7+qG�c�
V��������gX�@-�r$�`{���[q���ƶ���v	3n�O\�ǡ�� K�K��+Q��%���Y���I���c��3���K�ݮ�u�H.S������<r��=xX�]�.�<}MÄ6{PB�25f��E��g�QC��a�����_����U�w��Ia|Z6�vۢ|�gbLO�����9y��㲵�*gϝ��k���Si]J�I6�-/������.t=!h���ي7��Ʃ��<N-��ЀI$W�M���	K=�{�CY(����-��:�.��Z[��9����g���NȽ�'��\��jD`�����#�%�5"#�&�44^���1�by,+�&.k�! U^j� ,I�L^�.	{7�3P�=E�$EB��a)�	w�*i��&>ׄ�c���e�A��(�3&m��vㆌ�D1OEz TC��9��66�h8C�$k()��*�Z���<E�@M�����X�Gￗ��W�.J]ߧ�/�����ɧdljA�j�Ѽ^'���5���`������R'[_��+�?t�ޛ�'�V�5��E��4恼�^�[�$��'_���{��W?����^�e=��a�(��Nw5C��mv���P��"��M3Y]�:��X���Ot�= W91I�ʓ�.�І�Ĩϣ�:2�e~�[�ݒ��p�'\e$V3�;�ЧW80���'� <!?Z�����Y]oIT����;�gF������O=-��]���y�ܒ�>&��u���'�����X���=;35)�7��@t�{�s5F3lN�V��=0;.�y�Y�ڳO����P"�+?xB�aS&ƪ��_�P��Fc ��n���5s�4z$% f=j�l�Xk;2���͛�� S����$g/H�Փ�����eIsK�n��kMu��Iiw�!�[u��G���@j|E&�X7rl��d!#�9��� k1]�C�Nw �.����Y(�p
��᥄���/�3'RÙnd��S��233KR�~s]=�H7����c��EK �#�T�7��AάT
(��G����&ee���2�KY.]�J=]l�� ���M�/B_R�t刎�ӏ<(����w��?M�{�C����~���y������ӯ��BRc��w�A9y�QYy�4zO��5�T��ڔ�Z�**?V�b����u���L����.=0�������z=���K�3/$�����N��0���S"�a��������;4����Qx�Y��Cz���(�Q��D����C�2�x��6.U$\s��"G�)Q<����!��;�!��Рd�\S�W��0?����̔~G����G/��u����rhv^�!t���8z1)'��|��_�������S��Lh|��/>+�����++����{˶�>AP�	}��=��|�KOHe|R~��{r��w�pT�T�Gz�����V%�M�ӗN�%<	�Y^9� �{8K F#,!�&=�Y���h�&��R.�w�5[�r�ے��{N놫h�%.?U`u��o�F�z�ߔ(njH��ؼ��%����
0}Gϯ�:�����
;�k�kDE�y$��S�`�K��K� n��H�tT�1I#�	m��Ճ,�rh�� n�3+]cm����Hi�!זVI�b������M {�M��bը&P�ʇ�z�&�T�+�!5��o�x�`���=k)����a���2ի��{��'�G�b|���g���܅uY���<X{�Y��H��rč@���e~nB~��_�+jٯ,.�g�I/e�S71����:�]Y�o�"¯�\�����| ����^=��z�>y���8�+�C �4��k<��큉��E�<c�1�ِ�BOJ8[f?g�3�brL�q2����[ɭd�1K]��x$� 3#N��8#m�B�0���nI� �E���K���1������:tP���/�k��'+�/��)21Q�B9/�/_��^9%�)������G�;�zN7Y.^�&����'y即���C���}C&������N��_�7	Ջ��[r��{��~NN���?�(��\�|�]��>�����[�8*���7��W�"��KSD$AO�n�& ��!|cGhݬ��'�����!0L׫�˄��r�7��l�"�evK��0>=��v��������4� ��-�	�{ͫ0�+qp�	ˣVQؿ��^�$q��vx�~�PGnt7�y����ʦF���c�����_j�Q���3-�Ǥ�����+:�oJX���iW������gv��! r�0�:�����5�vZӐ��r��jS�mv_��H,t���ISO��ׯ������P�4e�0PO�ח?�*W�ݐ��]B��q9seY������ɇ��k��ƬjLa�_}ΦZu$���>y橫����ҩ�K�� K��M��!o�!0Y���_�^�Fz||VC�9�gN.�]ah��jJR0��oħo��}������ײe����r���)��9`�H��T�5i2_��D"�s��)\������S?FgbdO��bxQ�,E�Af<ĹWl�P��	��{�Y֝���U������� �UR閭	g����n#Z��zj��i�vwI����LMΟ_���Y���;��z��RQƯ����U��Ɋ~��_�ߔ��?&[�ii<�A�vԗ������rS�9��,^[���>��k򷧮H�_���?����K�z��I
�.O ���=� �E�!/��ϐ`(t>�Q,_f(d֘���X6�u�$�G�Q�?��rN�ԭ?xp�<��g������ƙ�r�ܲl7�$�U�~����4�'^�4G����$.�;��߹�NCv��������I�nB�CV��Q�]Ө����U�@�~%����=��6]��1�[�dnnF�y�}����\�^���)�uA���	���͚���ࡽd�$-c�%-A��v&W�#�SgllLV/o����b�Y��
�27UaB:tdTA�$0��4��gw���x��	��@�4d��NI���i�<���<~ℼrp^N�u�Bc��H�����Ě����:΃��j�!I���T�x;�s&��&�a=j0,����4�^�����6߶�-:�)A�n�B���~3��"È�Ì��?r�f�1�e�+�:�8n�좝Gᘔ���__�q!�Hl�7:��,�K��,��
��aQ�:^�W�x[>�G}����S�O7�O<$�<��L�i�� �\�df�A�`օ��o�E�}�&5P�U���!���F^yu����v,��1�j��riL�=���?��M]�R�w\�}yY|���S]�Z�z1e	�P��� j��o^���<�]��;H���4�NO4f��ZD,��W,�8~5�N���S����V?���QrrZc�A�.�^[o,�3���@LJ��$'*'�c���؁`'UHnn�N�0%��R�t �u�LzѪ�χ4N�����`�(נ�	i
�?�$�tS,--�5>yRff�enzZ�,_��U�1@ȧƷކ�ML���l�}�D�8�m��g_ n��;���9��(���^$qQ9Rc[)�$.������˼�������ޠN���+=�^�ApR��;t���w�+Չ2�-H �/&tL��DUjഝ0��0A��+��kr��1.�N�x��>�H*�=3��v �hX.�|_��!�%q RFF��s�Vt�O%�=����d�:#�o��ghŕs|	(���t(���#u��`��mv#��-�?�Xĉ�Y_�zM�{�}��G丞��<�����)6{}���w#(�2x��vs[&ǫ��3�׮]����j@&ɻE�'��o���I�f���V֍��0�y=�]Z�ၤTm �ٮ�[61lCE ��� ��:s=��Ž|I-t|�����e�]�,0��H��̏�a��k���ٌzWQ��~$ �)R�"i��\��t�.�ŉ��ԩ����Z�����h
�Y+� ��aW�n�����PDsYd�A����ǔ�DB�/��0�:9�нџϞ�@���?��ȃ�##����-!��"c'>I�AH���}ӌ�S�*Y�-��.�G����O�X�A%�go4e�  ľ�ol1��FM5�U������ʦ4:���0��r �E5�ׯ\�!���OȾ�^9z�5,[��rS��R��X�'m�,{dZ  .d[�aM5�g/\�{�bX�^�B�q��0_�w}fkԸ�F��7���n][+�3��'t����Od��#tMNَF�Wj�UR<�pLb��gR���2>&�Ҫ�����@�A�7G�o}�9y�������8�-�<�A���)�O=��<��L6��'�z�`R"r$�قWq(�i�\TO�Agn]]�X�՝n�������}�Z�J��m;��r�i{طN�Y��9Q��G��>yħ˱ 8U�A�K�HÃ��y9{�4!I��y�������Iy��G����G�MH�S`@a�����+��8�,5C."���~�kҍ�s�tP��x���7K0R`�	����mܴ�S\x��]�rAf�U�	q�~�iy������~h("V�������g���ǌ��ń�q���IRfP1�?��N�~���Imf�C��7���o�����X^^�?����W������6���ŗ�T����y)V���4�v0����T*vZ�!�B��[��6^#����b�0��w�������$7B����U2����p���)BqH�]�oD�ih��@�R��*��({��Q�58���gڗ��}������2��/�.ȯ|�Y��_~_.^�,c%(�������Hvc=�+�����}��K��$����ȩ�����r���l`[��lo�ʖ~�MI�4_"c6v�p5⡜�R�ӳi��\�Tj�BðE|L)�gD?�CQ�D�b�+��>�����օ���oʥ�mY����Ԑ���'�"����(���i�E�@}��z�D�aAz?���Ў?C��%��^�U�����tb��oh%A��s+�����ىqj<x@��;ߒ��bZ��<������{�܍_�]���	�����Sn���s����:Ф͉A�=�r@`Y�xlX��\U+d�ɉ���q��+ծ��gj��}�L��c:rLz͞������Ze��)��ln7��?Yf����p�Vr�J )ӾgI�͌�i9@�������}������#gH��U���}��_xX樧��}���`D2��P�F�Q�4"����Ɛ�ut6bH�ݳ���[�����VYrfh8F�͍��&��D�j���0� ��3��g!�k����L��ͭ�ll����Y߫�l����]���AT��o%�Ē�z����- �)��&�4�)	�e��ҭF':<���Z�l�q�a�����0);~�0u�k�&ґVo\�X��f�b���*�\�};�+]�je�S`�o�ޖ7o��b*]:/+��dqK�;5eT��=�ks��%Zm������`Ho9p��lo�`����@�l�4.�E���m�1�P���9���Q���#GeϡB�r�25Q�{�>,��A��sd/��Ylվ�����1g�J|�[x�M!ID"o�$%�%�p�+5�p�r���r߱y�B�H����?�����,��o˃'�������dz�Ei�78�h�k4������r���2��9�W�����g6L⤢!(���y�������0}BC�2u�����NW(��U��|�����-xԏ�H�3����λC�{�=);�H9-O�i��6�[�Hj�͝/<!�?�Z�Ѣ���!���	c�����QBl���"��1ft�hh21^�5& 2��s���2�s����e�� �caa������ 5�+w�kRp�J=��GO�@�L`�QU��Z!8�����"H���p�I�9=���g.�=/t\�n�������	�_�4�ٞo ? �Z����ܪ�Rq��!I~V��K��| �WW��Y׵��|��u�|Yr\�@�0a��)�	���<%T@k�bw���$]L�h_���=�5I�u����	Q��G�2��92{M�7FO�^k[�b�&y��D���k&f�}�qt5���rwX��C>�t�C�g����3g�����gj���l�<%�V��~ɟ�M�����<�����/�B�\�F��k���x��Քz7�w?�X���oƥ���a\@�:pt���b#eq7�K�ے���t�z��7u��)�R.E�fi�;>v�M��0��N�:o\����@�sZ_��'q_S����B���}��<�sb�O#�\L�5��3BP��r�I�3�xcok�����N�@��5n!gMG�QaD~�ӟ���5��(���9x�eG�8|x�ci脆�IV#�P����wtD�wP�:`�FW
�i"SS����C��Ϫ���[Ρ��8��&Dwh�V�D�{H�ڒ\�x�S���f��3
�d��%J�7X�Q��O�_^�4��@�&���	�c�"���:^[7�Ջ�J�m�Edr�"O>}�<��i9�F���A�C�I�h�B
;%H�;�d�6#�4��L�0^��!Ŋ�<�-���Ë>����y}{��#y鵷�/�|������<,'�ݯa���Fz��w�С�}�DL�9�t��������X҆�J∺�����'���������/<-W�_�7_?�F�&����zi���[Vc� 	S�b ���T�Px g/^e�}�v���k�"4|r�*����R�79���a��rU��G�����<������߼ 7ՐD�Ii@N��Ԓ��@f�}��9�I"�7 .%kZ@�Zb��|�0[]��{D�"g��ӝz�lF ��`�е��=F�6~R����7
��W����;(c3�����lm���Ͽ(�f乯=+'�[榦���	$*�G	�=]�P����&�޳��d�q ��!�M�(�<��C�	C���%i�g@ؼ�>�cǎ���i=1r��-�=��Ո|��{y�}�"��Hm$F{hD�}3��Z�f礏&�!��6j ���$NOβ��1����ɼ�i��Mi�r��9q�T4��I+*i�+q��,�)WŢ���b�1!�C����^
~i�T�}�X���)R,�s�Ңl5D�b�@�H�&@s�&�J�mc�!�����O��R]�������u�3�۲g�~����6�ޘ��]Q�|����_���KЇh~-w�~Θ���X�:sM�����ܽ�O�𿖯����ݿO����5ʗ��K��hț�@�:W.�;p%�h��������|��'%E�<��p'�
X���j��RP��7�!O~�i	�;~�����%?�����w���ѳzMj,��"�~g=�ϑ��OI���dq�Ӽ��,����3��r�1K���2Y8úo��|���׿�cX��TFKL��'��Rg<LG4�)Do�ב8�+�k��ڍ�j"��υD��ڦl�;�����+غu������?�'>&�{������EYZ�V-]��S��?��ߓ�͞����e�f�����-]9y����g�\�����z}/V%nmʗ�u����OdQ=������R�����(@�����Ѐ�~6o�I_���IZ�ʌS��נA\�[�˧�~���gdy�.s�w�g>����t�cy�7��Ǘ5��R$؄�P�Ϋ��!��!�dv��x���DIO������N0Y:39ΪL�r�eӇ�m�4Eb�\�fy=i�^�"?{�M9wmU�aT�G���o�+�ߒ�xX������_�\�= T��ɒ��a�>���5(;C���L�uׅp��W��޽,���|�����^���QV�Z�^��!/����go��1Ay��[���E�+7���R����Wn��)�=��D9���x<Uc"D6�4>U��'��}4|ْ?����?yI�u-�f�;0Ax�%���{K�z&�]�!���΅�R�� �;c�-�<�.E����Q�r'��c�v�Db�������Ǌx �/�e?��2,���ծ�<N���Up�tKh(*�&#	ʫ�ƦsS̗�����6%���e�ݖ�M��dρC�[���,�ɟ���%9�s�Q�η�(�=z���k�kP2S?���K���E9���|�s��s��?��L⢓�������'�K�IE�@��i�2�1�g�Ԅk���g����y��� �A�WA�{��p�}�x�'O����my�s��!�ɩY�׾�����,�/]7�_�@��4j�Bd\"���J`WʼX��.�!�d��Gz�j�^��G�I����Y��iMڃ!�K�iм8%�vN^;u^.�i�˒�RP�
��W��}9�a׳�~S^|�\|＆m�FIy�ڀ�o�4X�̋��cT�m�`L^�����M���-�/?zY6���|�n9�w��wח7b������g����3���P._��F$!����iy����g������ʫoI������7�&e*7h�_���k���{���>�����p�&�8/���v����v�� [S��C��ԏC:ܟ^�۪-��Z%c��x���1�7�;�`�#KT�&,���{��U%��w(8紘e+ZG��E����X�l��g�Ƥ���|�����Ĕ���4vGi�-�y�(:rei]�훓�?󐜿��u�M͎ɗ�����OO�Ζ�9��N�U1�s�����/H����'O�o�������|�_�{��/[ۺ�?:��l���� *w�I�*C:RF=��ܲ��&�R7��:-��m�z�v��T��z 5�v��������o~���&tט�o����T�[#��F7v�<�ɊR���}���,�.�[ ���I��V�Hu��i�.()�L!10�8�.]^�W^;-gί���p }+%H�v%�0pSC�_�������3W=c,��E�LBU�H�T}n�����̫����x�������o�{�D�(J�7�6���5��J�yS$�����,����O�5c���J��_�-�ﻭe9�j������>�ǲ�^�PeukU.޸&De�r4ă�0���%���G�>zO�W�K<�O��@0��;?Pl���x �_���R2�]�S�G����~�-ٿ�G�&�nrK�)�\,�����0�jlBM�(oz���A��s��^��Wbzf^~��?�s�/�$V����1��ruL.\�&?z�E���������wO�{�!����q=*��GW�����.�������˯$���Yy�c��/<%G���D~�ȟ�����~"˺�r�i��wb�zAۤIVJ�hŃai�ۘ�LA%AY�ס�t��ڛ�V���'N�$(��@�J��sꍽ��9Yk�u,��W(�T9��X&��8�Uxȕ>Y���#éXeH]Zp�^�~S��X�T}��#A'�Hy�Il^C���y��wu�nʥ�M���3r�Ε��ht�V�g�xY���rs}M���gU�o���h�)K�PU�����n�y@�������Mh� �ms5�箯��+���vxJ���z�)C���լw�'L���5S���:6N�ߵ�%��+XT�\���FO?[�!G�lP�$�w�������F�P�/�O����{"��fX1Ϙ��s�h�Qs�bȭ�gc;bD�\}��R���?��> ��}�F����ыH2�q�)AY��_�q�����Q.Bt�\���pa'�YE�������?�2Y��D>!��_�@��X��C,SXJ��Ѩ�X�([���ٟ�5�V��ܗdr��<X�$� ��~tU����uU�S/c���"W�,(?{�y�Ȝ�W�n~�~V���/Ͽ������O��7�<1E�iX9)���w�Ǣ;��0ƶ��!�<T�S1��\gc�ۧ5�����Bh#�aN?��.gGv7*9f��!�*2���8���"�zh��dgOu�9�5�Y+�F�XR����peq����E��Y�N���'���
!��n���[2П!q
��fk�\��@^�����M*��o� +�F>	�7�0ݹ�b8�vX����4��գ �h���T�p�r�9�X��F�L�UT�����5�h�eۡ�B�8����\"i��2���)t�S�=*3�'�	b�}"��%�ɣ[�&g��p�f?�>���=xOn�{�vK����Q֩�u8$0e_"���PI��<+g ����L�� ��e(��ۛR��N�ǥ��~���|���-[_M�.d��by��M-�j�'h!W�+:��( u�?4rA_��Ņ�.���/��NҬ��^׸zB
�qB�Ӿ�@|\���������\�����������)y_]״0&-=9�D%�*�Z�*o������%��(�26>΁<���r��"2O���Վ��K2dk�b��m'�ǣ;gsn>j>ESg�����2.t�~`�x���� ��'z�]g�/a�1Й��k�N<�4%�	���% L��P�y���rb�
Ati���<�Q���R���ؚ�1����艩߁���Lɛ��eX�ޮ\���G��xD��^�����Szz��3�
����a�9H�����O����U,R��s�{Uu��I�<�A0Z����uë���ݳ��`�����rU�}H�y�P�H�=~O{}k~s>`C��I�a-mLvT�p�B=; �KԳI����$]�a��s��ÁD�m4"��N���IjAD�6�����Ő-�����%��p��Z���I�����{�{����Edx�OsQS+2��T����2	R�!�G���||�*O-F��uD��
�Ơ\���������?��jjV6CX�C�'���{���sM]�x�j���+�����
���64SsRџA&M�NnC�ɒ��}��n���<.Q��.�'�cC�5�C�h��]� ;4���L��2:�����_���� ͞���{���i��1�_�FΞ�dުP���9��h��Ƚe��0eĠ�6~&_0t�|��8�iR��s�,�w��]R�av�֠6̟0���g�d	W.�lN<�f����^`m \���W�z�ΐ6���-/;�t��n}d�aE�Url!dy�ԭ�T<5�i�$��G@��7�'I�wr�ډFfmp|�-6�u���HGA��ʻ���6�hb�HG�h7����F���u.�]����NGj}T\�߃)��N(���drd�۱���E�Օت�y��xX��I.T��.���I�DL�U�~G��Ģ���Cɭ%�0�Tv�He�8*ڏ��H�+�cehF�LoP>QN����K�ʎ���=
�)yO�� 3$��������n�����C��1�G��IőBY�rÏ�*#ǞOF�|%$��X��v����X�������H~`�:u�&e��N�.kNd�F�n����|�4��۬0�?"νC��S�Uq����3�#$���n��4�϶)c
IWТ��׸�ъ�x���aD�z��7$A-�2���[,��,4$,@��_��3f��@��k�/��F�Vb���#E<=��l����	� C#p{C"�8�K�a�m����؀@�������ĩ��,����ý|
�Ɉx�}�94���	F���dhE$p�GɌ��ķ\�OR���10*���K �呰õ*�)�A�k:�~�}�\�}G��ݮ���~Ï��w���9���a'�Qx�G�d����7nq����o&2�P�J�o@//�'�������� n�d]��&v,�Q#���(t��+pd�6���,�g��o�V��ɶt;����`⽎�8f����z��ۍ���I�&G�Dth^��� &���
�)�Kve����y7CbU���PRoz �nNpو�8���A�
3\X#���a������ݮ8K��v?w��?�G�${?Ҥ;��~p=�����#3H�g�&�#�����!�� D���q^^�%�Л�n��޼w���ݭi�y���O��@�.{d�o4���3��p�YN���L(�
�O�8?��!f����k��'��wQG]F��`��g�6Hd��Z�B4gU �(�q!1��S�7�q����h=���Cw2v��8����b�`֊�줁�B���A�Y�2:��7o@܉(i�ХƸ���Y��3�\n_e3�F����>�q2�r`�,�..������.ao��+� �gv����wx�޺��d����[:\Ax���6��N"4�|F2�dx��'�y82�Y�c�c���򭡋#}^�^<H�Г},�*B��p���<��s�oYx8�0���ȵe�B}�Q/���P��!�H>"v�1�'�j$�G�~����%["C�Rܝ�@��5��P��um� ���<P@�!Z�K�7n���#�c�NdrTd����\$P����E�~��-�f�#�̵E߇߄����zQLzt�tg�gk8,#����m\>F�/X��Y��|M��'�F G#���,nghv{.�k���T@��S��Z�pKΌ�DO�fҐ�H�|���K#��8��73�'ޣ��0��vF�#C#�	э�h��稼z���FH/�uJ'�=ƃ8K������`xp'��n<3!E�<��O?�Y���$��r"���/aH�3@OU|�&��vn���\�v�.���%��GI	��ԕװ1C��:���w,U����8~����j'�F�$V*$\�]���d�ӕͳg�8� 76�B
E�7)'(�-.f�}����M&��ZB�6��ߡ�|2r�I��x��f����ܔ���.���dx=I�Q�i�U�x�`�1�Si��D-��G+���ω�����aIx�����xo�^\�7�q�%&!���Oy>����BO�n�|t�9��b����LF���r2�@��B��I�lH���p����\4y�k�Sz~4t}u���Mo�xg�� �@*�nO�FQ/NF�Y���<^ӝNdGN���C:x��2���Ĥ.��6�m��QK�ŪY�r��|b����6���n`.�����(��'��#�w��޸Ntf�Y�R�6����-���C��y
�d����&Ho=%�5�Ek�g�9wv�?eD�N����2�K��ڙ	��[�8��M'�j\(wx�hRq�{i!���c��,��Il3d9�$�����HG��a;n]��!ʝ�=y�m?t�Ӡ���n0p\w#�4|�膺��{K�¯��>5ࢸЇ3i6O�|�3�_���]�eȀ8��,�:�Z��a�əz����F�����At�7$��HuƢ�<C��c��x=�7%�G����hYVc!g @�p�on�G��ˋ�~6��Ѐ4]�`R���������~���Ro���19�-���_Ð�C���{�|�tE�I�۽���L��+vƖ�go�����H3��HO��d������}o��n�ѯ���od�uK!jw�p�;�Τ��`$��97�b-�14;�G�O�<w���ar{0;���04&lL�F9�y=�;c�3&��.�X�*����rsd+d�855%�z��'��'��e���In��R���h֗8�2_|�Q˼ّ��g81H�56�v�����5t7ԣB-�&@صm���i���P�K��u�x������8:@��щdG�m��|ʯr�|r��e'{0�aL~�1���w{��GcI���n�ao�ˎ�k�|�� ��w�̷�U����/BRiI=��6W��/��.۸>a���'��۽q�u��g�]gt����'������`8Υ��y"��������td]f��ޗ�������^�T�b��=a����4Z}i��1=�XMw|���;M�t�읉0����k�I�E�k�d?��I�b�B�%�vKX�h�ꁀ�k߾9q�||�l��Ic0��v����rF�oct���|硛���1���;��0=�yw���g��lM�n[���ɜ]��p�\�aԈ )��2�~�����v5�l㍖�%�����;p3J�
������V#��ȸ�u�O{�2b�v�`x�#'�O���B7���}�����tgL) �"5�>����>H:�A��B��%�(t�ܨ�
<5�p��N�~N�[�p��b����8֪�B�!
YYdn!<p\ A�$j�����9�9���V�I��-�x������o�e�ޕ�=�ad�HrGO~�G�iv�5��K ��q���./�`.�#�����c�O��ޜF�=�odIO�����6�Q����\��?'�{�#1ۋ�{C"w|�9�<� �J�#3p+R�^��+�^�w$��	�ql�;��:��+2C�H��3�B@o~� >LC^_�##�s����Xe�� ��t��5��E�-W��cG�!Y�=;o��:7?;IBq8��[g�Mj�fFD܂��"Y�#�2&<)�S''�E^Q�/�o���M^�9r��4L��t��	b�������F���Z�H�Pw{Q����޻yA���_��0�;�Β��^-�!z���com���I������{�ۈ�ݷ���#�7|Y2|�����12Ω7���t�da�]�U�\�ʑK�놣�)=�F�&kt����9���Άnh�����������'�2!�鴍
!wNZ�x,{ sjw�d\��;$A��7n"������	��&�M~�J|�a
�A�'��~R�q��i�Q4���SO.����ZX�1��n�V�b��=�-$4\����`��u<1R�>iЩ���
'��a1F.G��Ż�;:(ݚ�9,C���냇�Q�e������j����u�ЩK@��l�����ڎ��>���}X�݇]���cOS $
(��YYY�2"C�߽��^��H`�i��Y���|G}�"����FvZt�d,���L�ZS8w%2��0����os��~�d�=�����f}t���]�e��0��j׀�ٙ���$���.���#�yfF�Ppa�I�F����WC�r�����E���z�j��l-ܫ�V���3Y�\5�ő�%4Q�6^���o���{��oA�+g2���A���p���ѸDZ$��>ܥ3mÁ�`r��X���i`���iGg�D.&�r�q�7���#����qj��{��[�p"i�SQ]�"TD6d&N!&¥`~O����<��%�}\ 7%i�K��0�8m�<i�_����j�m�^E�	��Vh�Z����5�t١'�Z�4��׿�����`�p��jN4�0~-�e*B��{@߯�q��?���|�:���/A���'������.��9��3����-u�F5Mi�|�ԵdDy�I��Q(�ay�l�C�%A3_[�2�K)�3Z����{E��TX�$���.?�إU���fh�?F��+f�����J��Xt�kܹ��&wvh���g���e��W?���y]�v���\�e��3�y�X����L��9��+vC~mgZ'�S�Ee]���(m�v�O�D�Ӯ`f�W���(�.A���׊3�������
�3	�5���u�c���!����H����z)�k�S�]�yN���+��gK�(�d]�Gϳ:�Ydĵi]���E��j\�jS�E=χ!�B_k��F�9%,J�J F������(*�AK̩�exK���}_���R�ذ�S,%���Q�C����K�d��r=OI�HiSǪ�ZJ�o��\ɖ���<��Do[JQe�+��U_��?���`_�(���jG|����k]����GV�P(NМO��?�i��#�Zv��El��rG�!63�8�=��(�I��T~=.XYD5W/d��ű�a���YytZ��3���E���)"f�u�?�!{����%	�"���">�}lU\��q�	m7��N��jt֢IO�
I$�����|�\v��Y�W�}[3oK�Ǳdv�tS�fF-F���I�2��L>RjI��r��d�Ǝf�jʦ��#��<r�b�,6��DʪH��.�����F�Mh��(����=�f�K��fk|o}�i�f0}6	��S:��M#a�"3gES�	�nԂ2X�>�W*!�6
�(^��vw�B����l�w��K��E������I���Zp�S|�\�������=ymT���pZ�9>�3A��He-g'�j~�~*���x���73Zٛ����s�q���L ��)E�� ��T<��Rƾ���1k����H�lW�FBnS���?�	0d۷}.�Jwi1ɟg��8�s�<���2;��V4a�ԜI���]9IB��	G�P�qe��jtZ�����lb׌�w�Z�6���s�9��{-���!߁�^R�:�j�595ߥ��Bj�����/�X�5sm8�N��hĆ����|�IM�Χ�) +h��8#���Cմͧl���ƥ1U�K��)5�����FRp)�$��:6+$PP����um`�O�q6n^Q��:V�������VSrj���A[�x>�R;c��W�.���R�J����t���N[��������Kq�D$"4��i�.62O�!��i�c����i u<��q6���&2�J��L+�{�d���"G4�ܯ�b��X���{}�Y���q¡k��*iӢu��m!+>\W,$o�]sS1�>��d��q(�8-��H�)�fJé2+J���=qz$�-�e�3]3_�Q=.
Mk��(�A��G��$�9�JN�'9hy�EJ�?�pI�p��ɴ,��ֲ�K兴u:׮��\�ۼ�_$Q����թ_D�Θ��[��U�6�2���ri��X|$��h��ܟ�8�0au GԆ�"���I'#���L�f�c�v�CK%����%��ܬQ�mZ��,R���Mo�WY��Ӣ��ҙh���(��|]�2F�	������GB"t�mh+��s�%�@aQ�.���1{;{��tN���͞��	:��k�w��s��ة,��%���B�Ҝ������Ґ��6Q�;Nl����H������rs����ð\�Ψ\�kq?�fW�����RBʎ"�dŕ��8S�����8q����2h��pD˅�!*��.Y�����Wt����:�<Բf�qɝ��=�P	�ո�E٪hƹ�5>'�w�>9M���%�eI����M윘e���>_�[[[Q���DtO@h����oC'�g_�"�x�f�7٢�/���`i[5*L���S��L\JD��\f�j�\�|ܬEf��>x!�1y���-&�ETp�p��8Հ�UJo�:=���T��/�&+ĉ��Z�n������:��SR��Ao4��|�5N�����d�;�k5O�1]��mN�����V�� mA�eBM�����%(�<7Ś!�0_ߒ��[]G�� �--��̚/�,�3�H
H�y�A,�>��9q�ө����,�ﻑq-*�	���k��'�be�+ie���� ����C�d��ql:�B�	)�8Z^ ��,hA*�q��R���`���9jB��$�: ��lJ�ސǫ\�ES��K����p�!bo�St~{�x��B�3���wMЫv(�|�������$'Of�KV�k�θx]��5����]�� �ƒ����ĩ{��L'6a�����hTSC�pD�Q�jNG��X}s�-B�1��9��ХIڽ��#��0���,�['�.��M�ؽ�d^5�t��v�h&	[N���n��V)Z�zw�'�#̕���Qb+3���T6�X�B��.}�N|��ۈ�V�uPr}�u�I
����'����T$�)�k9oU�Gն�/�3efŹB����b)m4��Xqec,t?"��*�*�#<�߈�Q� \r�{�3�EAr_�ʱD%yU�AX�<3Pi�}'��wv{t~^�2h��W�w���_�{D^{_�G�)��D�$��L���|^q1+�J\#�d3�9KY��T)�Yc��ǜ�|���z�E�BU0)����EX�+:u�Q� �qb�tac�j6��	l#+j)	yk\�F�\�edXD':53D$p��˞��	���x�����\�a:�d��w,V�3p�ϥ�隘��� f-\'�0d��6�r����B�U�D=[$T�!/
���̚��ZrI@v��o-X_�e:w½�o ��1�)PBtY�r�8�Y�ZmI���n��4�!�B��\,�4�bG>E#�Wi�Z��Va[�@]��^��0(骚��[ԭ6��-��?{�_Ѡ�3��r��t�0Aa)��?c���Zc��0�se���y�A����VC��pA�^�B��>���@K뎭@j-hq�9��lOj����M'E���C">.r�i>�������%�]i�`9������&)xG�������K����_E4��]deF��6J�5��5
�l\]�|�#�ZY
R�ZӒ�� ����i�'?�=V�ъ%��kI�})��)��\��+��t�����Ef:~�F�P����R�f�����R���,I(piK�,`��_L����7�ﱒ999���)��3=n�U���R��4����g>�t���K�o(\Q	��89B`Tq���h�)��U���+^%�B��Q2��ݾs�v�:��Z�-�z����HC�����W��3:8s�(��졓a�#KWžцZ��eޢfX�Ȣb�&.ٺn�c�GE
1>gٿ���U�pF�$�!M63������<�vS�����T��7�.ܜѤ�͙|�3OH��*J��­B�V�U�0r��L���@�6�\1�]V�S�m�ͨ�gX��	��"p��O+��QrP� M�I |�,�{"(Q�P��|��B�V�Ưt�q>h,���9`NPo�)f-2ڂC�$3����F]0%}d�7��%+��*�Q\!ބ	�J��RmyC����ڰH�Es`�Xt80G0C��{�.}��u���eA�������̨f�����ҽ{����o�2ݥ�E@�-�]�F���rs�k7�hr1	�=�C/�y�0'P��.��Bpask�Iw>ZMi��L�Am2���������o���qAO_��d9��`�M�����C�6�����z���$w�`��L��<�dB��A����h��BDҤ�ò(�|b��9�?w�Q\T�.�9e����	��FG� ����%���6�dVV�tn��F�p���j٘��O��)�*(jqs��]�'S��NNQ��K��ٹ�&�a�|��jΉ?E�u�a�o*]�$�";Y/����JX���N�����*�ўf�_G�@� ��p�pn��ϠB�)3Y�NQpk�s]�r�����h����=-��{܊�+�9L�Fa
E+sv@���T���H;�ZCEv���h+J��R�e�2&�n���߿���>���V�vВ� �����~?n ���{k+�١[7�6�k��A)�XLI�/�S(�RUi��2i��#�@�M��v���"(�=���m���_�[zy0�����G��τ̻h �X8�㡏	n�.kҽ�R�C|{�[lQ��XU���r�I-H޲4���͖S)��
���,����B��a�RIr�|
�EXn�	'�8� ࠝ��Y��ՆF�
�X����	Ъt9~E��%=|xw�.λ�O/_m1�ovN�yX� �Ga3�1��U�/�F}MQ� K�u�@4���t�UA�`Â��2x���z���6	��Ϡ����y!��O�'׬��n�x$���=`��̴�N���d�����hwo�n޼��9==	��0K��3T��"5����䅮aN��Ƞ�%"�W7⬄p���&j#f����¥ڛ�Im��K�Q�$����;)se+��	�ٴ%��"`����fD@x���a<�[BՖ@B=��*�א���G������wz1e�\u��p4�dM,�gMH⃖e�.oF���g�˩�A;�t֌��F4AԄ{���)��%M�(QPf(qm��=����^e�룉�Ղ�x�C�t��5��܍�Xe���v����0=@H��#�<(eJ
hf��lr�wiBD�2V�ҵVAË��I%&
�trL?���������?�ݝk������xCG�:x��^�>���#�&�X\O�C'آ�7l�%7�Zr.CU����`��e�Ǧ�B�Mn8��貰�	#$��󀲒�S����g~'�d���,ѱ�`�Xc��;��償����=�א�䃀D6YXM&r�R���NJ�c�¸.�>�vk����Gx5��āf��$U��R,��Fl�(����+�J�"U�v���oa₫]��	 	!�W}rl����e����R\g�Rf2��Ԕ�w�u(�71��.i_4���o�,�~H����0>�_�?��p�SA������)}������=�?�n@�'s�M1��{T�S��p~�w62Ѽ&5#�Ikn��to��V0��C Bi7x����p*�`�u�}FA����.��$T'�,�VS2eיS�o.jn3�ś�����~��p�!�v��>��G���o� �I;ۀr�̙����O��{�(-f7C�`_���3/�� 0�ӫ��1A���"
��E��!aP����>����U8�����7tt���LT[n�l�R{�X��R�ђ���F�״�x��KD'trz!5Hlb��4Z��ߐ�ُ�>�$D��%7S��p/���P$o��d~��zI"��{��ˋ��R�륕A���K�3�j��'��2s���/_b]��ȅZ�k��]�D$��O)[9{7:��DuJLT�~A��������������$��F\w�]����_-!��e�FQ��Z��� `j��:�#�$6_��[�Wj�B�4�0o�V�_�0/�rz@�����7��ۜ����7�� ���m��"H�?�o��t���������q��{����8bMP9��i�&KaHZu��ˋ1�h�r��H�������� "�"��6r@	�4@��ͬ��>-Ҙ'F�ep ��47�>۬��D�.��E������^J���q:�&y�͋�ER��E��!J�E{��fJ�EO�dT`X�O!&��f�D��o��xֿ;�CbOF�2n�b��o}��	m��M��#]�Nd��L���q��X	��d���Ru	u��/"��,o�SdY3�G!��K��Y=�IX糰f7�ש��8�Q󰁧P0.%7Q�inVr����}�zv�ɯf�A�ᲅP�
�:+�L>��9�5�D�kl�矈+'�n[BU��q�d�q����ɧ�Q����$��#����:��f�� ����!$W�]fJ3s�}HL+�d(��A���(ex��+��}6[H2���\:��H�`iTK�iς�����l6��v�ƠiE)�4�.�8��n����{
�:�uEX�7���+��Сe��#(�n�.���&mִ�==���?b�js@�)gH�Q�*R�G�&S�-���R����3Ē �-TO�ߤ��BD2h˘���L��b[W���Y-�aN�}��e!��<}$0������>��	����T:�G�x=^��'�k��niy�FK?":Z92�d�|{H�`�<\S|[���Y09���"
ޕ^��rI�,,�6I�(�mQۢ��៼/��q�7�ymP�fA�јE����t}�h�%15�)���Ţ�0��b��e�"I)�I+�B�%�͹�HXqM�B��Z�>x�sR#/�E2
9_�d4�,��c�p�Ύܗ�Ė�����v~��t�2ҳ�0b]�����d`�b�P�8̕"���V�9��E梐I�^�[���t3�[Z�w-�zJ��B�5�Է��n;/E��M+�s�k��7A�j���i�7؆�:jF��12�L?[�q�8fQ�D�`c���xk�d!>���x�53b��蓏?��ڤ�~������o�3آ�bƾ<�$,VB��b�&���M)ۋ��9����Q�;	��] �;��''������ki�HL���ô��
Y��2�3H��GrtQ�����dcjy�r�:s���,���Z7p�LY"�}M��Nx��x�uq��_ח�(�pŦ��C����W���`�|�łCLbI|_2`m�7�.���洤�pd����r5-��vy��jg����9_.Ca�Z�ޱN7��ڗڳ�(��*E�\,���LVh
�Ǿ,��Lk�ōa��h�P�\�)��*q�-_��],��*ih֍j��G��i���t�	,���H͒D��oe�.5�b�bs��u�xO�WX�����K�3��2��8��B�FY���@q[ش����'?�+��������$(�^@,��L��Cq�T��ET@m!"��ơpΊ�⾳uG�t�A7�<�`N]��?QΤ�w�~B9{"�i�B B0=����2���$�m9e�޲R�l��1�i��DHo��k�B����2�z�!TZh��S� !Vx�DZ沰��M[H5h���6�.Y\�T��[ך�5&��̈́H69����>�[d����AY��w��@r�9��d�É3����F@�-k���1v*|.9#�ڴ�o��(h���6t��	�d:�xO�߲ע6����l }bQ+�Tb�Ul�T�s��'	mM�b_`/	|�%5�|*�t^�m�灔`=[(����D��2j�B6��$�N;=*Br&�2"gʣMZd�б�'��c�A��jA;�;���[4���tJ���ʬ!+1�{��"�4��Y�h�)dL=�t�N�(!DQ;�t���=ͱ�8��l���I�?�/ϸP���Ft�	�9�vr~��I`�/'��D-bTJ������~�n�4 �>�z@�p?� �L%=ڥX̴z��C��;DA"���&���o��w�z�W�}^�-�ò�<߫���4�7Aa����(�����"���� #��浚�QX*_��S���+����؛��k��uNM��\6Ȝ���S
2o���2�&"��HQ��a�Q��#^�SL��}#y�a]QH�����J2S��m�3Ǫd4O��$���u��e���7@��;��a�67aL�u��益k�|����qʞ�5��>��
��P!�#y	eC� =�]ϑ0Ӌ�\a���2dem�}6�&�)�~AQ���Ϫ��\�h$�ś�V'(��g���j�l��pH2IXh�]���}�2m���ޞ,�dh0[|���k��ta擙����B�l|�9�G#ж��ǐ�kL˽�υG"~M��.f��M��HL�|*}���Ϙ��J̤K.?�\.�O�]�E�Z�>C��L�0qz�T�M����>|�yr�i�FN�H�$H�t�&&Y��T���6*:V��ii)悐�z$9V�h�����9��"��,\�s�u���"��^��0${�!k\����e¼�dCr��0I�T���<oH��#���$9����jH�o;>J�֝�8*��!�Z7��H<���<W}?OOO�l����c4ߓb�<i�k��:c��6"6V2o2���(ֿ�)�1�h(�"�i��M��2!E�q�J0�
c���R�-�,�;�*T��s��pL�Ӯ�4��n�(Sˉ��W)U��ur�	+�A���y�ML�'��+Z���G%HQH�hk�@��Z�s�!�$ɑlװ�l�b��x�*�ʹ��Kދ�F،����Y1?J�kn��Ǩ���޾=�e@)x��#Rk^u��\�vm������/L7D�,˨6:I�,TIJ��e����2�gO�Z����5�N����5�}&�ii���"���������t�N���2��jU�w-$�Ze'�O�m�B��έ!]%����2�M��&�2ڼKfH6�n�}Mɜv^q��2i�/
I�'�1�j�U�Oϓ}W�9��k^��; Gq��M`�K�_���lkx���F2||�ƵY�rM���X4*{3
G^�E�oP
����V4��m�z{<�_BX>�z�s�y�8����m,�,u�S�n��>�on�VK�9�,� �I����O�\��AyA�`n���u_��X=�\G�����Y!�W�,��-5��D���X_���~�h�\��	e��5��)�����'�`Np�r�&+1Ma�
F�>8�A���&"�Q��M����u3E �ا���lt.?ֿCI �&EԦx�|��m��m- ?1�旜ޢe:��%��r�2R��M�9Q�����lVE�5�!��"����%�_h
zLfL�N���o{��ɳ��x��c�ؿ������C�o�jo�eϪ�'2�dk;��$a���dH��@�|9�yVw�s>J'p}�4��(�>���gm���ﻈ�X�fl,P�es�ԉ��)I�td|")��to�z�m�|�1	w��4�

׆֙JBdŋ��|޾}K�﫰�9QG�bw{=����kz�&H���ؙ���Z��5S�ً�)�@U�Y��J*rE�A�wd2}�+�ay�?�9�WJ�hzɰ�B��Q^�d�|���~��_��R�	��o�ɯ>��|������W
]��*��$#i����L�诘��2�U�)j�3Ea�φ%eB�e�To2�����6�v����_
F<b*g�ưK�a�#�%�V�~5(p���������Q� een�rVc#�&�XUD��О\���z��Fú�<�Q+NX�ӧT{=��#L��/��B
ys�\�&\�/�}Ls��m�F�	�[,5)}�P3���cn��|&�׉c�Y���Ѕe���) �L����c^tT�P+���,�ROgZJaLV+\r�E	��P��l�'�P��M�ʺ���暃�ޯ	�_�N����l!R(�$�����f����lɫP��o�a��+kc$����Ge������K���*�p��6��_�{���=j	D��S��޻����Ͱ$�I�0MB��ǫ�s?o;����KN�Lc�W/�5�+�(P2�B�s�f��i؇��zAq.;]@x'����b�+��Ã��⽋���{�)5Wj��������k����8������m�j�:"*�9ͦ��vQkt��Zs����LC�)�"���{�б�{�$Z̋~I5r=���+����h��p��p��X���PG#DE�՝�R�*EX	6}n(n/��0�ob��kf�9��E��X�tHS�c�`-�F�,D@��1���QX��m�U0�zcNȪs��G9J1�%�M8�H��������ЭD!T��m�	�!~v�h�w�m�	���m�KM#�%�o����94��|89�LXy-05��4~�Mh�nV���`i%��_9�u1*�s�����%S�+���>(jZ�b�fa��s�˫j�8�������L=�Ŕ�/t��-]���ԜJ\���.	,�7�~z!��	���Q)���y�XP\K��Eu���HHc!��A�k"c��^�@��,���g��"
R3��]�>�H�+�*X���ߧ�=^Cw����#XǇ��&�9��"�/!R6�2R��6��o�KZ�y�ENDS�B��ڐ1(�@���#��FZ�i,�ib
�yۅ��6�	9���|�z+���GC�.�#9���3#�V�o5?	��jE�YZz1�	�tv���%k�*α��"omI��I��c�7�N\�M��MG��|�W-|�z��K�c��`*�]>'�_���}��.�1���p�r�X�Z{���R�)�ڴ:�K�Z4�}M�2J;�=R�&�̅hʤ�Z�M�4C4�T���q?�	6{����ZNW�3��:�|�o	�:a���%)�.�n��h�W[��iK�G��n!��������D����tQeli�R��y'J-�B�j�U?��x�l��MQ�Ońv=��	Q2��J������������='��5y�\��vX�"�m�g�b2�9�;�h&�,��&ZW�r�I��m6�bxy����dT����J���c��ו�q�d�΃�(�Y#Ʋ����;d{|�~� ɯo�[v>Q.u�� c�u�6�J���l;��^5���Y?	��1��U}u��>�JV��ߣg��:H���L�Xt���S|c����څ�=/�yBՈ7۩���d�HJ���m��c���pf��_ju�\.۔-�Q|�ۚ��� �����S֦>w���lsk�&PD6.�3�i屄�H7�k�su��F�HC�4~|?3�H���v��!�Gm$ ��A���(~	3=U翯����}땴ǜV:'�wD^�T4��?�`rϥ���|gME5�$oF��.�F�����Ŷ7��LT��t�ST_0
���2vXӒN�;�yM{�2'�Ip�}��~.q��o!J�����Zќ�[X��ѐA�Di�t�!0�E�o��{-��, �NLǓ/���I�w�N�@K^�LUO)Z���*�g\��ICԾ�j?��j>H�%����NjFT����J�2;_����a_Rm�S��_��5Uf~$�!��cf�OFIޚ>yΗR�z}n0�%G.���omT�YK�s��\BkW-�vU7Q��� J,[)ѝ*i��"�U3�uk��;�ϑ}E�N�W�ML���"�\P��U��٥߂��E#WǨ��J$�L-�RB��S��X��	󲢯�?������?���]=o䲵�?�?���SHT��t�'�͘x�/Y)��O�D���b��(�m{Ց�B����bd�#��5�4DrY�V|h�,{�I"Ҧ��͖���c'"�!t��Dk�:ا�B����kt�3f1/ă�ޭ���Z��{�����c�ӄV�*��M���IZ�5��B�TCż�j�@��9�Ƨ���씴�Κ�K��y�e}B0�_�X�������U�����!����\�5�ū ;+�+���5��Z�Yh�]|L��9I�����e[�!
��W2����@&�ӹl���bޱV0?L�����9�-��׏6��ߌ�l�t5Y�@f�ھX{�(�c�4	]gJ�af���C9�O�	�'p�o��<y��N��HH9��-��p����|3g7����\���E`�N�G��&�^�lf�h������K�W&|�������1�Fͳc��S-���`Q�Rt%#���"$�����=٩a��X&:Eg��%�4.���g(]4����E3k�KqC�y���}ßbu!dZߨ�2a`���ߺ#n�KI�y��BɊ[9�"R�����ca���M�����	�q����"׉
PF͚��j1}��T�"�%���	=J)���Ѷ�8�!��:�_�%P�p/�V����fw��wo�jou`��Uy8�u<t���#���O�Ţ��Tp�Z.4�b�#�o�6����V���i��fӚ����&-�8��Y�4.vݐ��Uȫy~f�e<O���0Y�)�P;�r��'��O��ٜ8]m2}+1(id1 i�p#����i��q���0Źq�呓>w�:�S��=)y�{�_��E�)���#5�����5����x��f6.�n�86ƜD��]�6V.΅*�Y�ְ�_i�7��
��`4��C�uDᦹ!��A�ɑ�d|s�@U�>c�g �b�3B7ǹV��s&k��Qӯ�࿡	�L4�Z(�!��Tp��`��ԭ<!_�$C/ۺ3F.5�*�P�\��,���@�Ϡ�'SmWy���P\K�f�� �	��yгnmXP`ޮ���63x��M"q���'���	@u�����Zs�b�4�}.�����u�
a���B���f�4W��.i,f�/S1Y�dZ�/^�K��F���h�]zڲX��]6�^�׫ �7�NL��BD93��|�¿(��J6����Rp��b6�:��-���Oh�,���L�%�B1W��A��NUKޓ*��Sz��M��`�+}��(���2Z7[Wd\x�($7]hMD��z�4Q��X�&G�ū���=v����a0=׺��Ó6"���h��R!�2g4RGYj�'y�}�FV��pRW�mDC06)i<(�[^�<h�f7)��u�yr�Ȏ���(1�D!BW,r�|\�0/��Y��B*�*6C:�_rC�q~��:q�u��c�;�|�&|�e�N&���")�˩C�_!D��d!�����q.S��9%}fzG*H�&�B'˕af6mSR6>_��_C�~��i@]5`�g����]��e����5�zO�ňDL��=�}�"��Й�(D�e�h�%ݟr�yr;6N��c�1�n�6QUGz^��J�F7�K5��W<�������S�����C�n8���tI���'s+��䱱��DW�U�)�|������d�*�����bR4��~�+�C��~�W�4�'nb�~_&�D�[���;o|'�z���'IP��/�z�\v�\�}Δ��9/��Mb}���X8V�Ω٩���}�9A�Ħ���� �3CB4���=�T��/��"���a���W(�O�o��	J��Y'��ͷ�{!^�	qh�P=�o�Gj���b�]�ݵ&	a��А������6*8���I��	�F̛���Rڤ^��	�
�v>B�IK��ґ�EdmL[�[!˹������4�� ���D"΂���q����R�l<����eǕ"ϓ��?o���Z��5M逘i��H�b6c:�|��{]�Y��'Z%TB���v9meI���5��xbl�.k����?��A��&f���9Z��Ӵ��kyn���7�u���oɴ�I�8ښTQu$�����dʣ�V+:R"�*b���bo� ��c�?`��?�s&e�֑D� �ly��Zw�a�Z�%E��&8��[�̚H9	J�mޭ{QP$�[�,��M곽�iݙYK5ɎO?�զ��/W��&a�����5bϚ$�F��گ�$6s���=�3��t+R�jvߗ�7v4$����W!�f!2�w.��[R B��e-{����|���i�
�֡U�s����,�P7��ad]B��A�L~4��?��Ry�:#�g.%g
yZ[[�d�T�Ƙ[B�H�$\����[�U!�Wm�}(����wa�Z�Q�)�G4W�Ԏ(���IhM2@�jW2H,��I A���F����|�>���;�Ѽ $aQg-r�e�,L1��D���ޅH��u�9��m��Ӿ��xN��̈́��|Y�B�#��P��&Mz��*��u
eT�s�oE]�4�����,B͂Z���S�U��\��#�7���>���^	A��^�((�G歴z�B;�9�`��JF��>��^w$¸V�S4�+�$����4�F9>
�/#���?Y��I�sc��$ר��|���lܼ�9+�L~F�Ô�$�f���\�Z gi�{U����E��ۊ9?VA��E#��<[X�N���z�.��XR�����ˢ����8��/����h�yI����H��͍A���7�&e�����f�Ǐ��e˪UyR
Y^�=�����i|�dJ,���w)=v!�!�x{iY{��Y�rq��@�|#�A�j�/��u���$i��(����� 9-�>%��>�:����J��9�Ȥ9���)�/ʂ!~YK�� @�WU��/O1iU����$�ط,߅�_e�d��Od��J��/�@fW�~r�_ϳr�C`w�@\�|��R�*L�2��y�E��Xm  ��IDAT�j�8�<A��E����Z0�Z�Q��&��*t3�+Lj��ý"D���~�Z��1ZQ�\��+��%�����i��8v�p��1󣱢8<7�E��8�K��x�r���4�S�H��<} �Kd�>٦ATxI���ȱQ!R�z��=�����&��l�l&�e�2V�.����p>=皃hk]���EL*jg������G���r`�&L��`�ϋ�LS�$�\�eV�ʜp⒎��!EH?����퓆G��0؝�FҺ��&D�ӧ��l�9��/Ґ��zغhp���i�5�(�~~"�l"� � Ip�l�ο@��P�.)��b\�W�:�*ݏ�ڵ�~%�*�%���r�3-ũ.���Z_�Ґ}�0wE�b�Q;(oNT�.�*���lN�
JGtQ�	
F��y%ܐ��c�ϒ����ʈ�e��քl�2�۾��se�n��ӠBH��M��1eS���D�$�T����:�rOT�mݰn�P9B��O��Τ�Q�$џ��rh���f׮���'o%?e�����y�QJ��m�3�h4}�G��c�z<n��	�a��FN�mb�6�@SF�Ծt�a�oIV�S�-/UH����G�������a(�����a�{��[��ާ��ug�EZ��Lh�1g��^䡨	=Of�Z)/����H@�jY3�L�Ө�������y ǹ�y8��7
;\s$)� ���eg�\k��Y�kx�]�ٔ =��!�z��:;k+K�Nk��E�a�k�����+��^���-3�`��KIg`��Jᯊ-$�Dh&tI�dȦ�X5���B�0��<~xo{g#u��C���EH@�\M���k�ʟ��t�����+te3�}�BDY��sV����j[Ά��i"cگVY
���a���"��"I�,��8�4�B���洍�m!�yfL_J�)4�x	��l���b�4M�8Lֶ�i2��G�Mlm��� :������C�~RL��d_����p�/gR 7u��!RK�R���jJE�YM�st8��o����CMh��S�!8x�4�&���5{�{�wm�6w���3�-���׻}�RQ�2�p�L�CJco��#�.d��-S1�A$���:g�H-�/�S�N.�:
�=�� �{��w�?O���N���� D�����LQ�G6'��W�d�8??��A,
�Eר�Ռ��#8�e���3a��e�H
���H�bq����B-�t��� ���d6[��bƿY�4��s����2.�	���3]��aQv��R�#_7V���daTKn�ɅI�_$߃��X�	����#����?Z�/����:��8��V=����G����㖒uK?h5yt<��1����o��xG'�'t1�P���`�Z��f���Y��_�6M�$hRT��������G7nޤ���h�Z@){�4m���O0�sX��R�:���x�l�'nSB*d��<�B�[�isc�����D�}��ph�
�M�L�ڹ�_��Y$�Kٯ�]� �q|������T.._E���ƈN�����_�����tX�؇5�[l0�>�;3o��9:MҤ�O���F7� 8? ��p�n�^PAEӋ)�1:zwL�)M'3zs��&�)�-� 1a�x�ྐྵ.b*8ʅ
͍�u�}��=��?�aQ������߃'Z�9�:b�(�|����5���]�/�܊�*��2���y���-��%r�p�:ސ�k¸���ћ��������;A2>�"h�I�0�9tJ8j�x�O��GU+�-����̧DǇ�^Ћ��a쇴��E�?�Gw?�Kۻ��u�|`�xMB�xF$����tC��L�"O�Jދ�˷,X30�Ue��LS\��
m�P��8����+���S�w�D@ȍ&�149V��*��U�L��xɮN�M]k,����<I4ݣY��=(�^�GzAR�_��؈�lYQ�B
�.tM&W��<��������^����)i�$�{��&�������x����8;=���v��#;�q�~!�� ���:!N��?B�B!͠����٦��h{o7h�]���_i��g��ML^C�$Ĺ&�	N�܍ΧX��8KxzщP&���{��bL�9˻���w��(S�o��h���T���=���p������Wo���}:ºY4Z�KAXXh]C��R�V��o�a���+�F��Y4��|ü��{����0���ڷO��ݛt�΍���M�^�����?8es�2Zݚr��8f1�HfB�qC7|�N!�^H��R���^���t��d�m�KT�B�{�k��}%�c$in�.:���g�:%)ř�Ѳ_w"��5����PM(�$?�=E��x��k������-��s�� ���l]M����)
	�����V�.O23ɛ6S���`�Ӓ5;�?�X�Ɠ:=���9��Ũ�<؉K�*��G�E��0y������m;ǻw�Ї>d?���)���л�w4	����>yE�nlЭ;����;�y�&��n�f@-p�B�@"����B�5�*�N��N{��H*����m$��r�1�g&9�|\h"�
5�,�R��w�_��B�Tb��,�a������壯h��kF|Π����CK~~����K����19ʘ^r���4K��C�Юl��`*��9=s���߾F|x�>��!ݺ}��n@�=��Y�6�r���\o��	r�P�Q��}�Dg�mX�p	?��� i�y���7De�X��+^
�y�'��I�т�:��y{�|"�fz@K�ч�	�F��!�h�EF:�O&��B�$6�$�ԗB�8P��Z����z-������0�]t�
��E}�a��CrA��l�����t���3���v63�I��/�@	�g!h���[q�Ļ7���O��~�����7_C�}�-�ys@g�"P޾{K�o��,@���� �_������{��G�6�dg�+� �^LXHh�!�wU���6�f��
w1�R>�d�eډ7�9��0��*�?��"��3�9��k��ݽ�Ύ����+��o��O�ońu?o��|V�rj,Tj|�.�!^��i�%�"�Q�%Y��W�j���Rh�M�Ntg����6�����ӝ�w�ֽ�ac��{>���d ��n+T�0�9����c-�ώ>���]Q]�y������	 �٢�
�elF��z�z���ßǘ�Wc4fj����x���a�N�c
[���}8�_c��i98Vk��ƕ6~�쪕
)��x�������aCW� ��]�M��$ ����������+:>>�΢��˨��ك��jb����D�^݈'�����@?��_�������L���|=nͱ�y��x���^��÷���s�<@�'���Y�г�y@'׃ �H�L�>'4`n�bf�����)��qH�}a`Nt'E3S3O$dl�݆ӝ)����y�T����c�4E�v�!<���]�׏��o��t���O�i��J�e�!-#H���ҦSP.��S<gG���+��m"4�V'N��7�s6�x<	�xN_�5�;��?�S�vX��f���6Y����Z�"�P��O�ȑ:��*(���0� ĝ��/�Nu�u{��Xu��M��pʳ7�:��� !�C��r�,�I1�}�}�Wz�ȻPq��g��)*���{nd(�Ѳ�p�U���)c�!D�\�%��	�g��@�1�����/��gO���k4U�^�h��g��8����%���,�f��WN������?������>|�ܹg��樆Tt6h2;��O׮���)����������/�����>�w/�i��ǟ��w}��=�E=|@w�ߠ2�?s�I�[g�B��w�8�m��S�]���j3yqy�LV��2X],"�&]�� �߈�.�C�U
F�A�sz����z�5}������K��ܢ[4f$;���,a2@\�3�K2�z@AZ)|��r���:���74���xA8!�;2�6v�I$k�>G�)�1:|߳`�>��;:�����~����K��Y..��@�<�kT3*���&4��\D!�k�#S��e������qW�]v��s��8s�a���
sR,�,H�cCv��[��~dU�R�h��R��YC�2��h+(˝?��(gd0XLKG?��1��se�^e�^Jy<Oz�kDX��K�����g�=�Azr S�9:A�WM�����qq�I�X�Bg�DJ����/��~��'$�
{��ߍ�w��I��]��� qdJ�n���ӫ�w����t�M̨Ã� �_A�������m��a!��0Fs&u� E3��^��'��*�Cl�b�+A���>�iB�w�(%l�!O_+�i���el �'��ߧ���=��Ex���/�7���]:>=���Z? ��9Q��M~��Tz�0o=`}n���ƚ��3Sz-cq������A�k��q�E���^�(��&�n'���0'G���9�8��&��`J�S^;I֐&/j�"����W����c�����	�bX�UF!���u�C�[�+~�B�-���\�ۏa���m��
rdl-ٞm!�)2�����>��?�0xE-A"6�9.OgS��,�A����1
c�^s��������yC_|��~��?Ћg���5�6?W�jҹ\P���?\�IMR�F8��)����l˪O��ߣ�@�L�x�yMӓU�mt��l,�&u(��C�[7����t��-/N$��������=}��n߼M��n���&],�A�J�B',�%�֚W�2���$2�9�
��8�rT��� Ԏ�/�ۡ6^뮖�����{A�=�OO�yA/��8o������_��o�������Ux�;���>}��[z��)ͱ9{%���n"��skxK���ѐ�L���<�y���g,�p֍�qd��n��p�v=��������Y^�Og��7�ь�TI?��!+���"�j���Ea
Z|΢����|ʎ.$�diNV�aQWd����U�C�Rn�z���oЮ�{��^������ƭ���
�M� Hl��<�(ذ�~��k�Z`(�Tϭ�8�d����<�G�$���~��מ�$��Z�G�ƥ��ݰ̠�sZi�3�Y	��N[+���Mm�5�/��۠���?���_�l2gN�^@c��KK�;]6�?l��B9 ��Ɋw6�اZqZG'������.��!=��`wd���]�$9���4gu@�n�ҋ�Ϲ�b��`Mg���.��xA�>�]�f�R�Qm���a��Aa���7V�	Sjjp�UC��F��N.��{/�ϊ�4��*\�+4ZPح�~���f���+z��	��v@a=����/��F�-}�7���%m_�E�������>͚)�!���U���p�_);�|HH�Ӷ�����Y�"1
\@PK�d���e�$�0��'����.
��p�W�~�(�O�����DKX̝���G����-Wu�F2+(&$�p8h�H��_})2W��Q���U�8�]l���O}C����������O6���x:���!ݼ~�:��,w��<I(�bz�]Q���&��Ka�j�n�0(�_�n��t���`�4g6+�!8 ����Q�|t�P"�<ʾ]c[@�2�tMO6d5�������=�}����o��w������XEՓN_D +W�`6�)�R'�X#r+�p�0'�����C,K6�6$��ؠ�A�����H1'�m�x�p���'�U�;�0&��6��ڨ��"�p
����إ�EDS*���3�� q�Z"H�F��e0��`�q.��G;ܱ��d�%س�q��'/���t%�3�{�^��`�jHsm����J��l4WwDnZ��?<������G���(�n$�6^���:}���V����)������۰�����85��T�,1gX����fgЪh�m���2�Z�����@ns�?|/��9�1>��Vм���6�؞=��Q��{���`�J�һ|�s���g��f�`�΍IiȂ��	i�8̭
��J#�h���J��*6�/ �BJ:�W�ì�u0-O�bP�*�}Ce8k4��}����^�i���>
��7�]q��==���#�������F�$� �w�g6FI'G�������&,�)M�Ǡ�)�L`HA�X�\�U�c�	F(�-�f�WvY��:�5�%ݻ�}���hB/NK >����aL�$r��4���#/Id���~F�Sz������v�;=�,���߇�-��tZH:|W�F��j�
�B����x��O<>c�Lb��d�_{�a�0 $�A�UC:����g�i:Y����������c��H�k�f��i�ߦ�`Ȋ cr̛�����Q��	��X'ݠ�;\��y�cs2)��%d;������s>�b��V���\��A��4���ax)a��R>��T���?����~��!�{��thBoL��JYԽr%�'5���1zP�6���T|�z�?a�Z#3�H����G)����"���Q���Ic�/��N���y����X����8 ��T�D4.FL�P7hZ��@h� L��>��}���/����if^� )Y�0�6|+��
N]��"�
Mpb�&������3�F���p�.}��t��]�U�'�Dw~v�,sbq��oN�L��t����	Bdș�\�	���j���<y���1&����ܥ{ݡ�~@�-���:��[ �/lL�U��?��A)����2�I���/Jmi�cΏ!����M�ֿ�C��Gӽ�P=�9!(f
���5�?��Y�[�=F
����[AL�g�8�J�����ݦ\2D練���~��ń��UY�lD����0'�<�49-���cɻ���,�&�%���ˆ��Bq�$)s?���/�\6r��.�A!}��R�&E�G#�ڹ����t�%�Y�6�w� .�wf�W"�����0�K����d��	�j0l��1<If����2���!��OV($���v!�ERwe1C�� �AȜg''�@~���� ش�߀�[u��Tr��Y@����a�
����{{k3��CF"�j#��`�n�O?��C"v�j��@�Syv:��uG���n�������߈�ԍ�	����b�Z�yMG'D��:���&�7�y�(M0�z%�e����XZ�g�7��/HZlJ�JꩯA��A�l�/k���ï,�y��'stx�g���}p�^Xx���ANw��~>���j�p����ao��}g�Z@.���p�}?��.P���D���r,6��	S�@���u������r��I��vר�!eC��^���g���k:=?�q��M���T�W�Bo�`G���쌞����߸F�?�,�I]�聊����L�q��8S���k��R��m�oG����)P�"�d�r��(��D)7��#"��ZjE$�e�J��"�X��z�>�������m��r������>o��Ŝ>��#�կ~E�GǱ	�?J�{}1e��$M^V
+�Drc�o���f�S/t/\���pl;>��=��'��4чӊÍ�{�X��N ��Cju��{x���m:���x��Ԫુ���'���%=��ݸ�C��r|�Ԝ̅z�L*b's�6�ĕ�*�	�xP�)�1̢	�7�ς�[	�"��N�^�������}��ǟRU;:?:��b�&���`�5�Ԭц��8|e��Nէ����`m����=�M�rԇM��dg��
H�
�~�T[��i?��.��1W����I~���;z�����z��4�Po���#1�YּP@�����D"Y���	}���t��]�y�f�C�zN���u�J��E�"�r�Z�U�`� 9/��~ߎ�vP���;jb����z/ڴ��D���z���ſR/�Ũ�p�m��3���[�E$N'ī}���51��x�ٓg�����y(���֕	�;�"�)�=����8�R9Iā~�&�����b.�퍽 ��"�O���mـ^����,�c��S	hIH,sr[��8VQ��pSf�F���Ӌo0i�T� l�ex��W_��N�>���a����	�~Г��ϐ�l9M��5:�#���'¹���H���'�v�z�Iw������7����Ɲ`�푛�O-;�(g\XA��@���B�I��b*����95�D�3�&x���`w�t0m*�`����n�0D�ε����a��ɧA���ͣ��#�t��\�A��8�Qp�"J���i@N]I��G  �z~~L_>z����F��F%Iݗ
�d&�R|R��{�����u��?���B�S������cf\�}�V��Y�YJF➛�@uy"�1���g��l�E�ـ�o�$��СU��la�xa��؆�����È���8u2i3� �M�����������K9�J{��N�����lY�Ih�q]�=�.����v�l�p^M/�ݡ�7�� <��E{��	��t���x6��>�^Hs���~��]s��C��a/$�'��Ϋ-N5cm(tMfo_��Ք���~����~�>��`#�����1F���t^�B�&�Lu�`���eNWF�E0�<����_ӓ��i|tA�rD���o�ȿ̭p���T��b���0���B$����=��F�$x\`��y��&��0���C�rEk��y9	�\a��w����{���3[�����>��/Z�F���r�'��UM�Zȏ�pϳ�o�2�x/_>�'O����$(�!]�O$|�U�i7��R;jGϊi#{�]1�����D��>���{!~ƛ1�M"=���h�%`���� ����7��rݶ�R�A�7�?6{��3�4�5�	޼�X�9z}�w�D�4QyM���c�4&���!A�R��|~������&5��k
Su�1w��o�Eo����99
d@A�t���J���g���'�! `U��)#V�<�l�\ۻΑ���.��2q�e�y$S�0!θ�'_�.4C����0��w�`�ڳ��H=C^HW�����2(��M����k�n0���	y�h���	+m�D�B�	)�Zh�0�j�ֿٰGz�dM��\ 4>zwB�~�5}��/��hL����������]�
� <-���L���$,��M�t��*�I���p���4!,��,�suӅi��&֤��p~D����6�ݸN�nߢ��=z�}��#^�� ��Zl! h�<��I3~ar�}E�Q�e�lՆP�2�Ǐ�{�N�	7[�3OMUZ������#��J�/I���N0׮�� hu��o'+4�%o�U1�]���VҌ����t�2�*�j���6�^h�����f0%%�3؊���M���J=��K�u0
�2x�n�1V��<��8�ϣ�6��$t���$� ��74CQJ[�������:@ ~)������,h8R��b
鱰�J+�W�@���ɺL.L��3,�k�׃��
ς0n0�:�`�� ��@.��9ܦa�M�w'G�~Nhs{�����>�4[ۂ���ѐ��<g6��0cx�ͭ]���9Z�֪�D�]L��L����+��� Qp>Y��o�F~L;A����.'�-gBm&��A�w��Ig�bM�ٓ92E�����_~E����0{/I@�?|I_<��nݺK[lS���3}s�BNm��<�ih�� �H�[D����>(�;[� ����5����N�F��yi@Q��5�����~��p@o޾�O���`�"��u$��.PЈ��osh��cF��!�,����?�l^3R���&�o^ѳg���;7���$�����/�Ȟ�yǿ��y�!Xm�1r0ɹ��{��B���[,���(�����_�D�6��-j�ͪ�Ǜ��Ȑ��d��9E)IG�i31�2�'3�H4W�D3�\�$����U��B]�8����SL�$@�8=����4����z��9#P����)��;oK�Ae,��ݲ�!�ͭ-N��[~Qq�ɰ�ɭ��&l� �P��a���&m����䌾z�5���k�,D�Q����3��X���q�FX�[��w6��� �w��3��Y�`'���t,�iH���v������k#l��^қ�wt�>�̥�gWH�IV֗&3c8�(~F�.����f��;y��j�z=A�A[_���l�9=}��nݸM{;���ng�o�܌=�
L�Y&̝��DU6Fa^n�pCf���tt|D��<s�o�.;|W�ד�����sp�	x������d���D�=����qZ��k��i`�|��e�L��B��8��ޙL����k���3��|��El���5� 1��i%j���et&3%����L������3�
M#��Y0@J&�)�}�^���b@[[iw�0�23R���0�l��L�5K����a�!�m	�&:��n�<�d���%F��"Lx��B�BR����y�R~��	}��K�堅��gg%����`` P 8 4F���:#�0�v胻�;�9�sr:��@��d�� �՝d8B{lmoS�*ܣ7��BoN�^r~���d��p����q@'[���$���j�U/���~�2�� ��rV�w/�Sa-��������-������	}���~�����³i�%?o@���f�f��R�q/���1�x��[dG}q�g@#���	}������t��u�4�.�����������f�C|`A螞t5�E�(hlO��?�P5��Q�o��y�NOi̕�0�0��s�#�r07���!@SA�̗��^,�Bq�qs�M�@1G��AH����+:E�*���zb�O&��& �ͭ>�V1�2?SĖ��/#su�N�K�
*@�Y��2���6��Yө��XX�3x��̆�&U
�F��2��e�@o&f�Z��)�e��x;-�7g��-�"��d�
��JrM�<�9u|���j�e��P����4��Q��,���F��w�**����O�aA;�!��!"\,��* R�N0]�:nv����޸K������Lض�7^����q����7����1}��[:��x���Z#Cu�o��{{��>sIX�5�{��v{�������]�w�&M΃�<=��p�l�
���ss5�M����0�=}A;�w��m��3i���[�df��5��Q�S(��0Ϟ>�q�昏rA:�����|�^���?�~0!�v�@yw(hMX��M�t�`w(��H+���YR�klw�U;��X�/4�.�p�+�߇�	698��<�gΎ�r���?��&'͚ʭ $z
������5��%mo�r���LN�Q�?d�4x�|���wA\�d��-���ޱ�`�	��`�RW�4i�_q��������6�Z!���-i�!~N�c�b��Q��n�4o$f����jN<|���h��W��l $M.Z[�Y�곛�e��A6J�|0��u�J��;���{ce�ݱ�D���C�A�vAA�EP+���،	�Z��D`:(�ڠ��nѭk��@�t<e#L�� D�g�`o0{�߾�(���K:8>���� �%:`[�?8a�nold6��{�ѻc��O8�]�vdl�`�LΖa����~�3z{� ���rY4��]%���q7�=��~����E$���i�֐7�R����+���9���6��3OG�����o�.�NY�:�8uD���O��;AH���C��Ϣ7��l�!S��s�:����c�Y@��vi�
P�eq^�/x�n��.��X� rg7iL��I�>½�d�V�tN��QZ59-��aY��W�y��2�;�kȞ��&Z���s_�ߑI8ǃ�89}�E0����-�`&���{ �����c��J��Z�ؑ�2�a�B��&Dlޭ�������X�1U�=v����������7n���zv
�j!vNrꒋ�6�N��Y����l��˄�.fi.�E�Z�^�=�,Uw��y%���'�=�$ɒ�0{�3R���]�5=j��|!���s�� x�XpwG�.]�3C�ڽf�GVU�p=9����	{f׮]��^�����s2.� uQ��3�'��� \�����
Փhg�+[���X�|.w���� �����ē�[;��j��O�ի7���@�w4�2<�j�5�I�әY�H#}�z'�j� ]݀=h�f����;�������ZO�|��;�ۭ;�tJ�5<(�� ����k�:����r���<x|(�o�(�ʔЙ�!�(6W�e^�q(Ûr{.}l� ��l%��/��⊆ �%�*ҦG� �c� :�X��7��^ts=y�HC�w��j< ��,���BeK�w�j�I\�7F6�h���P#����w���J_Kƥg4��$ᚐ��'��{�Lg��cB�d���^���4]�1�wu>'r��rV���H�x��:��^��b����T�c�Z����ayi�{xa��P4�bM���E�j(�xp��6$��Z�]��+ￋjf�u�s�v�����}+/`�i��ࡊ�/��GB�Q��.9	��5�:�`�s ���K g�t��j��V�Trv�/���vWe�	s�fa80��%�����J�͈ๅ�ޕ7���]��ņr~�VޫG����z %u#���a�Jٙ7���g�ɸ3���{�������g�0r������A�  z�+�ۛ	A5��k]8g7�Ak����)���A\$'�k�߯������I�i�}��xwO����O%S���]���H<��FO��X�<��<<z-W�S���aŶ�RZch�����M�j�1=�칼�0�gO��ѱ�H�U3C�QЇ6�gG*+>K�20K.Q7��~0"�:Ԩ�!a��q��z^��*�)s�{�A|T~ԭaG���~&���9�{���ͺ�@�.�j�A���x��O�f~+�z�E�fHׯ�3���v�C2��w#��6g�-���U��>�f�A,����1+@nD/�5RЕ�~�Hm.]��r�pq�b��*`Wֹ�iAc����\���K9<��}56/HJ��Ʋ(lU��;��*����,�����t�2O'���@
����l�A06u�UR�c_� ����8_�{���a�nf�����-�����B㉈$b��cuA#Knؔ�n��N��|"���Tl��Qѩ�����=Q4%�N�4�F+h' &f6�ʅ���ł�V85#���n"�S�ڠ�m<ڗ��9�;�d�P���TT-�-�c��M�(r]�!�r�`�qg��h"oȍ�k��F_�L�l�ް���8ң#00�#g,Z���<��z����>�Bޞ���b9-i�Y��Toe [30��i$��7o�Pxz�d��G��i\�t�Eo�=M�pY����[����h�����S� �۷��=�ư�Ps��~��?���_��<��Z� �c�-6�;�����~Fy�)HF����A�/ a �5Q ��w[C���Y,��z5�e�(�յP.|�YDO���F7��i�vp�#��8���%�cHL@��ox�m�@�Xnc%[� ���rEp`�'k���\�3�CB6����B2Tx�Hk�qϦVhLRO�#��)ߩ����Y�`u��+�i}J��J.޲%��t��&&c����{4��1�T�OQ]E��������WQ!���z(T�\|�4NcŖ�d��:�>g֣UOQT��<�Ǐ�]�_ɛg�L�g�P +���� ����q�Ҽ1(��{���N�����R3�`�ú!�G9ŋ���F^C���Tޫ^�n$��U�=�2���DίOe� )M7wXA �[�a(��!��(��b��n&�z�����r;_���܊�ٹ��W�k��*�.��;�'��4V	��B�(��	�T�~�;5ֵ�5DA��F���q=@J�Iby<N��}�����H� ���L=��T�>�TCPdE`���eL+o�5#ŋz��P�:��J"�)x�*�����+�c�鯄�Y
[[z�xMX-��6lQ�����@�#g|)i�o��+g1�p����f���&�	����y���Gx��?TV\Hlư ��7 ��ȯ��|���=K�V� �U���ʅl픍��b��">�@�z��T�O�������zDBxld��s-O��� uÂ���X-gl����f+�c��5�]�������ݧ8���lv�����ꕞ�9�2�zp��� 4���{�x�b��z�C�P]zxx�8��`�����W8��.��p�qT��|�d6��)J��^�wvI5&D�w�3����Խ{�ٳ����{�2�<���N͍^[9���\`ab�`c�(q��s<j72�өqM�*�� q�+�� �w�hT��\��Y�Fcj��W�i��px�G1�:�u���oe���`I�' bҦ�$JvfFT\�L��ɭ�\�J�wr�!�xgGn�Y�S� p0"P�G�$�	��47WCe.Y�c��~0B�\"�쫋y�	q ���X ʃ�I2Ф*o`V��t%��sE�.G{� ��l�����փ�rJ}|���ǥ �ӷ����Vbz�zh/F��޿���9���~�V�g25O����@I)^�/�g�kBEƢ�2c�ƴ��O�اTn�B�rO��eXEL ����N�H����X�r~�b�Ք�F��:����q}f'����kW��=��:���y��	y"��N"���l6��Ò,S�!	ނ ����Ya$6*�	&�J7��-V�` ��=Aށ$_]Y�M���V�2N�rw��48�*#����ǲ��/�ח2��������+�O������YW#�d�	�^�P��HL�GO5��̴��>[<�{�ׁ�@�������Ra7o�tk� ��N?a+<�oo.Y�Z�vbuo�^k`VK���f���Jج0�,�б\y�5�Z���t���C��q���������� n�PZs2������k��{��	�#����(���� "��������T� ��N�N=8�y�}�EE�SW��Kq��K̀0Ԫ���%zf�kZ��u���1g�?wI����4h�q#�׼QI���`hL����^P��K����ܐۿ��c��޸��1J�d�RZ��x�x�	�$#�0��S-�XOa�>	҂cdd��yz�s�У1jx�:������C�'�wPӱ��`��J7���9��ǐ�CCf1���W/�˛�7A��
�[�q3�&�>B��}�(���r�c0\ B!�x|t_�n��ZO�X��%��;���Z�x�N����*A��c��Hk^"&�kbɺ��J${� ��!e5/ o��C�P���x[=�=Vծqx����\-QDXz �W���z Q��7$�"}<�����Y��֙P70>��U�ã�F��N�|�jm���-YS�{zKϾ�R��ߕ���r9?7�4�����H|e�$3=���5A_E>B���k�#C�}�X!�x;5��ă��}|����-8!���3恘A1յ� ���2��E��-D�x��XI*Pժ���Z�u"�a�;�3 D���n�&�b�2�_H�^JH�`�l_) �75M�G����J�qzb!�h�b���Yw)5ر�n^�P7�����DNs�������j�BS�^�4j���Q����O���������O��S�\��;��ѡ��5{���`g_p�}��R��f�!�|�TO��E�C"R�{z2!.ES!Hx"_��s��e������ژ����b���C��z'�7�����] <��M�%,l�c�6�,*���k;�;N�*\�G���k����Gד��y�W�^Ӑ�H�b	�:��q2U��9�mk����-�HG�r��"�l��6C�`/�Y���>�Y�c��L���om��'O䷿� @����V���#�-2�c�m8Ahډd�o��JTRgH���n�p�[�tD?V�F��C6^�<����<�+�S�&DT���n�@���r ���% >�ma#;���\�Br�H�fTu��F��L����� ��wbhޙc!�nt�ޞو7^yLZ�MH,dȾ���:�)�ɩc���ĺ<�!�PרOB=��б�_Lo�A�Pw���xg9_���O�9����G���w���A��b����B�3k�����T��?�o~�.�P 9q�������c��4�P��'���U1�l���7�)��5J��z�k=��{$�}����z��<�&퓬uqvE9����@��rAc�5@K
צ�e�w�r\���.�9%�'��\+�1�W���c����ĮX�����jZ9N���3��Y��\ZX��5��	&�Aӿ�o�4(�:��A������B(�v!�j�F:�0��EA~��V"Ãb>���C=>�����|��,��;}5�x�� v����͖�ڪ|K�,b|D�^�?�t����yn�3W��{kW�J]���*�(��������1�F�/���1��B��J�4���;�e	$��34IS�]�dxBH����
�ƛ��<�=��k��n���Ly8�9�6P�����h̢��Ex"��S�ӭ���50���d����{ ���b3#(���{��r}sM��$x:�^EN
=�@���}N�
HlA����}����{��a�D=,�bP�(����t�+y���+=�.x��N�e�{���/on)��tk'kj+�p�v��w_�4Ǔ��YTmi�7�D�X T>�y]2���B�5t���mZ�
��b�e���tl����Dˁe���ǅT����d2���Cv^	���g�5U��xX��������o��`�(P�ﳷ�+����� �7����Lcp�Ƚ��\�}$0Y�$�OS��e
���Z�g��3{�l����)&�����Ad�-Jf���54�w�ܵ��(�\�$X�y3$�u&`���6\���w��aJ�V�Y{B��xO��;Ҿ��q�W.Iب\�3R��*�"ܪ~HziF�C������}��kC���>N��Y�J<7V�z�$v�<�6�� ��p�����{�B��M,��N_�w���7D�����^V�iM�\4��/笿�ʌ�(�xJ������B7�6���D��<b��r��E=�Z�L7�4��5����8}q
Ϧ�^�{��7C��|1��o_ғ1���Ǳav��$�桯�v̠�{>w���6� �>�1��!����g�	�9]o�3ln]�b����!^������J�4[�Vĭh�Ԣ쨗,�b�H%xC��qS��2S
@�W������,<j͈U��[Bʟ�d�VYFݑ�7h�H]X�����⩋q����O��۹�h�͵��6vՓ2�&�w����zýu�yӡ��QxH�����R|zsp�v��&�������̌��<��/v� ;���`�@��V�)�Q��Њ�D�&dSCo��BU�*�'+Cn�XD`��ݭ�	�V��k�&q�R4�2Ab%i��fX*<�T�B0��B7r�IAJ�+�i���֔��1�(-�r�}.v�G������b��Y0B�!!��LKVRN�;8��a{�rw�y�衯�C�A赡�׶ZW����:�L��.ӳ�-�� ��]��`����l�����6�/^��4(��չ�_���;g(�Td���7PzܮA�&h��҅Q�7��$��6��d1m	��Ct����!�7���Nt<�ڍ��1�������9�p=�^ݺFe������Nfv8Q̮����p��@
BW�lF�`ǻ5�&�#5�Ql�=ThD�4�W�ᨻ�1D�vta�v��3Dx�L���>�:�׸W,��!~Z�-/ܺǙ��p#M�2��,u��5��n��XU�bh�g�H�2*u�X���{��b���!5Z�B3v4�v�l"���=�7Rq��ٙ�[N��Y�P$�]���a �G"ϩ:JS���1ں�D�7�Gz�\�mn�,VyǲE�b� �"�%���TYT3���o!#}4'#����Aq6Ӓ�FT��UE�Ϝ*YK~N-*O:�l�,���+u�54���%�;Ԧzuy}#W��L�p[����1h;��jk���Е��s��$;���=u�{Lk��=��:�չ�3+uG?N�d~)W���(%�He)�<�q��q�3kh��г`,����N*����z���'�fTp� *�f�8�W�vLIY� ��j���&� 2��Y�oX��A�;�Uzyc���e�p_v���F�����!��q#�J�.��W�͒�����dwo�M�YXX�֓F  ^���4^� ��:0����lqĺ�i'/�N:��*�y���r%;��KP֞�h��!\�E<��ǄEf��ާ}h ��� U��%���Ѯ<~r�{�Y+QH�Q�����۲|i3�B��$�%�geo1����`���`I�&� �i�!��G)y;+��];��ã*
w���d\Z�����S���L�o��И�|P��M4���
�uĈ�� To�y��O>��b�|���}�tf&}��~9YS�)�w��š�9k&�~�����d�|,v��uiF�ɨ����n����������Ꝩے�Ӹ4������w�+��}3��d$yTE"�DN���6��Kdulm� ;B \#����pu��58X�(vCI¢�ac�%[�17+,��x.B9\�s����⇗���R�j=cq���Gx��^����[b6�&�1���F �>ɘT	Ln��fX���ص!K"N�B����ʪ�ҡ�1Ld��h�϶���!���q3�M��		W淭�iL"f�1�D����_-���>��ZZ�a��������s�Ě��������X���f�VB�<�8��FZZ87���i����C,�hMfx�f��%���$3�Hlw`�x��[��A�d�N6�F6��H���32@��<��i��,���j�`�Y3�� V$臢�w�P=���o����с��-~�����淿��=u�QR�Fc���㖆Oy��f��!ٯ WxB�"�mGo /���,>����5V_~������F������Q(���x�FƓ�uL1ǹ<z�4G�@;�J,�0�	t�-&P�v)�PI�~���#��t1�'6�꘩����ݑB!_33�&�%;�o�b��3+�k�twx�6E�ʠ7f�
��8�Ú@|�Y(�|��`����2�D�7o߽�pf��AU5����Xkc�R���n�u5-�NҖj��K�X��g�����M8��O��Z��P�R��mI��3�MEs@G����h��b��{F�OΙ4`+T��//'r�Z�Ñ���ލ��f��֒�C֪�12���^ǐ�W�����Y8�cDW���奣���KA��������׃�:���pCWsk瘲���uq�����uQ��r���kV�2EJ^WG��/���La� U�t����n�-��-+�!�w����-�Z%��@G��_a�uz̶�3��=��W���o��o_~/�{���o��'�r*t��`՜����V��p�%�+Sn�-��8���&*���j83C<&r�0O=�<�����~�SD���sOѣ`ͺ�]_�R�u5�π&ʚbN=nZP�!�`�_H@�����K�?��
����a�Pǫk x3�F��ͧ�n]��@&��:z��<yз��+�J��0���^t~�/&�zBN�9�G��h��j�!J&{�C��߸����R.��Nn�d8�g/�uh�z��Tõ,�, U�/^�d��!02X��핼:}/�����\nt�/�x ��I�8�V��HAc��=~�F�ׁ�㍜��;wJU��{�h�ޏ�5���jIC����Y28��*�F��usVv�U�S7�u������澴���-<���qc�������M�v!V�:��YXJ0��ݯ�F�U��GrQ̔X~:K���R`c�]Հ��۶	�q�`XBZ�KصVAa��d��A�Ѹ:����ا�J�]V�ؠk�����Jd�̷�7
\Q`*c8�:���ɂ�%��,�t�A��Ew*쨈�)rvy*���L���<��Xn���E7�o��Q�����n��eܯ�4r%|����E{;�"v0dqa���֫�,t�vv4�ړ��D�J
c��B��7b�3t�-�B�-�?o@t<"�׿v~�������j4S5���`� ���k4��X�8�Fl�	=S���w�j@.�~����M�'97Ef�+l4ot��QW���y_[2�}LtN�WK��줗�iy��|�����,C�ʬ�r�����h�fQܨ��_��x�v=��Ț��*�EUx��+e���4%�,���r��K��1Z�k�s�1�'�&�.�ql�������`x����Q7�8I��30�����R7kw��<]]��cp,�qhsfDj#���ąQx�j�	�֯�*�e��A�b�@��<R��]/s���X=B��P �0e���ՄFJ!N��X5QR����8���XEZg�1�x��1�ْ~$�PSC��M��{�F\"�@whm5��A_����iy�����{9�x���:	j���,�:֍����.ޛ�+	겏�KhhS�wV鹺���#���&]��ɠO��P;;R�yrP5R'��'��bc&�6�[*\S��a���g�/km�+ߍ�����7,�d�Lo5��fӆ �����O�]/u1���JFz/�.��5S��� (
53��C��lϩ[ߔ��b���{�Fj��ɂ�4��h"~~}�B�>�ެ:����v<�@j-�/��;@�ռf:��A×�аf�s�"�?�b��[�!a�g�Wx�#=� ���"�M9�:y�16�"�9R4����n�y�L{Ͷ���[��l}hy��K��1���2�^n�ũW�6J�d��V��,�։'Ҝ��˭�u�GH�]Kˎ�%K��D�`�&]����O>��iŇ8-�
���Z��V��cӖ �Q�ɉi�� �E\�x��u݃��JnW���5ӊ 1=���߿�D��xF� �M������5�Y�����k΍�艺���LW����m'� ��k9������H��w����[]�s��]�'Ğ��i ��z�{���,Z��� ��\&K�|�k��ߐ�������c�h[��Y�����J�;�\��c��	-B^Q��@�!]Y��:4p��FD�ca+f����^2=����,��jB9`"xO�|4��U���  k�(XnHAO����rӟи��y���ș�3v��1CD�<̗zES���U�9A`T�R��e9@y?�|=�˛s5�z0\�'�	���l�X�^�C,]��%>�ia��'V���j��6�Y���6��\��}|��u�=0���?�7qf�����rl��� z���zgG��3Z�jݷ��P��%�b=�O� .+��3uhY3��rqI��F�C����#�uѦ \��ջ�y��%�"d�!Tɂ��jAxAO|�lNBx'CZڎ��z!�Ս��|���m�|�ݿ/�}���fCy��7:������r���V$��$Z���Y��v�Cu���/[;��(�h�}�Z���w�;�����Q���w|���TϣbٺNfa{����@ꚹ6E�����l9հ�B�TC���� �*փ �7���K��V��p��g�h��c�89��,��1iE�H�����63Q������W3���[Ӳz/�	�RÄ�kk�����eM�*s�o��P���a%7���_J�/����}9����������vz]_ݒ��V� ���ͮ>���z,�a��kp���[ 9���B�5�1H�_8�*W 3�x�Y��63�4��tז`��C�d|"���$̅��3�pN�~K'����i�9���~��w�C��]ց��Lsc���k�����G/�i\��/l��ZY����HMO6$9e�ŷ�����G��TC�S�~q\�V�] S��@�64M�R�e�u�x'ju:~�Ȳt�#�Z7�TOnK��@����޾��z��AU�@n@H��9@��<ؖ��B��3�/@jU�(��f��<�B$�A��?��u��7���#�wr���s��o����1�~�t�����Vc���>O��h,c�/�7X�*�=ݘ�/^�v�
�jC׳�0�$�9�l�q��Ѿ�����RX0p����I��h��{��>#����D(st�s^���-�-�)���)L`9[Y�y�"���L�x=�h��d����8.M���G� 33�hxU��n^��9Nkdo~x�R��5��8��(,��D
.~ֈ8?���� m:6z@�W�y������0���)�ĭ���a j7j�#@h��?(�ּ���u��چ!��x��LcR4���w?��#��}�NL���p����A�WJ|�B1�]�Y8d� Ȣ�s<x@����a��r�,�wɸ��~UM�}]7�Lb:��!Z�;�n�~⼴j0�2IJ�XXR��^NCH�uc�[S�����
�!���	�[�0� nf�o� �.�zJN�.$w��QL=Px)hq��3��?/i�..�t�"Ɔ�Ƥ٦�svzF�0���?��w���L�1o� ��*�O�yU�No"QzZvscV�vM��7���{��j9�~G��L� �4��If�#�vv��y%H=QÙ�W�i��*�r��9�M_B�7��q)\3��5R秗4"l��r��7��/tH)o�o��Go!!�K��Y(�w���1��rf��k�*ge�zk�\�B�p-�e�*nxC�6�W��I�$>�H��X�]�����r��Q��{��FC䐫Y�x5���;+�3�S��R��ͷ�v��v�W�A%8=4��ٽ$6bd���`2�0�mN6�X��!#�0Q��=	� ��ñ�tVp�3T|W��3���D<<!�Ւ)KS9�=������B������f2�k�!���5|�6���)CA{��T�YJGs�����ጉĬdwo��]��;�ذ�hK� E���=b���B���PÃ�� tz�!�/�!�A=�Ʌ�5�X�5 �)��S�Q,i���cn�v�v���?i̹��5��9�h���A�8 ��"��N���t)�^���wK�(p!�s��C��.�L������%�j��-��`��q����d����p;���[���2ș]X0 ���s9:�gX/�G�%n&��]݄0������\z��83�*Y�w��	[T�g�c���9�p�� 蛐������g�¤<�I�{*WFg�vM��t�d�[�52%���Q$����-�KT!�3Ș�fJ�0\�`x���4D��u��: �Z��#�1��J�`D�P������aΞCd>c��O�F��W|Cc��P��+�"D��s�X�*z�Z��	�rYMQ��	g8EB�5��FX���^���A�'�F�F�2�V��oZ/��A)�8����]��a�4JW��&1���R[��3�* =�UN.�MTZ�!���HDGGG�I\����&����h��7*=)ֺP�褍:����N�9h�\���L'y�F�Țjb�=1c J5(�&����.���T޼|C�����r|r�M4��b���,��� 7�b͆5��'��sX��l�m��fI����\]�uN���x]_do�*fbHZG�:g��H�y<�k%�ދ���O���{��Y;2��9Ѭ#s�8��@�.ҩx��~�s�ʫ�������.�3d`@%Hv2�]�W�a�c��������9���o����YG�G`�����$%.[�3]"剛j�1�|q�0��/nޓ���hde�%�(8Pxk�ם]h�ɠ?⁉/x�b]|�K�7�0���m�v�����O�Baڙ��B{�Z��vPi"��ZT`�#��X��c�{��´M��FG��t��	��=���4	�����ھ"h׎	�b���hېx�8��ϩ%�5���I*o��7�z/e��&E8��-�cAxS��%�:���[s3� )m������1�qd�x��o���t]�3�ѯ<7h�`�"�D�+�׃aW=�.�@�!�2�;�Br>�d>Q�����x��[�ecsH�[���{�T ��A�y�K��ͻ3y�ꝼ�ˢfI7,�4�qxt ��'_�aF]���m:�i.j�I$���'�鐨x TL#�:<>�����w���뛑MZ1�ӳ��<p�ⳏ�����~�����z�0�
�آvm�� s�c�ҵg�� *�! ��qG|F1����i�`�t.�!��:_Z�h�OqwCy��^��S�L���G
��Ȋ���QH���jX����s��sj`9/y����jJKl�#�����|�.�������*	
��qbސ��p/��ЎC�&�Y�9�5W����^5�+;Us��3`�{���b*+rJ�{������d�{#$�qa�t;a)n@�7�� q���pa͡r�ZV�"$	 �V{wȏ��
�ɍ�v�����N-�<^���[tc.�V-������bq��9��1�h]�� �q2Y�XC�	�,w	H3Ǽ/���1�����sc�^�i��_���L�֥������!��������b.56�X������}y�F�·�дGM�d��e�}�.��|�?<���6��l��_<�������)�z03�A��FЖ=;��o�y!;�{����P�����i�X���j���$����wl�6�8,�1�c�[Y��D�ؘ(��� �xhL��ke�`�:��P�\�䶿}H�6h������oȚ���둥�7s��C5$�4~��0d�;@@���{7,Â������Cɬ���GSGs��v��2i��q�D�	��A$�\�P�>��4jf��k�L$�h���Lg��6�F�/y�@j���~�0dhRc��N��fȒ{�yW���x�z�ℰ���i�v*�lvM�(�+���<�ݳ�w�P�=�RB%L�x4�12;��>,xAL�^�����z�D�V�Aڽ�^�G�-8(�8�zȐDʌ�7�i�29���{��qԀ��xN72A��>of{e�,d���ɣ�t<vW�^f*f��B綩Ց���N��W�E���;�x=g����[0poy(�M�bB���������d5��_���ʽ{����=���5�5CA�f��� �
TN��1�3D��`0�R�S\4$>�K*bK�V��WZS/Jw�j���h�DC�.7�����L�"�\�x"k�X?��y�����.�I�e�p-
���Xh��Q�1gA��٬�4EAf-�
W>��J_{d��$��Bf��6_�&Y�@#R�� �+X��� o�{�e1�IlH�'"���A*ߜ�����m�Bb��,~�??�>Bl.hH���HjS�@n|Mz�J��௅`򛗯�o�����0�BE��U���l���o��V��7�x:l�F.��낛5,��0Ђ�(沰�~U�^���s%�m-jaM*��v����|�����Np
��U���ˋ�wry�N~x�g��翗��o���-
�N�u���|03���l=��n�G�,����H��ghf�x8&���Vl��ޓ�P����o�7����������t�t:�?��?��E�$����+���\�3�������P����8�����o�5c�#��-A��Ye!�W�?l��� #����.�,͜��[,k����-3���2S�j����� ZB���_�������f��r�~FL�����L�Z��lǐ"n�O�DxlF��j���3ܠ�~�M�{D�����Ͳ^)�^^������U0���bB̆ ���ۂj��&@���ݕ��I$~�E�ʬr�TS&�=�ט�o7��J$�~c�[����T�G��@��왼y�ZzrC�{�V�7lƒ��P^\�3�vrU+�!�˚q�ɶ)��o��V�π.�``Z{�9�.�Fh٩�n�:�C(e��f�g��A
�PuP�wx
 LZ�gts����7rv�Z.'oe���M�j����^/��]BOsY��@.qؑ���_~!��qAV�|N9Foe�M쪝��C'��d^��A�S��4�B/��O���5���$W�׵R�D��仗����������xoe��ҝ��s2p�֐]7t�
fQbLɅ^7p9�������0��?��7�a�����{'2���@\�;�A��jmz�>�U�H � ��'���3bbH��!�c�M��g�|I/�W]t�c繌�T��,�L�Hֈ_c�s� LvbJ�5�[�U���f�%� $/�uK��l�o#��8|!T�3Ó{�E��~�!�CDܔޓKD$�UsM���A��Pa
F��v,UU�p���p\��or^#��k%�B�2�}��Ճd=-�u݃H���/X�\cD�-�?�@��ضQ<%��Jb�&6=2�Ǻ��=���������l��iآDO&(m�댯a�r0̯����ƴ§��]*��V���'[��P�����^�qCL��'�B7p�#DݷFd0��
.H&�n�����r �J��]y{�F^ݾ���XL��%�����⌴m4�^O��ƀu�SQOꋟ}.�������z���������w���հ A(�PgF�fY{{Suo�&b�Hh�[h�fln-��_�Y�+����аa�׺䚀,�B�rI�u��J��������_�gϾf���r)��ݬ��
R$N����w@'�T��P����ˣ�;4>���\�Rؾ�[EP�Z[
�7�!���ҸA�Ff�2R��+b E�b���|���z�,���T�sk��W_�=���� j�O�m	&�vY#��,H�C�8��-��b�[Xq�A��mkc����6_ ��{�$��q7g�K.I`���ag]wY�	�i��X���圼�>$# ���uh����N&.v\ΒRh�=�qB��� �[r�o�i��%	�k ���$xռ��:l[W� 0�گV��f��"g�l7�)K������ #x�F��/���wr���i>H񱓻Bwu�`Y���[�F��=4KZ!�p�wF{�!vdO7���.C����f��߱�t];�\����cMxE�6E���Y�0tpw�&��
7���zB'o�^� �����0���{:?O p>YX�Y�h����ή��_�R|����uQ��
�Vmty�5oʤ�7?7'X�e�"�Z��R��y�WOh{�+�����U)��?ӽg�/�!�b�3o�~���ǿ絠
���C���	��QL�����n��J�CY���Q��٭�}}��הnġ����\^��-3�g!��Vo�T�;���ϫ�2.|]���,������ٛ��%�����W����#�Z�ā�:�lW����� 6;�����t:s��B�Z��}�"���YȚO3vCDim/Ɗ�XH�����PP�G����=��׆YH�j�ׁͻF1�ǲ�7�gS�m)������7u��]��R���JkP��bH��b,�i߳��ױݨ)8�j�b�ogo[=�gR�i����ܠP�j/�@��X@ݐǠ �P/�O��ʞ��l��B��pWt�S3�6t(����D�.�5+��޽�^0�~���4l�� {V7z�.Pf�_gg���4�9SO�k2
�uE}|��fF<d�����x�f��J��W2�x��a��h-�&����T5O��i/��]�%�9��:f#��<�����=!+��h���� ��x½|�B�ݿ���o�[��g��Az��G���e u[릞�z6����]�,�1�Ɋ�F�9�4�PLב��4�T�0,yM3�!�9_��uS'�=mxH��c��y�ȅz��dC�W�s�o��A�>e&�u�~�HcEc+��KsUo���d-�@ı��8͏A��=J�G/���U,h��,�S�3R)����}��$��%N��ߢZ�HZdm��1���l��`���@v�u�h�� 3qpI�u�e�<~!{���W����T��������@�Fh�LJA�.Id'��t2��� ���^`��f��QzR�_���Y�;�>��{2������\�)Q,Ƴ�`��r3�dmZ.�S�X�fL�	툪[��@&���X\h��W��/�d�Y�Z��@��%�p�M4rB@���S%����1O�р���9�,
+��}�a<5T;y�P��_�K���x��7jn�6:W�`�ڼx���y#;�fz�"E+���d���R���c���t�#��<�������5�=������S���:�%���N��!YI	N(�5����^3s�{��gxv�^ޟ��n�pk ���������䠸'b�n#���GYV,gK~.[ɂ1.F��,혒H�䞈���!���&O�;	��xt��w��ٙ�?��ƈ�б� �N]��bE�rZ&<���/|�e?nD�Z`�{!	d�.��f7;S{�[��F�V{P%ofÌ���x��o�s��$mЗ�o������Iί��&,��g5Uڬn�)�2X�5��- oe�=�a>��- {))i�;���>'�Zcxj��h�s.^L Do�n/���+p��[YT�73��Ph��L�jiEgp�w�;r���N��bEA�}�S��1�N7�Cp  �-��{Z\b��A�dP�fQ5h��&�^c$SY���R]�S[�U������_Qma��WoL�a��tk��afM�M|��ݸW���Mݗ�.AR!pq��7a7@e=��s��GG'����Z���7���Gu���Sy�^����gT��
����Fpc�ߪ�xv�Vޞ�&��_~)���P�*jj�z(�����k�m|E�QyX�"��c��N���X9�~���ꔢ8s�"Sui$ʹDd������6z
��hl�\ww���'�.�P��!M�|�U5v���b��s�3?�~-7�����@5YEod����)�g�o����\G��w��ˋ+YA�&�g���r�����F{�aw,�ۇ�ea��̎U?Ԉ3Ό�Y�7��K"��b��F.�Ϩ�����
�E��| �Kd�
F�?[�hP{ן<8��_<�|��-���)I���%vU5��r-�ٖƐ�0���݈�����ю�kFVW5��׿��S��F���QpB�B�4W�L.��U��Ny�g�1��wd�Gaʮ5m�5���4��b^r��e�[�&o�j���;����ׅzM��٣G�LB���w�K1�<x���~�B=5��Z<z"O��\ƻ�d�F�����\H�\ˏ�1�ϼ�՟9��g�8���➒֜��F�QQ5�e3Z&d�!�����N����~��hJ�!���E�X��G�3
���Yҏ>~̕���l?�x�!X�є�#4��N���X��w	�.�b�w����K���zb�V	��?�?�I]��n5�[<��!���u���'��C��5���1���' fŭ+G�ײ�w̌�nY�e;NdI.n�Ƽ?G�-�˛3����)i���<�Փ(����cf�#S �������y��1+��u,�C��-W+����]���6b�#˾�=45��v���z�Ø��:�t��X�ao[��o�F=�L��?�g9{w�pd�k��q��@�Z4�z� ��^S<)��X]�e2"h�[�Z#P�����$������,1@��
w�|�g9F�+��x��0�I�Nou���ūԣ���ӧ��WOeg�^�e�g3O�Z��/�؆�P�J�.�{�$�Q7F��܎��KHkK����r��6�@8KcSuvRW;4uŚ�M� �30Q�alɱ�UW�z$�X�|���c���kɟc�<��/E�U�Zal�A:��S���M�	 �V�Y�kŐE� Z��O%*1aA1�D��2v1o7�|�Au�����q��F�d���/��������I7��R^xߠ�4c�}�+6GկI���~!�#�ᱼ{��y`�v���0�d���]���}z%��� ��o�z��o������
��������E����.���-u��@Xɳ�?կ/���'��c!C�!��2YQ��H�c�JFB*z�+��	���w���O�����y0&�԰�(�]Q��g��Ø�o���� ��Z��;p� acz��\�4��<���3��u�0G�Fg�+���#�j�*'^�+6���p}q��H����z�g�R�S?d>��HXC��-�����\����1�D�<�6KgW�2����8�7�)Y�Ðō7Ѱk�[ ��Pfdb�!=�{'����O���G����<y��V�<��|���]^��#�|S�:&A�p�P���	���%�O&rxx(��m_<M?�v�B��Fm���/H�"D���1vN��X�gM�r��,R���C���1s������/r.ײ{�'���_�����z�vj�b6`�r+�hh $+�+@rc�����9�!����Bf�\[zE�!E��?��~Z�y�V���?��?|+S��9�����[Zi�1
Sig/�,�]�{W�����ɉ�����#�pL����X/� ʌ���ӧ��!�U�d����_�M]7���Sh�Jo S���0���G]y��g�/���s���0u
��Zq$�0iA��f �^Z2
s�,�Y�f�U:�����Z�M�Ȕ�q-@a���H9��=0�1ٷ6�����\�x ��~���X�� �W!�-V&�U����֚�����1
/���E�EJa"���Z����F�q4Rhc^bUI"�Ƭ�mi˪Q���J�~��5ъ�Թ�;�9|�'�[�w&��=�i{�@�&+U�$Z��!I��u3q��6�ȕ5����������ӽ�������<?_Sj�62��R'Hc���@?���A��z"�KS��5�&�M'���:�}�ا���@L�\�Խ�\%_ ����LC��r�k��#�#�����z!5h�������
QąL HS��H:�� x�а���@}q,�'�rx��Vְ\�C@�hg��Yj�ڳ$'Ն*%ށx^Y���c0���Ãd��֭�;�ks��%q�)G��4�{��gz��ʃ�����{����3�T,�!�V��Q�����1(;^��Zu-��$�����a<�S!̅a^�
MU�n�,O��P�ҁ������T�ב{���/��y�VxW�;8�޳yJm ��U��N*s��рx%��n��)��S�q_��k�=��#%8s�]��,�\_=��t�{�����<l���?g��w/�򭪉��6/�@�L�u��5��kM�\up�硕~j��q�;���0R���
����I +zy����F���l|��5ݻea�8���t�lr���h9��.d�c�ê�|)׳KV��C�����u���3|y��;��_D}}	f$p_��(�[�Y�d��]WsS����{d��D���rn8V0����"�e(�lNc+,iV�+޵�W�Ʊm�811�gڰ
nP̝��5��j��dU���ў�; #�?�ɩ���CA9�`0�ڴ�.������(�>p|
�mL����U�Z:�`��.W�Q�.����ŵ�~=�ӳ.���ȣ'�塆0�?zz�0�U��y���Cj�����y�6��S{��H;��D����F�Pf� �����QR͓�Tvu�\�o=R3���0��Ǭ�-Rh�B�Ǆ��}�2�7oN��m,0��.H�C�d$W�� ��Y���	�!��r0uIu��h�$�c�Oz%u����(Ԭ���� ����/ƿ��P����WT^_y��� � X���ANX������(k���iM :���.ȁ���������s��/��+N˨4VEQ(���V4.$>�Bm�ݽ @�c���Gr���լ��� �$i���j�L��uCb�G�Q�	c�R̽L�U׮�ޤc�!�-T$T�K��\Zuv��؜
�	����@��G���_���%�7�Q�߼��UT����2)¼��A��4{����r�Q
K�D�qF�v�:�����c��a≜�u����p��d�Z����P��?m�h:~<7�9p<1z�^�`Hqg!|���]'c��l��4�7b_>���!KT��|o@|Ţ%�b�}/�������#K|3��P5'�ٚ[�����[aQ\T��	�O%�#vL�:���l2,��P�n��g��8��&�;����c�Y�vK��;�-y�职z��ّ��aL��������ž��[�>=P���(�2z5��;Â�u{�!�P.//�z"W�z�M�NÈ���kg89����#�s��Af���'������g�a$�� 4A�=[a�`i�xD�j�OM ����2�*�ɽ̾jyI��_��I�5$(�A*I���VT
|��AW��TSr�;���`Dд8�z!�4��-ꋼ�w���M�����U�1̬Ґ� ��U��f���ܿO=~�^ȁzc�vL�tz`X��#� � !�G���G�-RG;�ш����v1�	�ߣW_��Z{�=���;��d׊�a�/�袶�gG�(-w�f`qB@�}2�#��;.'��������ͺ9X�I��-*�I�J�O�� ����?��f����h�ae4���:$mM�3���eO�kh��◿���������o���8([g����k,�+ (�$67Ĉ����e3��Oe2E�sKY>�� J�;"4$O�uն`�������5�䳧�dC$L�u���0�{M��;�j�(��Tm�Os8�O�{{����T_�@U���F%.�����\%+7-Lк4��A0���>��ףJ�l:��4Fv���Ws�i��CfyBtK%bw�)ja��Jo�l���l��N���H�AA+d�@P\q�X+��c�-;�%�^l�]`�	���x��f�Yk����r/_SǕ�Y��.�=�Ϸ=�;A�����B+4�G�8l�:O`�������Gx���YgX���R9"�rzz��y��,VTJ���!Mx]����Ր�������ּl82����<��}��.����z=,������5zz(�(
K�9Zbn�ֲ���3�Q27Yl���Nںc�e������������o������m�a�t>a8�T#�ng��*�!��4�헧g�����M�J���]�}��\Q>qkw[��;�XO��s�̕y�Jc�֝ڳ;#!<2_�6��W���ͮ��'��0�o3ΙAh��`$��5�����	 �B�qG�Ŗz�cL9gvFjx՗�ñ<8�����;���gL���W7_0��E1�Cꛄ�\aBQ��mIok(��-z'�'j��)� c�|���3��m���{F��:l�eR�~�I���p�u�	hef��L"3:�l�뾻�k`�'��Ey�?$!��Ś�aN�=rt�<��M��`���[$��isv5��?���)�j��U�<bn��X!�a?�r*��|F�	�q+�3+�Aʰ�Sh$U�"%�����<�7�B�Ւ�)���x��x��'�
<F��E[�u���&Gu+�� ն�r$� m�u@]�%��2��E�'�(���=]lO>��K=�R��aP�.�������`0��)�?�,�L�ń=`�X�4�Bc�
��hح.=� ��׾��� 1��U��f�Z���[�T'��6��Gf�~�o���j���) ��LPXh���t>��v������������6� a+�JpL�Ҿ="��Y��Tn/�I*��"���jm͖����:Bs��OP��Q�(��vS(���+H�R�����ܘV�oی�q���z�4]$�={"���6L5������^q�LYS^!ς�X!�Y���c�3���vx�VD$�o�>��!Uݬ����iA�*^i6�4�������ն`I�-�l���cDpJ[�ߺkU%����7���%�ގ䪐��&Z6'8�&���j��B�0��a�����H'�7�v�M�fL+6��C�W ��>X�a^\vz�����^	�ĭ���G�,qG�;��{[#)r˒Dp�W[�d[D"���.>�+2l�0�b�'XQV��~F,)a�{�J>�Fp[�Fk��1�gЋ�ZI^�_���l��"�;;lJ�}n�HV�ELLs)že:�IG�O��Cu���S��+W��TcP��K��	�y1�L�h��ejcQ�����&΍���Yf�U�A0E`����$��f���ls��z���+��!�rZ�Cm�D�f\��njgjk���b$���	�d�ټ�����?��� 6F��p��v�����.)ؤUT�����2G��7�a�4��,^��N�����/��p)]���TY��`�Y���f�cwkV?�9�(�9g��?��^~lr~�.?�dD�T�����Y�HE�ɝM���՜U�H{���'x:����c/-���
���eq#W�>�||"^��a�����hn��PY��\��3�q�FZ����ժ �����e&��͎���8��(e�t| ��w=\i����n�p�#��q=��۲lty��މ�&6����:e��E�4Ұ>G$	f��
PK�1��2c�%��fU��gT!g+���h��U��e��^c썼��R q|�.���5z'�D�)Y�ED:���GV�_������2R�Y)�Qj�?�e�i�6��x#)6���1�݅�[G,
G�'0΍Hv�f��<�ku�ʴ�-�����6�h�H��k�	梣�PA�6�4��p���8�3.y��	.)L��r�j��R��n�ߩo����S���u*�] �G 48�/�%���{��z�1�"!y�q9�-�mV�>=�5��D�h�����;e-��:fa�����}3?��:�s,�CCҪdo�sq�9���x׹�~����:νM)�T��^���QY7�`��񞚐3�	��A�;b/���J�cm$5k�v�C|<�ʹ��ƈ�+�dFE�AG�����܂���x�=���'kQ�87�����<��]�u��c���P�R��Ҍ��Jޮ���`����&+�����T3�g����8Jg�fh�P15���*w�C�F$�Y�Q���Q�P��������f�0.U�n Jl�x�ZR��	/��u��ӈ_�ǳ����{����S�1��l���Ҧ���Bcc(�c����%�����-lY�������h�
J�%o���j���Х�l�ih�hź�:��n�#��1,� �%H_v�J�`��Ƽ���-�pVۻi�y4eY�VZ��joB�3:�@/�dX�/��PYV��ݷX�Ǿ����1^{:������]o��W=���씅����0�Q�1��N�oo��3��kd-s,t#���~f���j	-�5s��$Hu���^:��G �tM���&D��pܷ�Ӆ����Ǡ
�������O++���9���
���c�3o]��7vel�,B��ޗ�&f���G��z���M�EH.{e���j�Fh���@�4�?dH�0�&��F�b:�k�,+d���zM�u�1�~�u4�-�R�Λ�"���g洍%������}�����BZC�h�-�&�����c�{_o��<L,� ��<T]s����B���I�#�+�U^K�Z�b��y�=B��0�qR(��1=��k���Y���-`��˳T�w��D.�n���f@�3=Mᅄ��H��)����j�eW���Ї����r��)�Қ!?������yL�����m��+����V���DD�`\�ĈҎ�����zx��d"{޴��?VwcF�f�d�
]����|��(+�/�)��w����'ߤQq̲
�,���P7��/��GP��Q;3�薖t2�-��E�Y��~��{n�;���?�h����b$���6H�b-LܔQ�3o�n%�R��O��y��5)��ѽ���=���G|29�呴�G�;˚����0�S�0	��<~N0�d��;�K)
�%�l8	�U�����]����@虶��,90�������<t}���@�)���U$U��mE�=z٨���F��
2-O��)�/��B��+Y�^Վ�!�ʭ��x����Ra>?�Y$k]Rċ�İ,��S�k��@o�߀1<��K?d�}�c���nm�t�?����@r���"�74��2B��y��z�����j��s�;81��ͤ�.���g�ڣ�_�����Oτ$�$���U�zvZ��<;Um��w�7��G�ȧ3y���aN�Zi��8w�'ݮ;�}PI��ÿ5��m ӎh}F�5>����F��A��?�94�Nݡ���G���� [pK.B�^'c��h����aZ�q�n����;6��ښhUe����֧[�<*�٘����[�,Z3��B����C�t ��!�F�;����[�{Ћ@���(���g1�\
GCt��닫��}��+��.�E�r7�&��~�X�E�j��S��	^�O��tm�O��N�8 � Hr��F���d	�w�o>�����\
 >�1�C&M�<����n}����4i[�������l��O}��
|�\eҀ���Ec ���=���m��N#�N���n-[��Th�
��w�5������{��~��=�����q�k{VZ(�U�I�Ӎ����I&M:�μ��0�x���XI�v��A$���Hf�o�	����p��B4YIM�)�W�W�]�i�����:w0)~fD�r�L�{�㈸NU7!L��7B3���".��L3"E�
��0��4F0,hqI42�1N�6�˺��B�/����H�l�	�Q��~W�%>�e����5��x��_9~�'�G?ߟ��nȏ<��ҁ�|�ϲ���
�ߥ�}�z�A?~�E��	֩��^�N��̼s�!�B�a7Z�֬�Q�%�3U#�@�L�z�Ѩ#_}�P��L�o'2���ߩQy})�}�^Nϯ���ѽ8hBn���r[��|�|�iT���D�:�������'L�rdD�߿c�f��"h�&ZL��+���ӟ|D�$�Un�쾳;b��{H��vr����ll�BE��Ӿ�ۡD�j�>�݈��ӵv�B�p�U垈�f�T!-�A�����"�'�o_G�{�:�uj����&[�2��?������7U�wN[���h�)��������������E�O/��O��c�6��iu�ޒ������G�ýx0l�U��Nnzc����je�"V�M [���)��o.	�qSr� _c��/����������=y�n"����Y����_e��yۑ�!bS��2.��u���������TC#�n�넉 ��3�c�2��� ׾���_0e��;�C#���jW�*.�^;C�2o�Hqqp��N�X��<|{��Eo�XS�F3��^̮$��x?�X���㦍�E���i9�l�������������񅑖�D�:�ƃ
�s3��x=Y{A��}���3փ|�Qן\*�1m�WC>L���̻�3owM��5v�{� ~̴���7��וּv��c��q���x� �{ǽ�q�3h�@q!P��!���dG<>���3���2uK<.�� 
��	b]&E"/��ôCbwH&Vכ��x�o <��>3�89���A@��Ȼ3�&��^�����^�O>����n(/4������ܸ4A��/�xQ��ǉ���o�y�����L����l��0j�$�x4���l�NY�l8�Gb!,{��$$�/���bkD����݋7k�n�8[��č`�m���3��J�<śgy뵑���Ne�(װiP��}0�?v�Tѫ��fo�ʝ�����ּiA��ҽGc��SβJ^����8Fq�ic���״�S�ٻv�;�%@A/� �ԭd0�H���՘��z���z�m}�\��t�cVg�k�B�#>C#6F,f�l�"�^��Hmm}���Od3jS��.fS��R�JVsb3v�DF0g>��CE$��P<��Ӈ1���B��s2���a�,�h����ϧ.͆p	����/z�t����G�
P��s���<;�]�,U�B�Tl1P�Xq�fY���b���z�SYju��N�G)~��p�r�lGWÜ�r�V��1ɳ<�=��n+M��`FЙ�Z9^E�Kg�]��3ظ�@�L��{��S��~"?���U��lzY2�LG���P���	���˜Kݸ��Mʼ]�qF�Q�BJ>�������y�0���m!c#��ڐ�Q7R̔A�Uؚ���o� ^�!��B��!>�K�7��e�2&3]Õ�Z�ꁠ��z`��X���L�m�����C9?��vֳ�f�RYo�[Qc<,�w����쒥eE�*?�:��v�,t��c�"v �{�4CYqQ.fK9?;e��B7pH� �x5Ol	5v��?���ɒ�;73��j�@���X$.ZF��-��������'a�G���_��G8ƚ���=3�X�,�X��(R\�	h���ު�ַ���>����W]U���bUW�%��s����wV����56��B���*G��'��[ȭ���0��L�%���.�v���=l���\W�D��_٬��4���a�4��^�ddH��i�ЅJ+��މ��! �Ȥ%-���#iIѧ/��2����U#e�Se�_*��1��_�lY*C��Sʬ��P��׋�2�THv`-��H�R�#
�H�׺rp��W^�kQ��AH�̴�(�\ɒ}�\S���H?��i������3s���.CU�+tH�R����R�x^tTj�ew�_[�b@Q�ו*�j9���P��DDT��eՂ����M�X���h��9�8��3�4+�4e��e�k���LXL@�����hzdk�NP7�#u"���5./.���$��M�5�-�y��-ӷ)]���H���{��I)Q�� �lPB���qtR�슀�e��Z���u�WE�K�O^�+c1	R8X���>
_@��D"�I���jdC56m��?4[S!)(1�ǁ%��Fa,j�n���O憔5���WA?�i_W�B��zi�Q�������ZMF!��;0�|���I�0�CJŧz`�o[`�&�����∪��$Af���eӴ�Ϊ_����I�"B�0��MY�B�IP�kҹ�2�U
��B��e�o�ܘk�5zi\�
��f���2�g֚�Viu+R��%I:��6��X��+��7��4��p�F�A�� K��X%�x2���8e�b���EK�����
#�b��̔�8���bIQ��Сp�l7 �$�*i�4Z�<��aix�m���˳ƉBx��V�4����	������q�)�~k��*[��±���uު�z#$&*-���3Q��0�	��5�����$��j���W��?�%
�.0ٺv�M��؉��A��3^�Z�F'��	q���z���5�\_7�����5���/4�6��u��	�$];��A�^�CB�V���,�X���4��ûbSQ6n��↸��o(�.���v�bİ�x�nrT.'RI�W��nIA\f����v�� '߅UZ�;��xӧLr,�W=�����+JR��x�5�����;D�9��{�Zs��ZV��.P&*C1bT�)l(�3����0.�2�e
|~~֖�-(��`BE�S�c6T�aR;�!nJ�q.{��w�FP"h=i�S���� �t�%X5W�X"
.��d%��j4�F>�GyD����dmXr?TмM9�D+WQ�M���v"� jA�O`>	�-l���%l�D��@5�#P�ݧ�
y�(��I�p���G�Yq�r;$�Q�F:�gtJ�� ­]�: B��u���|e���i6�*H-(q���k�aǡ��م����(�#��I]�u6Sr�M�K�Qk3��5PB
�����j�nҢ�n@zp�5w@b_jĢ��E��|�P	�:c\X�۝�F�Rom��@箔������~�~�2E��]���gȺB�=	5%O�"*5�=d��נ%h�F���m���p�.+��|(I�h;I+�!���"�p��3�@�;�t:�BFH����o�N32R�4~/�r��%-ϵ��ބ��cb8@�F��EH����K30qs���5�<c���~�B&S�2%�}��wu�B�����{�)�T\�F�����ϥ�1�:����M�9[z.�#�,Uv1����p���#�� �7�B���~����fD�����|)�*�<r}H���k4�1�^[]������ _�X%jnF]����.ď�P��������YED\��@5t�&t�0��igڱ�}3��G�S�K���v.xܵ�g��87���)S&˵�A9Hw2&�yف�?�(��,K����	� o�Dc�®$���Z�X#C�/OF���t1��cS7T�֫-�V]�x���5
�ύ�$�Z@\�m)��L�3m�
�Ftiq�R�YG���@�N��w��R�qN��=�Ï$��N�K	J��9F�
��"WV�:���-(C��۠.��'>�
�$���w�ޕ���Y�Ox������*�r�vŢ��$>����f!�y�p� ks����e�c�~J,�n*��3��2�]8RDy��!��_;ĕ���'kk p^�����iȐ{nQ��kVOeS32��J�1�{o_�G�h���>�~�vXZeyT��(��4�஡��@Q��t����{Q��8����2NV�8�*�T�:���}�r���.?P��J�A9�*���E�0R�-M�ƣQj���2Qv�;�(h����:2n�*pZ�e���-��P�K�b2�� �L��$X����&Ʀ�����i��(���<.�}Vh��oIqj_������%Wc��g�rS��h����˾ļS��;��҆�?�|VVK�[�܎wZsg���&���N�>M�����f�_��+���g;=�"�e�|R!AŞu�ˡ/
��B�Յv˪�e��kc[a�=���-S>d3[�3Ja(�7�˓h�U��]p�^GJ^�%����Ʋ��]�Ȏ,&b�m�m�����C](����0�z&�!Zs�{�Ғ��Q��5GP��	4/���w���B��`eR��<�V0϶��%kT��wJ�y�4����j`�\b͒O��pAB�n5d�-Rx�(-�I�V�=R��Re�P�:�e���)v8GY/�YQ��0�ᇺ���[��2N���ɣ��8��[�0�J1W_�rw$f�FKF��E1�S�16-ɒ!����%3%�����"�:v'�¹2�+�3.7&���ĺ�z<�#�$�F���krX�#Z�[���K���9���7�,�vM8V,���|O���(�pIO���鰶�ei����	�3C�<�Uݲ^�I��Z��2Zw�h�!�f+r2;����k�r�(i4���}�9�A�㕩+{��D��5�z8���m��To�����&���8{��v�{^Y>y������.��*,��i[��4)e`h�C�ܟ�(��gu�A:�^R	��!��N� E�.?���3��+���ݘ��Վ~B��I��	@͈
Ic�3��ד���Ե��Tt�x�6d��v�۬L�3d�4v)���w��V�f��z�e�L��܍A��+ֵ	���Ռ*���i��o����[�ҷRU�Z���r���*�)/:]/6F��:�J�C��<�u>Oӄ�0X-��2"N]/w��B��S�t[6�R����BO�!�Zf��!O��o���)��i��B+X�?��P�jUe��%��=	˟��_V*��q�î�j���z������B(�۷LJSN�����'e��'��r����z$'�hi��qU�'���=��%�\�*w-L�21nh���ٌ_A�n?Ԏ~S�!ɤUk�ԵU&z���F֥y��vd�2*	2S�l^����LM�����TWx�^i�dI�|��'���쭖�W�&��n�숒@�\`m��my#� �&�����^,�B���P�
�Y�Zd�Cs���ڵ���YmeW+��A5#R��t4UZ*����Q�ǜ ȿ-�f�*Є���Y	D"0�:����b����ɂ�R��އ���U$IYS�F�Z!S�0����}�J��R�k4U	�5Xv&�.�3��<�N8�T<�wQ�h�XG��Nx�ɟ�Gy�9�=m�KD~Hk(���W,*Q����<!��B��+�E��cH|���1Jt�DX1���⫰z)wіQO�?��NQ*��Oያ][O_��D48VYk�ԑU��Ѷ����e���MS�˖��
����d�ZTun�|>����Xs��sRX��~NJd�/�
<��ț�E!Бr֡W�)$NcA�傣CBTV�]�hV�ZY�y���u�����5[�_�78��[4��[��G�G������Nd\9�`ǩ�.�f�����?�<�A�!9�����8��'<���I:��ŭ@���J�#=?�D�ARE�IT ��;�j�q".EԈb��lZXk���Ī��m� 4-Г��%٨�?�k&C�<Ւ�>Ĭ����4���E^&wT�����h��G � '�@�k`h!��
;N�vhO�b�g��<�D�bV̤�d��ٖ1�T!A�"�z�BZ���K����C���y�~�`�G���<R��ψY�R�+���%�A@�(JS BʕI��+S�P��v\�N8��hYJ��]�F�#�+�c>��>�}��5�i&c1]\ϣ��Q���Ӂ�1W��X���o|B�D��ֺo#���.�+P�X�V��n�4��epE�S,��)�Z]�6�{gWh;���qQ�m^q�XT�v�I-(��f��<��)e%I�[�Q��h�d���nذ�Z��]Db�N�7N��"�����i:(��v�J��v��KM�
Q,#"�1(�Iu�5U�5>��zJ\C��K�������w^�"��"���!��Ј4�IL�[eA�4��)�h�&�lL$R�����%MQ��c-`w�#䚛�aB���?\y�0������E�:W�7� �h��>^���8�p1Zſ�y����F��0��R�&��i�|��D�P��cM�}�M��A��ͮbͤ�#ZK2�H[M�M&t��w����vvX��iF�/=��Tz�}t������C�ĕb�>8V!�Ҵ�s��Z�X'"L�c�&FC��K����՞�e��8ԟ�s�ŉI����D��$�ј9KQD3��Hi��F��s��5������plhD*�>������ �+3W�V�JU�$�t2��R*��T�@��]�������Ύo�߬=���?�-�����ײ�V�?��@�/�Չ�8�Pa9��I�[�]��
]ܐ} D)�ɒ��[����f��Ja�n\T]������hnl,�:S�e~d8I/��RPEI�b_Z���ڥ�%��"u���o�#4K�1��O�u�A�؅���P���l�����������n�ߧy٢�h������E�22E"�F1pצE��q�-Iw���2�
N�[���d<�n{�.?r��p��d:�m0�V7TV��ӅWj�
*"e�,��DR��@�-r-,"W�e�>|���L|vn0�ea��~��z��T��.52:EM�d&k�ȉ�5*��	\��$�J0�۠�SR��҅����c��s8�QM�(�F���
������A��=�,��h�x�2�Ҩ*E�+ۖ6�r��i�_�U$�^RՅH�@��z\(TU۶/K�j��kjY��5��=|i��gY,��К%���<�@��g?��]Wo��J�D]�N�C���������>�w���ΔM,���6��2b�)S)C^�2V�n�������4�]u������`�<�������p�L��-��3�3���{pf3�|�R�Z�y�NgV�4�O����ʊvM�s��K�:,-1�W��.&��u��� � H���Z��ba���B��T0Kg��ϭ�n?��ǃT�Nu��	�R�Ry5gi��ˑOrY]�)��<N����-`N�"��-]���ˋ�V/�#�=��\���}���{M"z��,������s��^ ��7��5Q&��K����8Ȑ��5z�^���G0�_�&�_�_���2�3|5��_m�u6����l��ikkL{{��*su}Y��� 08-8���"�gxS��m)��~��+dpZ>%���!ŕx
:Bd�u�*ة8V}X;�x4�7�@c�+���X~�h�C�7jpV�HA#��k�Je� u�$xT˯��������B�슬j�V�=C�KشV�E�k���,��[� ������"iaY��]𴚨,^���$9���u��>N~�
'=|;�4TF	xJgt ����z�M����֎pҚ3�(A�P�Q�{�[J��C{�*��6(�3YK?G�|��!w���
XU�UvU�DxQ� �b�F��,iQ��F�]���R:�GKjA�������$���<6����+w����7:A�$ʙ 	�E�4���2!m�l�䕚�<d�)ބ�aggG8<҆��:�[J�g΋ ���*Ҡh���ʔzЂ����Mi��Z��4�tOK	<�`��̯�j�RY�t4f^�����s�\y,��,�4x�ĵ�h�f��Ճ�A�E=t/�k|�5�-%�nprb�4{xm���$^�Ïz6��?��O�����R��e�]Hj�Z�"��J��-r��
���邴��'�j�>����!���_w��wҏb}�lX���3�P�)/�_��3��jW�9��M��8K���Э���D�U�%���`S��tt�>DQ�R�^�%�{�_�� �s�j�漤��B'�|v��~C�MR��{�Qc"2����nUp�TD���S��I�l�M?T	^��[� r�"h\#�&�0eȆ9��NJk�})rB9|��^�v�T�N��k։g��8���*�$5�|*�"׵�GZ��2���楓�?{]y��iU�?������ֹf��xh� ��(<F`����D^{�Z�*�Q}��(����2�i���/X�2�|����'���v&U�NUWK�T��K��Rɕ�֊!%��H5�fSQ�":�]ǳ1u:��X*gTms�7`�]�s��̭=V��ke�7���̤��xd]�ҹ�i�DR���T�\1z�R��6��Rݠ�ŋ�[ظˋ�.��`B���m���Ƚ������t�;䆙��%I"��/��&"/2:d�t�wBg�lХG.
�FY�c�!27�T˶l�
Nn���&�+��\��H+A*�ZC]b�Cb�_I$0
=ǫq]p��/�]0si0��=�c��$�G�-ђ�T����+-��٦��V�&��gj¹����G]��Q�
�?tMV����"���e����r��k���?����eM��3Df�.���J�g:���0�1��`�4�v�BS&0���耿�� c�sC�-)㷞��Q��e�F�.{��P�q9ph	i�e�-p���|�	$(4��̻xIf�¡AL���A�s?��Z3�*��?�b.� ��(E�HJ<U�D,H�Qh��t�^�-�M�*t�-x2���v+iR����F%����B�~%a,_�%uN���FeAe���z\�J���W��v��u�5J����8�Ru�}�tim�U��m��d��zتz�%�Itͨ�)� qiRuZYW�	�X�RZ�Ӵ!��P`��5�"8K)�)~��!�(ێsk�9U�s�꿡٫�3�P|sd�r�/��M�"��#~_Q~���Mx']�>���gZg�^S��Ri=�8�,�~�4�E^�:!GU.*¸g�C�7,]�r�[shP�f��6�Ўd��m
mb�.6�1-^۩T�%qO�����ۑFi��]3��Շ̪�X���h�B��SJ��`8��I��m�G���cw��\F�F�����t���u�I��E�3�W�V)&�-C����(���g�$6�P�E?+~H�<�,����5�C�.�NK�e��I���$�/#t�k��Bw����˒x�~x��5���j�R��俊uS2?5��u����q@b4��H<Ъ�A�q*������_.��ƚ:Q,^�"b��iqY07���誕�V�)OkbC�2�Y�{��:m-f�WD��V2f�L��D� ����A i5��� "�\�'q��Zg���� �I��|l��GC�'��uǂe�����FK��b�'�!�H)��m*�p������!��kÖ� B�W�H��H.��b<��,�ZJż��JK���Cblp�E�r+.<%�7yq�W�V��	f���_i��U�-�n�����Q�3U���Έ6����aJa���m���:�ܭp�&��_�D?4��L�z�k����M��gBM(�ht��Z��j�!��X��� ��2V��<-*�+�M���f)��ɚ�W�H�py?GDb�������I	t�-�ǂV�"��ku+Yg����5��[�l����R�y��b�j�nG&͂X��&�%�;�ҏQV(��+��-3{C-0�i����@����	�g�Y?��<���iA���%k�K�2�����34Q!]T��O+B��rOx�N��#UZ�cKs� ܋��^ �3��`�	z��R����+�X��G}����ڊ��K���[
1:RD�bX)�ч2�D��D3��jCR��g�tz���|��KV��\��5���D��,ȃ�e����k#������e}\-��������I��V�\�\�G�y$���ϟ��pJ��ޓ4�r(ms�N�o*���*�{�dC�T(g��B=�jpKRFl�:]�!oH�z�U�����F�e:-�F��N�5ySK�>$H4��6LH��A���R� �A�P[����}��;vߢ���7���cv��G�U}���82f��X�d�Ln��O�Z�2J�Y��װX��$�r%�*3Aq��z@����$T�Z����:��ьY���qYE)te��Å��&!�b�ԗ���P�l �Ƣ��evo�JMɽ�ʴ;H$�����~3�5��Q����`c+�	�q������D2�U���偮����dτ)_�Z��@�7�q�@[}u�&�	{�:��KnnoJK���� �ѳp��`�ʧ�~Bx<��`Ȋ��ghúsWio?���#6�@K���(h����m����
�B�q���|X��H��+vғ��A�)�Rؤ!ݖ���=�$\��*��7?Y��TȤ7��Ċz���Ϛ+Y,�)=�dVR�ʴ����ht�;Ӿ��0~jݺ)8[�ơ����{Rh��ZXRe:V��F����+�(�b������M����'��E!�O����L}{41jK��.�"Y��Ù�pP�t���R@KU�*%-΢���6�I�s#&��\�H`�j`0�)�j��sA9d����A��
f:��B5Au�'���g>-c�JLqAI"���٦�������x�ַG+����Q��S���6ap0�V�QD��pi��N{�>ub��#F�SٓiQ��t�1�*�v�j�)��*�F3���=#�{�)3�C�7�VO�Q�X�5��gK��_5��2�l�ß��T�@���gFe���Z1/'4a#��CS��c)қ��"�[�%����Wߡ����zN�K�q8VV\���ZQOn���V�e.����zlmm�d�#��e��x>���<`u!�G ��V�+�+5��E]�D&3�\����al\5�F���#��.zڒ�v��\_�T-f�`�`�M}ˉd�<Z�MwXm�c�*ZPn��h��V<��R��IĴ����L�\�}J�.�z���'���a}��M��X�>�zc2!��A�Y��6*1�u/�Il�0��� ȍua�K�eh��Ue�����s6k|$�R1�l @�x@e��w�^pC�F�`�1�u[�	.F����Y�](��-�{o�R����`��h�'w��I4ږ{��V�P���M�P�ڠ��ca�o>I���w�����O�F�
c�}��:�򃭭�t���p���BQ9�~�����ؐ��G�zr�=���*�(¦���H�K���(�����Ve	��"q� ��E�kJ%F���.Tnp�������"���}��`_ZC�,hr��*��+��	�����e�|<>Wx\���q���D� ���UoR��^<�@oJ����g:�`�[w��Ic��Lס����kŠ�<Bl�j�?�̪�yL$��7�!x5������ٌ6VsR���howO�t�#L�uv/�����m����$S��F�Y$�ٜ|tE=��5P �&�`�h�b8D���lτ�Nb8(��F�F�+�M��<jp���RB@� �9?��]���Z�UcWQ
�/�	yS��:��	�^f�����Y7|��Z��%�u����q����C��D\����GA+��ӎ0�AF4���M�,���>�6�1��J�vy���V�d- ��{}0�g�<�Gݦ��;�����9K��&���aq]�N�&l@�+TS��YT�I�݉�o�.��{�4�Ġ�J�O�l�uX�Nkb��4p�1�=˾1���J��� �䈕H�B�lgPe�Y&�l+б+���`#���K��jPļ�Ё+���G�bpYq>,\bAm<|�t��g��r�����'��ؾ��_�2'q��3��&zM���<^����2�NS�h`.�+)��,��\o&H�Su�����P 0����bL���j��,᝻w���{4d!�a��t|8 �S`�X��ӛ,p٘5���$�<h��ć���Y�� � *[��6J�*��g�I��C»ߤN��}��Nw���������v�O����x�=N�}Djq��t]�����t�]���2�������> (la�
��b.�������N�]j=�Y��y񷹐?'�ըR���{:OH�&I���iPLBv�{���0v;����2t)��'mE�1H^թ����y���4�W��"K=c�����Kj:��]�( �~�}Y��:JEje�dR�jJY�X -x+q*�g`�G�dɲl(�y��51�^��X�Tj+H���%�-.�����쌒��l�Ca�St�O�F:1s2l��Lt�����e�Rݦ���Uz:O�N��d"o�n��NIh��3��>y�9�vd�E��rޔ��bg��@pgk@���~����v�������x1�J�-y�Y@��<�k���Iz@�l*�P���E%@U���G�"x7����Գ*C�7k��+�����wߗ���+2�,�����M:�~�6������t��.��:�dS-Q�ǘH7RE����T�L3Q�����Jы��Ã��u�N4.X����b-M�M0�-l��Df�\�2`f �2j4�{F
i�D��f���~��	\S���c������Dڭez����6)~��* ��T�����
���nM�]��E���r��(�61~9TY8��`.OY]�t��' ��e���@H�QlH*8M<�_��U1ťl�e�J�HI�)�*�-��3ֲ���X�Z��k�dܩ�W+w���v��uŭx%�qP#ba9.E:k�G@%	q2Ya�\=#M�����{eYC\��tP��$��ڒ]��-^��JW�`�DZ�T�؃�xGV��	�>Iԝ
����CVZ���Y���DVϡJ/b���LHY�ݝ=y�˗��/|�g����?�wg{�?fH�.Ч�~��\�H�w���m�'�����P4���J��[9\�V���`s�XT�]A�Ź��1������vd:r�����%p�P�~��&ֳ<�Υe�c��]����G�JhQݏ_�(��ǫ�BJ�
�k��f�L�������RO�S��"����F2є�{�L1�$W6�@�=�6��ҟ�k+�v6$��0��0��E�|b�0��i�biO��$:E+��3���#�;]���Y�>�R�T��Ă@R�f��(���&ҿ�Ȭ�?����J�;���Z��3�ه��4�u$#ӌS�1A���vl�;=0�>]�	8�OD2+R�l��H���RwU|������e� �K?�]8�J�\>G�^�>�1�z�ӟ�g�}�>��E����t�����0Z��c��eR�վ��
K�~/��!�r��{BJC�`����d����C
+��(-�B�PYV^w�j"�T8k�[;t�X�\!Vʯ�4J��	�T���~(����P��a%��BUm��"%��,̴�zV��%��t�I��)�@���z;B�ښ��^����T��$���dec�Rq��/�����,�-i�.��2W'3ɲF��/Ԡ��vA�E���;��:2��D7Z�坶G.�E�$57S����M:z�n�7�1b�܄Pپ��/�4���Hƃ$��8	#5Mc��c���"FϏ; �m�"u��R6Q�Б���DI5�,l��1��7�I_�����St�˴�Ѣ�����cOЃ�!}����nk*iI�	���$�j�[TV��Oot������T�F#���D�/�iM*K� �K�x���^���,��R��j�a��H�)��Z��T�:aCD�VeY�w�W</�<ʤk���q�\_�w?�X�ݰ�rH].�x�����H�Xz��$�O�s<�/ڰZs�jJ�jʥn ���󵐑L�ں��^�k�T����j^�uu�����Y�����"����US���փ9u���p���������(�UUІ�07�h,��S��+t��˴s[�6:�5㵝J&'�Qj�`��^�����_%BԬ��2�u,�	�1�"rk)�(��+r��(�@*H	%!`���7��[�g�]��~�F%�����ׇt�'���֧v֦�xD�F����'C��f�QW*�� }h�S�iZ�3��L-�g�en`�;l�\��Zծ��g&�N��R�>��J�k��]Z�zQ�3"L4�R�b(�b"3w#^G��a�#��"��q^i.���p!� ��&�����I��С6�zZUc�޹�.����q�'����D�e�]rD�����a��ŏ3o@*��ܠ�0DZ-�W1�tX���T���٭�D@�s��ud�՞u�S{�����I�+s"+9P�٩RLH�J�_�Э�w�����V�-Х�.�	�=��B�o撡��g ��h��mD�O6>?��@��6_�����������[}�Ib�������s��S�m�{pG�D�{S~N���UQ>�,F:iL+8�tm��vH�,jǭ���m�ۯ��4�A[�%�v,$���%Ή���5�Unh�M��A�=t�����y�Yż����`{���w����h,|��f���N�r��*�c*)��E�QC�⌮��_�:���h��e�I��^ڟPۯ����xm�PJ���>���Dj{����K@V��'b Ϟ9�Ef5��z3�+���HP&������Liko��_V�V��	�C��O�?"�`�;[F�f����� U����}o�:i��y@�XJ�n��P"���D �H��V[���B7����(�\���kH��*�H�A�#؜4:4Ї7����(��"�)mf�m��465%P�r��e��q��Mm��/���.$��w�#���Id폱����z+���D]b2�;�5�f�����a�!D��0���9�=st%YAg0Wa	��kHwQ�	���JL![W5�b�k��S�-��$&�U��8���-{�$I���1�`�u�~}�52Pƺ�j�Nѱ��r�P5�����b��QU�\B͕�2P+m�=X�;�d��V�#�<B�ɂ��݌9~��hJ.�^�ڭ��%���JO�ˊ�*,iy_D=�8�4���:����P(�(�qA���}-
o���0I/�?���X���I���� E��"�9���Qf5�,l�@J͞dvF�@�dU>3��B�X,�Y@�%'-�E%5��%Բ3�~�JX�d��I܍��7R�-<'W�������V�t��JEa��E���J�����}�vY���Z�T�!��l|�á��i&G[v<f�]+ ���yT|i�-�j���`�Kd�J!�Nm�����l\?��V��2F��m?�q��Ȑ�\�yR�b�£K2Z�"����F�����ƣ9��k��	��z4Y�=D��U`��*�2����2S�q��B��2xDf����ڵڦ�;�B�Δ@e�N��R-�IB��V��>D�t1���ڦ�J��_"d��'DD�ju:N ��C!�� �E,�u�XEh��Ҟ�VKa��@�2�\�KQ�0K�o�o�u�*�tx��<]��9�H�����[$��@�Vө�=�c��G3��`m��Z1��`DQ��:Ѡ�(�Z�)��|H���YP?���i.�-B�H5��Jw����2������z�Hn�L��9��T4m�(�M��:�@=�h)J�(�t�!�JǮ� Zo��9�ǊM���Ί9M�cVcF��J��5�T���7F p�?�[�����T����&'��)ă�g:nW�P��H��Y��d����#$�8��6�mY[�X$�P�m(-�־�c����ؿ�]������R5�Ȯ�b�D˞K˿{���F�J�e�Z�ݺ�~�{2����-{���tI@�
����`(�Hek� ��RћX�tiT�U��OkǫZ�E���ׅ�s{9����\�C�̥��+~`�u��$��1RRr�K�^�8����ʸ׼�2E�ww1�I���
��������r2SJ�x䤃�B�W�\��kN2e�<"J�(��X���>h���f��w�����5�L�T��6�\���k��4�	M�d��W� �.�rD��^!�*��ò+�7��p,�70�Y7�/�Q�<�{%�U�y�iQ/�+��f�����[�z�o�}��&+X��4ұ�*$���4�*1M���স'�27��,+Wĳe܏��3����O���.��yh}A��*�����?�{�+B��J�#��H�M&��,AJC��>�w���C�+>l�#�(g��>fM3��}@i�z0)s��2���GuZnHxS�ȮG�1ŁNfg;j��k����w��~.)��mx������}=�����ϓXS���c��m��=��U/T�L���g�ߣ.P�3Ҋ6I�ǕT��t�f�<��V^n,��{j��[����k���hT ��ayu�]��//�_�ށ��c�1n�?ɝ��ćL=ƲCJS�BЫH��$DAA��R�TX�Y�&�����Uȭ��k>-��u��a��O{��a�|�&}X��T�kP�����X�7�~�
�P)��^�n�z�.�>��9M'cZ����#)�{�#XÅp�}c]F�G�/�:H��f�>�n[p�t�iu�i��BS����)� ג!~b(���ȑ���8��H��0;v�S����
\�����ֿ.�n�E4熈�ca�b!%@VR����-CK�B�<k5lXxBUL$8����Up	L&��.� �`G�>����Mc"ѝ�2
]�2!*�jB�A�?BL��Гn
ě���7��@�F�����	����	K�衝��Bb?�
d���i���>G�l��?�6dJn$��@,��̲��x��7�@UJ�������Wo�N|]ޡ0���vk��&8{��x�t�V�>dثVk���@�������9+�i�9�$��J�QS"T��_^���	�,^��k��L�.絍�E�Fg8i���f��j��"�Iu(FFM�A�7Ͳ�h(���V�WX���"�<";#3cwXPY8� ��e0��eK3_A�h����Y�To����x��S�
���k��tH��|Bik�:���Х lI��jV�`-�	\�j4W����Rf	U"�`���~�B*�߅��G�sXx�Ȉ�Z�s>\V�K��k�p(��j�s(��P���.,Q^M��Mp����"
Tʀ���䃵˂ ")��
S��}
ʁ�A*kc��` y +р��$P�_.0a}&,]��N��@�R��ma&3It6	����h�V0t��z��{�5A2�?��x	y�V�S	��JS���a
Z��s���Ҽ�_��	�(����(@> IN��X U�C��+`~V C)b����f7̄k�������J2�<��	=r�=��%����t@(��!��D�RK�c��߯ðܽ(�tv.G�ڒ�g���A�~Ȳ��)�������
T�&H�0J{N�=C�<v^�����,� =h8`���$�56x(�����=����2H��h<��?����i:�p��8h��$m9�^"].�%�,B�8"O~h�v!q�T�ObW�J1�յR/�BԖ�.0�l�z�R@C��9������P"���:����u2��v���-f�����{8� ��Y�tґ�c�r��/�.�x��j���2�\�\X�6J|[(���8������ܰAf�����%|p���t/�Ԡ���4�M-�G�^�a=<���� @��bVh��0͕�z�7���/i6���a�x��Z�|�y�(^Sa�����n	IN*��BD��	�یmSj7��������0�(E������+�D�V���|�XPڐa��l��XmW&�'�A^��ېυ�O�V�wHź�xO�R8ܔ���a*ŀ�4I�r�Do�~
m-����ayy汋����}��gx����h��6�,��B�Ӑ�G�&H��.(�u�7�R.�p�U��0��B�V2���{��;�y����"E<�! �C��ޢϿ�,��W>OW�8'��%�j�9Ș���W,f�p�6�(��H9c{�~�C�߱�O%� ������N�?������WY.Y����h�X���NsAe�^<S����CN�KU�JAI6xh4�&f�fb	FK��L(�w!"
��4�VƫEN�6k�oh
4���В�.�V,���D���;
�t$�	X�:�qk��dL�b������_X��j�f�����l$c�C����ϩ��X�r�_�-�������E��̙Ӣd��v�Z777�LNh4b���P����������xJw�������R��"En�
_�=��e��Z��Z�]��A�]8���[0jhw�������MFt��iZ�u���;³�h� j�z���m꯬R��I�!_��._�͛w��h��y��o+��N��OK�D�I�PyR����!�᱔i��i&͎�DS�b�aŲ�"մ�]H�@-o3�S�S(�D.�k�(�+�Y�NᣅFC�/`���K�����K/~�׬/��>kð1*M���N ȴ�o�?�zɼP�� \J��VW	59B��Z?}��Mv�"\Ē!�.t��mJ��}�˿�_��ߏyJ1�s�1t���ӭ������0�ʽ�W�B�
�e�e��d���R1���t�A/�>��7�d���S��"z�z�*�P�RGz;�`C�V��
�B�E�8yޗ�s�-���Q�+��BU��l>�7#6"��=��P�Ж��Bֽ����L�,X�<�@ra5SFw�E��W�|A�KJ�anP*
$X���~w��/t&��'�HK`(����� �D�m�3M�z���苯�LΝ�w��K;���?���f<^�S�N�´�/�x��yY���}Z[[�瀁���2�^���׿�������x.j��k0NK�a�����hө�>}�g�g��m��h�5J����=���<}�ÄƳ+��4��1�\��1_�xVbǹO�2i}����۴��uF�-��>�!�LB �8����T*���B�$=����+_V&�u��΂e����E�/�Gl�M�M� �����!<մ+*��(��q)�em��5�Ҷ��_}�>��s�n��mL7>�Kۻ���o�.ԚÜ�1C��zT�s#M��g��>8 ��P�V��u�}r�}��@7o=c�|�J\�T�!X��$�ݽ1��_����P���v��#F20�B��DGH���E�IɆbLm6R�N��:���K+֕v�>��%:�ާ�z�V�|�1>��O1�!@U�������V5��baV� ��e�����_���
�*��F��]K�b���ǢO� �Z���i��9���첑��!��g*� ہukH��?X`�&~��\��"h���Z*��b+X�#�$̕��	1 hkFD}D���
?v��ǿ���g?%���}ʧ/��s�S�b.���EA�:zWĝa��m��
�]���.66��Ik z�SWhc����}�;���W5��F��o�7��g���~�W���6��{lQ�et���:)���a�@�|���/��P" ��;=��w0�9N�D*H�N�ҵ�5�vg�~��M�'�K!���k��`�a�U ��1a��CD6���y.\1Z���(2��Hq�M��{����7�M9�+Z���� �lŧFC~�9�Y9��-q;Q�5�2:�{���l5��i�õ�0��2��U��X��~�߷E���՟�)}�?@����@-^�{3;@�;����PYFc@��vW*4�4Լ��g]6t���X���9��kww@������ݟ~�e0�$PCb�0%a2��a�2��ø�_	��d>�V�C����- <��k�X^>{�~��|�~�K/��BZn���&�*0ˑԒ!��zpX�ׅ�{�eD5�9ަP��J�Vf3�J��3g��b洽7��R$"�C�U��f�rՎmJZ<_��T"�����!�PR|�L�abA[[��fZ�ZW >h���9�C��C��NX �}�pa�^�����?!}6���z���/��"蘂��H���AA*P��X��	b,��(�W����G� �������F8j�?��˹(-Nw���
n0٣W�|��}�Iz��ρÞ׮Oi�%լC�N����+�F�b�;�`�\;��X�~g��̈́��1m���ߜ҄���_���.H�d{�?d���E˦��X`�:�P��ʘ�D�"�Q3�u*K���Ou闿�E^����u��^��Ya���<4�X�@Y9ޥv���=I_x�z����*�J�R?�6+��^�K��7�O�+�2�
^S ��]��|�{��;sV���oн�}
�txK���TH���
F-;�zJ�1s����C����@��UL����)����`�ЏV�J$���\�����Q$oM�5�q,��|W���d��������:���`�5�O�X�>�M?�ʋ���� ��ֆ�k�X>`�3�u��	�CyQ+$Q�	v5��	�%�z��j�NDw&vS���;3~)v&UZ,$KL�2e3�R����:,��ǂh���y��B�C�Ɣ,���pQ�$]a	�
FIT,$ց�o3Xak�0��"�+u+�����;H�4ׅ8w�]{�)�t�B)c�֮�\W���.��y�z-���#���"8ˎ����
�����X��
���v�-�o�K����_}Cf�H#����|�ۋ=��	�護h�z�;t�]Xւ��]�[�n��}�y�p��]�p�����xN�=������P��N���"=u�,hje�A����Ɗa*��ů7%�%ݚ�\��jk�s[	~U���'�e�Y,c9x�_�[_����:�m4��������{��r��sL�G��x9�g�z���o�
������as'��(
��x�=Ɗ��|��؝�zz����\���?��ʳ%e��4��X��J=�},A;�[�e�TG�p�c?`Fz��k�!�O'Iő*�->��*��CMwgV_%z&Y[�6I �`}5n�8���!�7/g2�6�{D҂�+R�C�G���Y�����抸��,�zk��?<
R��S���0h��$ҺD� ��՘�&�4��ȞD���x �&o|���1�5��D�p����ڂUB���#�@k�Qy���!#��%lҙ�5��T�E[�[4BS���#�C���PF6S���nSF H�ic^��{�ZE2M�9e��ȣ���kO���:�eo�uhc}��޾O��_�1}�`������grOR���XDL�
��B�Fk?溲�3�ɇ|��?��/w��$1M/�^��p#���_^��Dk�$ 9K4�\<���J:w6zX-vUF�dG:�T�6����Y���z��&#�Q� ?Fpe>�!VNK ��-�iH, )�v㼵��E,�W�T�4P�Lk+V�DW٥[_�K��M_O��eCq�������/~F&�m1r@m0>����!]��9{�,�H_mK��d���#8�Fu[`��jj%�tx�2��ߵD��Yj<��̦�5Kl�5#�n��(�"��6�|�Z�YS!U���@F����d7/$�҅��h8�kj��FK�J�A��8ę��h4��m��sq�JV���:�gsQb�_ ^\Ĕ�r��5-fu�EJU�iTue������Ae�C��)�)꯷�h�֑Y�k��\��V�J��h�P�h�C�J|�&�i߄�JC!b_�~�BH�%��R7a-[���L���=I���_�3�}���l�Ft��-�������ݹ�W��dA������/1��mVd~VO���9c��v�)�}��7h�����;���闤x��oH��{���|���w�@�� I+�h\��+����3�uXS`��P����O�n �O>q~JC���.L���vKBG�x}&�1�&�fH��,r������u5��rm[��2��=�uX��}�[��ƿ�3���MFw�q�>��=`�܉��"�Q�jp��`�,:�U_����!�+�ѕk��J��{����ñ�����YnZ���K/�~�"�0g4��?x������d@~�w�.���5^�u]A�d�\�&� (��+z���X�0����T�k7��i�5FH7���a�bG�Y�c	��A^�	%D+�׊?B�Fc�t�����ϮL��d��P2|I9����B�/ϵPK(9-�4��z����X�S���=vu�(a��KRD^��)�  B��E���`9UE}�)�����u�b�e��T�c���ȯ[9��(:�wp��ef3dV`M�*"�>����vG�V����f��RDd����M�����z3����_�_g����cmE>���lH�����ޥ��_�	}t����R�����7����|�������滬��R�1���s�_���n�Y�'�����a%q����^~�V7z��m�O=�����;�$.�ɚ쯓���f-5��g�92��3 /���sd2s!5 �x�@ԗ��o�"U"H��_F�zL�`��������Bpp�u�JV&I�f����a�4�A_��}>��;��Ν;|螢��}�.�|2�@uF5v."7j���{-8S�PjC� ��/	�-f�K*S
�̒I0��W^��s����xo�d���������������,�/_�g1�Z���I�DhJ,V�*�[������1F��Pc1���k�L��wEadPX��qʹ��8��h0�Z�����%��!S���**%��c�������>�?��A��;���s�=#F�7�5М��`$k�j�V-����2A��5�'���Ϲt�]|�=��S��&}��?�����G�O$�a���w�`�k�Ο�a�Gl4��b�����D�z�̀�$?����W4��W�~W��U�"զ�Xw��1���w����r���+K:B������گ�m����ߣ���T���[�nҗ��Y:��e8ۧ���z냛���W���?�ڦӛ��ܣ���/�m߹M�>M�+�/}���⧟��|��Oӿ��?���wiu��ɤ��k�
�+�^?��EC���Ι׭@�O��74� ��POQ1�bB`S�A`�#��I�Raһը��`c$F��K�Q>���٢#uwa&YN��V�fE)H�6�m��~�X��9�Y��X�{�f�9���b���w��^_F�����ӱ��Xj��A�9�A�k�
j,& T���p0��%�*h��N�7�R\�n�E�G���x�:u���h1����[w���S�b��=1�z� �nC�͙����iW�� qMpa)g������2���&�>�������&�cM��� �L�6b5��� ��X�W>�z���i1ڦ�H�FAO_��nـn����w#����X��(�کȇ��=�t��W�=�\Mh���Ͻ��r�y~�	��׿#׮�$J���T�L�ϛq_�fU?Ɏ$(���t(�:���*bū�T*r�7P�9��Q!������-I��h���hj7Ɣ)XfX��e9CZ.�����J��F������^��������������?�G�Aמz�DI�]�}��?����M)?��}���׾D_����W@���cI��V0�RH��m������t�B>�O��[�>�O�o~�pq@͵M���p��Y3K��iw4��VL�S��d��)z�^C�E�� �����)z����	<�L�$S%�Qx �	���p�{�"�yn�ۖ�}X�F�� �zv���砕�3�^ݤ6�[:?��ו
��MUT���&\V�$�Q<��]�%�h�IR������Pjw����@Ej�ݾ2cw�����ެ3z6�����/����)��!��"�������S�����X��*�Y_�wo:���O[�R�9d����&�2X�.��YF<@�R���f�1�T���5u{�}�C�HZ$���uN�R�Ϩq$�X������v]����_�9�5{���#�7^�Ϩ��v�C�Ncꭤ�z;
ﳦN`k�t3���CY��Z2�y1�㏜�����%��+��(<�V0��Ʊ�N�U���3�xXw=U($,�M�B�&8��o�b:J�3x����%��l���2l?x@{{3�}P��BK����GF�&�0d;�S ����O]�@X�פ�|�5�/������x�����?���R�ߧ��?�mz��S�c{��|�����������_z�N�=�J�s���|��7d��+�$��z}�+�\Ã��Ōy���Bz@+�>+����f�	+��� ��>Kfr�����V_���A++}�@�a���>+�T�21���y���F`�mbm�Y��sa�J���#�~����%��H|tF&p|��:��uh�Y�աY٧�u���/�pg�@:NS��}��/L�Q�,�ZձQ��$s��wL�Dr��$Z!�"���N���'w���)>��`@Ü���nbs]���@���ҕ'����o}�{��Hb�K|ό�XQ����[��W^�	�%�ck���}*X^0�غ��5ư����v���ح^Y_�'�=AϯӽO�����?�ˌ�E�w���U)u0�S�U�A����K����"�WN������nX��P���-���L�G�����ݻ�nΓt����hc�O/��9)����uzxcҦ�l��k�,#]q�ڍm�¿��5FӯH���o��{?`T~�n?IVR�iK��� �"6���X� �:��3(ݕJiԺ�#��PY���Y�ڕH��`I��?C"(jBP��7�?)bsSb�1�baiB���}ѐÊm���nh.�`�
�>������������ҭ���Y�w���g�e�}�V�X����Ux���������K�$���*�2`l���h�ז�m�d��%�+�bTO��+���NO_y�N���ƛ�w��o��T��z!��v�6R��W�\y\b!���[۴� �ҼH��Z�&D>^R`��*F:��a��+�U*Z��\8}�?c�V�[��v���"�u�	|�&uzk��ަSgV�٫����4������ߥwo�+���{�|/�vw��5+Yq��Ű�F@�]�Z��։-��¸�_"��1���|�����#�����u�51>�6O��/�,�34.��5�N���[��9�O����.��p�Wh��Q�}�J�l K2��I�|z+k�[]cٓ�wS�������/�k�[t���|�]Գ���I��R�e���0�C1a�ݭ�>���W~����/Ӈ�����џP�O����u��֫����UZ�ؔv��v'��ʻ	��鉫��L���ޑ֍ ��2���]Zm��
����Y��|�E:u�4���t�'7�=>w�����i0DBg*����nL�����iũQm�f�<���z��%�[Z�=��<��Z-6s�B[�4D0J�cK�6-lZ�v��f]����[P��;�V��.<@0�ņWa}s��͇e��نlp��wcʖ���]��3�l�\�v�n�ݡ�����+����+O_�rC�-��
�,��!��{��NP���.��b$��,K�#2��W�#}�~�|�(�O/^����84�6��g�ң�]b(:�[�;�a���g[G(� ��Tb�;�Y?��
�U!͌��N$#�n��Q���<��;�����]�6ݹs۪���˄
�&�>+�'��F/��%z0DIy�����������=�O���J��}��lcQ-�ŐGm0�)��̋T�����`t���Ξ9ǖ���
�Ev�|H#�nȈ��.t^;��>�w�Q��2(�A�e���׶N��RjA�9�i!��;�I[Q���NRH�,���9}t�=u�<}�ӟe��{_� \���W>E�6N���.��P,�+�/0���������o���-:���qؓ1#띳���	ݾ�1��[������q>���1ݿ�M��6=v�"=��� �n�|#]Fh�x�}�F,s�����W���Kt�]�[���3�2) �s��m�	���鍧#�Z�38��n�z�}M���T�(D)D�s��PDU|�(�^��OWf@�*�����&����7+bpE��u �0n�� U��TʿE���Rڑ������(*c_q�3&ī�,��կҏ_�~���F+���>/�C�9]��m��
V&d̊&M��^�~��|�c��W����e�t��M������e����n��F��O'�4F	r�h��v��ak�9>`4��l���f�0�t��h.[a�ʕ����GX1��<u�	z�܇t�Ï� �+�]�X�"�pQZ�!���|�]���P���>����E9�	k>R�ۥ�6��(���;��O2�@kA.>��޾tw:�t��eF,֗���|_�d��`�3���ⅲ+�~Z4�+�|lyg��q�����L�ϔJ JH�X*�F� qZ����%l�[y_���.欰y�d�4G3qM�cd_�m�Y����(��iZ9Gk�(2A�x�"���y� �ltX^2��Nh��{�t�{�嗟�������ߠ�JA�~��x��c�[��h���?��N��g,@{[9����"��mz��R'$Ty������γ[�O�m���r������	���N6W���^{��h�[�$4_�9F󛼯��O�{�ߧ��l(V��>O�>zY��	���m�'RE�e���ga=Fڼ��J��t�,r�ņ4��&C�yI+V+�YS��͂#N��m����]��R;�i����}��e�n2�%Z�]��*��*t������P�0cT�>8���B��Mħ�A�˖t�akwH�=�i��~��hr���~!n��O\���=&Ux��m��~Ҥ�a!���F#j�sZ�z��|�E�d����*b��1>Pl�R&e�ht���_��4��l2�~��6�پO�A���p�ۡ�fG,���<B�Ξ��^�������?~]�X�^�FW�>���(�/}��,����o�������ˌf���xL����Ͼ�]�~��/^��Oh��	A�n�ɨd(���Q���6V���i	�=�C����J���Xʻ��pp�f2���Rh���4k'1�QD ����K�U��K�Kbd2�b�	��~���g녢�n���@:sR��L��̴���$ ��f���bړ���@mG�!��,��IzRd�A���,��e��I�� @����>uX�^a�?���oӽ{��,��~�)nB�������y�͟Ig|  ��IDAT��F���9�ˌ�[|P!f/70�s)�{�]����.�#�Q�:\r��B�0����B�]Fh���<r��>y���5];���lp�V���۴{�i����_G֬��z9K��{�V"v2__[���b":SY�ϝ� �U�R���FO�J1;�o
����Nqg�P�MD6��@����}̪@C݈-�d1��Ҙ��OX�߸�M���'��/�,}.o��!�;}��}�9:�v�n}p�ݓ��k2"��)���=z��t��cT�4�ҳ�\�+W�����O-�8!���5f!o
�Z���(���/�����������L��{/}fy�]ӵ(�o���-i��9;;;�w����{�9;sV+�32-����mؖށ  ��`
��g��q#��e@��޳	�J���E܈�qC.P��SG�x��p��I���a����)���)�p��7����W4)Z)��j���$�P�Ǝ#sW�쵲���޷{7._��S�O)���_�%|�K���� ѫ����k����k:�Yl޼�*�V���7���:T����i�yQ��(:�n����ql� %6��Zi~T��x>��]����kzeT��~�
�?+t�B��s�k�lG[��60W]�~ ��4ٖ���$�gv�aK�-�T�؛�S�c�����9��\�9�cc#r�ƵJB�Q�yI�c�.^��`�KK����;�^f���
9�U�q����b����>ec'��Z�9a�Ed��\U�'�1���"(��|�����d�m܊v2$��W�Ʀň)ö^coQ��1�V��213�a8���V�nQd��ϻ2��܄���������~(�5��Ȣ$J9"?�ԅ��a����"C��^@W|�v��(_>�3c�M.ɨ�J[ރtp���d�������~�]~S w��y�#ذy#&ĳ�m�ͥ[x�����7OanAާ��H%�@��};'��_�e�O�Z��44�<~fۗ�M�eU���]��F����شy+r�ḱH������lGiLz��a��U�c�sK,7095��fii^7SV����u��5jk�^�����"�VWΟ;���'5&�x�Ļ�,a��<{����䤄V+6��DCbX&�Ʊ"�Ei�&�@*C�b��2ʦ$ZP�Y@^I^~^��4h)�T"�jbP�Y�-��\83@��������M���^��В��Nz�����=�=VBe�.l�8�2���`��q�Q%qL9��p�XHe�Zz�^��31[ͦR��P+d��IhB�]o�b�C��_޻�H��(/T��+��/c|\�����EJ�<CI%��"ehk+�V���gDٰ��'qc�eݰ9�^y��$�#yՁ�����*��zc;.�.��h�S��D<�auS�	�̗�Úa?bt	�X�V�Hݤ�@&��xxVk��y�I2���j���5n�92"�k�kJ�2�r��[d��*���h�أ@����E�L�*`���M�$��>�2(���(��	��š�͐��w����G�g���X����ٱ��5��wE�ƕ�p��1<SZ�봚(�:�ݯ}	�����`���ƔK+k(�%n�Y�BS�b��|�E�9���;]�r�՚�p`BP����ط!l߱[�
�D�9�	BXv#6��˩�b�2�{�Xꮉ!#˕�4�SSӸv��6�_�v��Fh�ٸ�عk�?|.^VT°I)�ԇ���d���R����F K�P�\BF8��m�"*bS^Q�Ԑ�3�gT�#y�d�@Pa!�U﮼��?V"���%�TQ�`��	g0�e�������P���-�{LP��G�G��-\]\�29%�y�.>�?r����󯼍��:��������˂*�T�!������˕i��/�d��hq��a���<�1"�]0><��<�7n��w�k��H�VO�D������<��\e�УldC_��Ǩ����u*x]M�����I���u�Ne����lFo�}�ݾ���gA�J��Mm S� F�#X�-��\YQE��"�rot��ғ}P׽�5G��݃���OlA�x�οp�b�lXÝG{����U��wD��TW7�=�pf�;o����ԫ����2D��j�RZ��}]��s���j��"R�X�r{�ܜ��͘_��!�'��T-7V��#{��[[�J�Ԫ.��~���g��TŹ���k��x���-3C��ӟ���i���5j	*z��3xu���)�a0�#����bqD;)9t�׍��B�:�!ڷ��㞳�=��:�s�xþ�ZmMB��L�z��Gb��{�����e1M<���Z��0+Q]��?��H0�
Gr���b��
pb�6���1���q�&u���\����k�~830:��.#�ͱq�W�k�����ّ�|� �U�����035�?���K�����N��c�&H ntp�}1̫1�������Ĩ�7-ES���UL�����ؔֱ����̼/	Z93lN0��&%��#�,F+�b/sJ����yˋ�q��%���-�V�ܰzu�(q�t$do��8ge��)����4�~�X�e���AQ64V�e�NS���2*�4�$��O��ݛs�������jوf��&��^��H���S��"��׵��TA����cD4�8^I��Ab�ZS��<{�vM����&��P˫Q��u�3Fm�A0�d�oy�祦G��'��l:c	3�
$��,�c��r��܇�b}��S1�����8���{va��(&7l����ֻW0w�V0�Lo£=��mn�&^x�%|�;�	,̡#����p`�<}�� 
a�!�a�u/.�XN��Tf��mbY���������H;�ؐ�Z�bj�mh�}���,�#��w6�P8+_IZ�=7�0�������ٍ����+����z5���d����o�b��}#�i����	[�1�� �xa���7s*@̍M`���ȟ��"6V��v����:�g�M%>�u�؍GP����N0<6.������b�oj�k����$�F$�@6��.�'o�g~�A<�O���-���It��U��iA��7����y5�~R�"��5� �Xe�L�S���
T�)�Eb�$N*�ɵ�}�>?s�4N�{\C�ё1I�l�j�.�>���\ �?���Q�(�p����é�8
�`�V[et�5S),���p�	�AV�	����Nb��혙٬�/��NF`n�쓮�\��Hy�A�%Yأ�tT��ihV˅%���4�@���r�6xΞ�U_�D�g���63R�R�a]P���2��cڪa`k�Vg,�B�C����|p]ar�c�����텒�S�:��.p�-�Yn
;/c�&3p�<�������J�z���/�]���a����`tz�����e�ĳ����$vD�4�=I$Ri�2'��ޚS�­0�*"��ZV��3�if����9{��rr1Z-v�6�ڲ*ޤ^o�0P&cYi6{���"}b�l|�U�9�R�X���c�6lP�i��y G|���*ޗ�L����^�Z�~k'�,<n���g	���SO��ο�6g��*�&k���M�K�<��ܚ*U��>pc zZ���d�y$w�.͌U߈p.�A�*�,����)U�2:��Wn���8����d
hQ77W�����_��z��'ݏ'�~�=���"�2�JA�D��F���b�R��x!`�:��E�Z�y5 ��92|����zi�a�
�,��Ŷ�;���ʺ�u,ǕQ[]��p�zZ��!F���9v6�Q�9�h6���(�)�#��G4L
c�v%���Y��NI�N����u�(��5�<���:��Z���Ҽ�gQ�F�^C�VA"�H��*bX2T��&�þJzo5��QA�O��#g��t���%=�@u�ÜC��i�F�Fׄ�k�x��XV��u�<��"���Mby��̃���l�0�L��.��Z{�se����axbXU̮_;�k��CPŅ�5�?��������%��Y���U������o�g/����bۆ�o���r�Y-��b��fu�fD$�eL��=0l�ZYZ�˂j��:�<pP��bM�/��Ȉw�[���:�TPH˛�MV��鬔��O�ڵk�pf�֭���#��۷�t���J7m�c�?��^zQsKYG=� `��T�\�weuM�}Am�sTyY��33� *a��cT��H0��P���Tc���6�f̄n�t1��P:a�7υ�Sb
������Bڼ`���^Wfia8�+����y���5��R����P�'.̢��bU'�ޏ�[�+�(+F>#a�WW���ZOGL�������l:�V�S�emlA]P��*���lA���VW��P���}h7�^����)�p��{)7dx��ak�c�r�49ƞ�T:�/\eũ���A4�$�g��d,R�tLy~A�c�<�Mr�	�ؒ�jw���WV����� �J���妆9��a9[�_�M�lulz��o�K>��m����=����$��bu�0�&&'��4�塊��43rGT�I������2Z�����L�Me��������b��@�%�	kU�q��A%y<�O�W�����vm�����#�F-�M����%�u�6myR,x	O<���_��Pj��}x��~��U٬e䊡���E�)����#��lQ�V��<{��^<�����Q�w�.E �j]U�)y�y�ZS�ÄPIl�a~��؈v��<��4�:95�h��X��_��Ւe[��ƍ3Z4�����ÍUq'73����xi-�M�|@�%��Qկ|��)e+��f$��b}?D��2݌�G�N6��B���X�&��M�����C'�MM:}�*~�қ���x��W�����ѥ�)o2���fK�8sy�/ω��ء�ȉQ�%\��J/;��6�*�N�ތ�M�9:�j�zG�VW�ŎJRp>�����.	j)a׮�0.!A>K`W���D���d���*�ǧ�Qw�(x�r�m*፺�l���������n�q�(��"��!iOR��F�Jl��+	�8��Y)U��n>+N���ĸl�2f�_��S)���Ɨ�}����ʵ����W�O�:��}0"�����Jiu������*����}���|�����U���ߪa���qt2� *Ѩ,�8.ɸ��@	Oa>R��������'��/<�������X\Y���(6M�+����f�9�Zsu������q��v<|�>AEl����+s��Z(�8CC�z4x�ծ��Ҙ��C۫�fk��:�`��U���˸p�J-2�bl�&�dH`(Cn�3�rNE��A� �0i̪ʅ>�rU �l����������\����)9�(F�֭E��	$IG�7Q�+����[�44(b��u�!���c*�az��;6����3��<uZ9o��Q��(��$_����D#��Z�d���-��95��ui�x�(����/�M	I��m4��UF�d��NE����+�␊XX��Đ��Go(��"�5ٴ��.�xI7D�/l�w�-�����`ll̚%,��ڜ�B���kx�����'5������>�R�%���ݲ<�q�	a;qCŒ����ih3���PD�p�]�D{�b4˲6xmXy��+&Ɣ:��4w� �FL	�� y����s�.avl߲C��NT�r*Y@����fC���ME��������?�BD}m�f)+u=��[�3}��AK��U���mRFe�ձ��C�H���D0��DR��+���`�3�	L�,��͟���@D6�Fq}q��7��ɯ�� �l݆���c�Y&E���7����kǨ�#�������?�@��W�k�r#ȕ۪A�N�N�8��p{~U~&��xAMR�%��N,�C��Xj�ڌE��8/`M%
xj�r�l�f7�8u0����QO��С��c��&�l�|v�U���жqYH��&����Ф�X|K��ի�033�I��\�tY��;m��?iq�[fD�u
c�ϟ?��ڒl�%����Ҹ�-��Z��Y5���o������$#���]�V�U��6{Bc�s�"M֫%�]���B���_z�ZͳMC�@�p���8#��؍�&�[�uM3Eës�
�.4Y�01��^�W+���yE�CC�*�h�e��o��T�������oi���}��ݚ���Ϝ�51��r�۳UQ��;`���G�"u<2�������@+&�3Jl�(�e�����^
|}-�3�EÓa�Q[��@�%%�-ڽx]�J�ʵ�_�P<���'�S�s��^�zy\�]4+N�C�2�J-�d���>`0�i����܇/�j�W�g/���P��?��]�ӫ����1��| !b�&F$�����$I}C�n0c�8��'k����<ʤ��a	��Mx��-���������vlbrPŒx�<�S���|�ow�����_���*�_��?��/4����e���Zm�� �8���;wvǎ�B��h�y�zRպ<c\��Eݺyss���	��"!πlA(��a����*���_��~JA³�)��)��ܐ�,^^s�XbbYP�!�#1���v!�Ğ�fb(O�7�9Y���୬�h	����� *�sR+�Z��[DAm���̔ݻvbjzRϑ��ܰ�W�IZ�Fiu�+c�\��)]�������k���ձp�s`j�ln��h��ގ��^Z[E����PX���M���'5�^u��`�+�3��%�H�GmQ�ϰ�$�?�d'L`�$�˚av�G��ٳG��.�}SQǡCG�O=����j��~󆬏���9#��#��@�P�/��t#�2䔸�wE�������4�5���ҕ��h_c4p��6�sˈ�Y�v�:�J�eANM���#3ro�����q�6{��2����췴b��[��bsk��������K!�j�=�ɚj�WcE�N��q9���e��&6 A�8�����h*�������a��N����Y�i�g��c��Rkh��Z��:����#�87{��_|eg�X`���7���K�q��*J�W�1�H�M��K_z���bسgFg���ld�V�
��\�ko��"�YUO��Ȯ6R�`�l�?���ő�>7U�D3�ͺ��J|N�1&�ò�R	?dR�Rm�q�q���Z8y��>~ZC1~v��U�͎
T�AN�Il=#r͆G'�m����
��7�>&�6a��mz�u&C*%����_�Z>�Q�r�l��I���㓞<��Q�Y�2 H5)"um8�\C%�uذh��"��j\b/k��E�[�}�������Urhu�0�is�j���9+��<20Y�*f�^NGű!�'�:椾آtn`~f���'�;�p��bM|��d�,�i�]����D�9	�r�z.^��͹4�UEm�k���,/�0!�W�a$a�ο��{�\!���]cИTd��N�Ve��CR�<��=E�H�������r�&.�nb׆��8��W0+?'��jn��eC�quaU�xS��<q	�.��AyhB;Λu���|@�q��#�D�����åW���=I��EE��`�AZ��W�����������O2�(՘wF$��7�0�!L'�.@�"T%�F&���[�UG4u wNe�r�y�hwFi�-�g%�\��ډ�8sIbU����E��3b�:WèƄ�=�Q�B�K7.��K)Ԋ�����U�S�Vb�aTMk�"��
e�<r���Ł�;Ѣ8/+-��]���5!��3Шq�pS�hZ��j���a�'53���^������k�|�@�)�����;6�J;*�L���ݺ��M�S�=�J1�/�������ʄ� P��-�D�aR��?�n+�(ȄNSTu�Tb���za��_�K/��ڒ���蘉в]Z�w?S�,׹�xq y,9'E�w��!�d��(�W��=X��U�H��Z�^ͨ���3�H�Bm]�Ŭ�ōR�Pz����%�l���w�JzU��������TP�paE6��y�~pE��%���'@�d�fMG�,��jxZ�f�3_�pekD���m�.k�)��#'ꔊL:$�����~3�&eQ�n'��j��IA�[Ǧ�]���^����b�k��C:6#���V11�g��0W�Y8]1�em9��Tt�QA�m��F�R������� M�����n���Di8��BW��s�Mx�+��;{py]7LoБ��N���D�6��˝���*��O�/�$o&rZ�x_��%o`��#��Y}�n)��,9�:!���:���(�Rę��D�)KSK�z�GjY�wt0/4q��D�X����
�7
�2)�AB�#�dLQ�����+�7�F3��4�Sn7��+ީα��l͕A��E8xN���W�O�In���86�56�*eH(�d�qNk~�7ʂ����H��o���HZ��s�MH�l'�.�8�<�p^�&ٟ�a�t=e�^�|����୓�Ja&��؝�t�~�߈�z��\��8���-�Xu� �s��U�TRQyצ�1i�i��j%�ς���?L����(�)R��[Ҳ͆6Vd��ft"}S����[�U�pe�"º�|�acm����׼R��S��S���n_��Ӝ���!�O�HH6���fh���������O۟C-;w�:0�r˷�U'����ڊ�� ^��^Ǎuu��Ba�R�+�G�M#ąS�,�������N,�TQ�p����oA�IA�&��p0�F�g��?�Kl ��n�D]gQ�S�R�ՙ�5�9�*R��Tp_ڍ,�:�\��dP]	�'=�~`�$5L�F�A�ґ�#+�\o'���Ƭ��`i}��g%ih#�l�j���	��x��ydJ/���{Q$���]m� ��FN5U��0�G�'#!p�ذj�yqv�Mpg)�3��߸�˳)*�p�ا�����sY�n�t��5D?|	۷n�a�,%g�${u��Հ�+
%��nR��em��Y�l�m�r�9�������+S5	����Tf���e��70n6���Q���m �1���;�Zz�15.Uz�(��8#��x��ʴ��	�/�?����H�kŨU�4Y��a��|�_ġC{��X�2-Q!�U8�sy�4���UX��:EG������V|*�c�"4�#'R�5qe��ܰ9�}�P�U��@Y�Aî: ���2��ʯ��g��!�S�T!�;��:�VFƐɗ�G�\H]ǎ���k039�ݻ&�g�r�8��ِ�:��80 iF�]�4�x�����I��+>�M��c./�G�D�,/�Q�`�)���.�������q��܀��5Pe��F�[Q����	L|�h��Zֆ9��yac��rhwQ�uz.��M�"�Mȿ0���g~�=�����H�ެ�P���t.	�Y���ﶪ��d�M���3�lѧ@cbv^��h�X�U��-��}�[]{~�8��Z/���:��z���N�~W/�ꚁ`��P�%H�tzgDy�N�p[L[���B�L2 Y���Mc39�ph���\��T�9p$��5�"�&VfwA��Q����2^bS��*$���4|PQa��Ⱥ��0Y�5���QY�uG��� �>�p�m4"&�hȭ��,k��i�0����$&�WW�,YV�U�8���[���+oc~iU��D����ֶR+�w�.[��8�o7�=���6ʡs��0%�flp��ӂK0�S͏�9A���1I��v
�b�-�UY_��%HCۮ��O��.k�ύ��w�X�JUШČ�cߧ�M�������v�s��`O�N'��R�VkR��X�w�4��/��n�u_��"2�TW7����x`:�r���[l��9/�1�ݫ$��$�3|1�H��z6��Ʊ���r%��U4kk�jlR���B݂x�I��F���Aj}3�r�f�T�v�5t`�L�w^7uL���&j���E����H![�v��23�F�H�|M㹘6�m��3r��q�8�4��
ٲz�ƚ��T��`�	�z�����{���nQ�@�"� ��/tÚ�����H*��y4�d��/4ġ�،�J:��~���S��9���%����U,�t1=9%�>�Xŧ˳j5dK%E��J��n^�I�(iWW�Y���^��5r����z-)U���X��A��d�Ƃ:#�(�;R�F�Y��$�.�m[��ч����+h�H*�P�ӬdF9J��mx��3N��h-dd��#o���A�����rms� �ZI}~Ѐ}�I�w2�#K�\z��&���"�N�#��	EN���'z��՗���c��a%��7v��P�<sWE�SD�3��h��VJLd��X�ӱ>M8��A�P�av�|��}A�0S��гg�j�'V=�d�Xˍ�tvKV`j��gܘ�Z#��3����K��h�p����
�N��%8��i� t?,pw31�M#D��V�	��N�4n�9U�D�C�&���}����n���t K���&�E�@]�.I����^�P�GI1/ ?����T�X���ź:�M��{�|Ǥ`��Udy�$��k�Pq��Y�y=7�B��3�C�������38 ^t��JEPb9��w�g�!7�X-j�b��mxh�g�j�DQ�	p��4�@Ti���x��%�4͉D���ǚu#I��q�X�RT��B�߿�������XY��p����!�A(��t߭S� a԰V��/�q��u垐&���l�d�y��~�%l�h��w�6l�_��FW�����w[�~|&Q�G�]7 >诫�&�%�}BO��'q�Oe��.8E�?����E'��6�\G�[X�CG�隅u{!��X��9BT��Y�G���u�>r��f�,竒�ԩ���h�=q�Y)0C�B��P]W��L��:���5�p�=��M�(��
��1�V� �ݑ�J����GNPג�М�Ec�J�N
�"#�1/�ʑf���� �eHbR�����a����zN�ØAF�_��0Ս���~��W7���[M~�'�dޞ޵C��[�����3�����h%T�-�Ov\��U1=�����y�y���/j��\�att�겛z��M��zLH�ښ?�h��N��wY�i=!]�~(��Β���?�����Zm��R� �@�DE����9��?�����0�9
rg"�GlH��s�1ӱ#�:�KC(U*�~)��!q�ˋ�[j^��B�K@VWz�%���q�|����A�dƦ�s0����Wg��om�ʵ�B%-i���!�ǣ���Y,Z�0k����X��Ux�0��o�2��.�4q�Ӽ	7.��t2-eqQ'BաXfd��^�����N�B�(l��u�3b���z�r��Sw�=�e90Z��J�@����	���@���^V�ZzE2�lڵ�%K�<�BA_�8q@�&�ZJ��+H��]��ۼST�����6tH	������3�I����wUߚs��,��ͅ_i�Ī/��/~�f�����$ޡD��A���reMJk���Ls6���e�[Gˆ]+K�zZ�W��g1��|\��*l�;ZV��'��l�D�b����.G�jҳ���hkM6��\���`��0R�ރ�Ɗ�{�Y��V�n-��/���u%�IC!*��^��z}Y�|�G �AT>p�V�� D��|k�:Ù��Zb]��D����q�g� v���Q��7���>梇���{<�o{���Lqodd^�%H�H���i
�q$/"�rS;�i]&.wa�M{ad���Xl��9O��L�J�Il��K3k��Uߞ�T�3��5{q@�lz�dg"���"��MMW&#���0������k6��뤨��)���i��	Pg"�{WK�P�8rOd�f`����V,9��B���<���t�
���$��.AM��S>%r������8��4����N��,o ���� "�H,��Ԉx���Y�y�_�H�1q#1z*("�Ƚi�V���9	lvc�;�.�m�P�.�5�*�ҡcD�: ��X�jq�_.��~e(0�5׊9#m��]�
��PPwq�&�Z}m���@z5�^�B��yb%2ju��[bJ9�<�&�Q&M�3$f�f��!�z\�*��-\ޡw-��������S�X:g&\ߗ;0���ׇ?"7W*�=�u�����V�^w��0�T��)v,3�(p7`㧩ٛ�2��7U(����l'mg�E��̧A��Ŗײ��z��fم8����7A�$��׶�	�1'�Ü�r���
�,�6��6�����!���(La���43��Vl������i�~A�=K����u�FD�ն�M"w�{n�� Zxh��ڇ=�������:�9�r��:�8�4m�r�p���
�ݽ�H��4p��a���J|��� ���9w'i�]�i2:����q}�SWA�<���8p�>�m$���E�x�.^��3�$ U�EX�Ė�ѹ���!rWXJ�Aa�u�x�\��N.t�������>%������������VI#W�'�	��ح�k�U��ƨ�
���K�j������Y$��XUɧ��*�����)�p��;���Sz�k���<�ȴ��h�y�}/��)̉�/IU�WU�JN��jkytc+*t�!��jm�k'B�,�dT	ͅEL�Ɉ�b0��)��,��bz$¦�3S����2�^����blk0�-��)-�C�������qƿM��A ?c�kת:�T��Ht��`����A��ǵ�$_����z��]W�]�t�!]�����MRh鬒n=u�P��.J�-a9�z���JY�ػa]����}����;�JQ��3��;��bq��Y��$PH�6'�zkx��Cؽg��6~�ӗ�s�LC�Ń������q��}x�Gm,�캦&<�8w�^;vo��>N���"J��#����P�D/]��ˬ��=[W���f~���Lzh��u�݅ۡ�¾)�3B�-z�Bq*�"��%i\�/F�\�Z��c���98Q� ���8P�����v�?��m,�]3l�����u���cR#���8@�!gM�Ė�3A#(�4�Pq�y�Kg=�4�b�5�q�7n��]qMI����e�-v]h�kЏ�����x/��Q!�ZF!����aۆa|�3O�Ǐb��~��/�^����J��Z�.�!�Ly�x�Zh����܉/|�(�{gΟ��[�	a�B5"�[0��հi胡ϓ�|L��H�<	s&�8��ԃ*�	̛Ʈ�J?�%CU��t#����3�0�j�9���v�2_��Y"�%V��{�|8H�s�4"A�A��>�I
k=�U��M����'⁃{����p��a���I���۸�$�M��#�������u��/.�#ze~U���9=���x�𳟽�?��o�(� $ѯ���>>f2HxT���5
c���d@��6OƅwԘBFL������ӛ-���R�j-Vy�1�Aj7�)�fK�oV�b��5D�V���rg�}���vV���Nr���$�C����2��-,�2~���?�?|nſ��ۺ����5A�H٨���A�ЗH<D2N�TW��� �e��%��Q���gzr�k�+I��,n��Fd2^丁fsY�V�ٟ��كᡌ��r��-Gpt�n��/���sx��W��oc�~��ve��"Q�~�0~�W>�H����U�5�`�Z�C���_[[�Z��a끻)��.qE��]���
:՞6!��>����4#�S�]�!��&fP�_a���G{j�b�㐐ħ4㖖s��έu�}`�H��0Ėȵ�[=��H���Ƴ��R�`�7�e4��ݛ�ç��O~O=z@����j��[p��6��o~	O?��������?~In��WtЯ~�)|����3��/7���_��?ʦ�_p!����U�ǷIB���lX�#����^�ay�g~���u���%S�h�7I|��쩡&2�"S6Kܮ�����*Nր{������n}#��H��05����8BW���pN�!�;��:��1�С�~Z�X����" ϑ|.��IsM�C
@��r��)�#^{�ΜEIN���6�3tcC �=2A
{/v�Fn!���,�A�H-h�������A�Hv������Op��.��-?yQb�5�,H�;16���w⁇�`���(��$����	�JX3=1���!}
�Zkmb!�$vr����Jq��>�tZ�����ZZ$^4_,#��<N�KT�=]`j3\",���o 1
{<�Ĩ���4 I��kr�E�߽]fN˄ډ,�re�&�@��Zʡ	�e�Ke�xvs�W�&����I���%�4{��$0``�W���L���'Ã��E�y���̿��k>�_��/�yDc����o�/��o��А�So����g7.�ş��ױk۴67�I���C��BgDLr��*�[.�*8����i��%��H�q)��GiH8�����I��<XIR�X�[Z(�ЫВ�Q�����/�l��}�S��d�	��͢�����u��A�Pס��Yb��?5?Y�e��d����$�c���x���5���@�"��	�Aѫ�E�Y%��ژ3Ȳ�����J�r�7e��ʎ|`�]�Bdfz������qK��ە�Xk,a�q�ɟ~�l�������+X�����頜��s_�>�K�a��)}��?�^x�m���Y\�]E���rmGn��Zs��L�V]�"_�͙�j��U��l���(f��ੑ4x�*��Zu�{P,�*Z�52�&�)�Ƞ&�p�":���+6��0�+�P�� Duq���w��%|��UI�
��5��54�Mܞ_�~�^z�}\����E=��6�5r����X	=��~������~@�/�C�DQ� �|��v�ީ�}#b��BO�L�Hø���4a�!f�jG�b���}!du���1��w�o�5��#� cRp�P��&|���/���, SW0��y�箹�Ę��\�<�8�Du�S�	Uk6-�B!*��Ċ4�aV%@��$����=�#�n����ǃ��}6&�H�Cg��4�:�4��}�G���vۋ�م&���zZy�f���=053�+�D�Ы������<8K��'���`xD��~��@��^��g����ZR�ڙ�*8L�Ңnߺ�>���V������t��E��%���G����ƹ˳���>��Byh;�m?�;_���1�n�Kx����V�-�Q����!�jmN���ǵ�.��:~�2��$.�û�m�$ŐR�s9Bc��\��V����6�|��D7o,��714����o����P*f1T����o�7~�K����N^���uז������3�y/2���c�1/�}tlT��O��i��2�<k�\�x�2����4O@�����psP��!��µ�ؿo���[v��Ï>��_{m4�_��+151��[�p����|��b`J�b\���{{w�QO���v/T]�L�I���R���'鑃&,=1�!?H_?����|����xf����q���i���h�����dޯ�
+�o�;�#w8�د�;��;���_Q������k�^1���6��
01=�9:�ܙ��g�3&�GR��G���d� �o݉|��{��<�+� ���fy�����Z�sK�49$�M�7L`��&V?�΂���֎�̏���+����p辍��S��4�7���{�`��	����	�@AQ��(�fW,L�FC4N�wsV��д�qCY���E����C|t��i�MH��eu�p�S��/؟��Ó��8�sضu�K�%l���_�>�/ȩU���K��� �޿�ReG?�/?�vN��e���W�������%C������>	��EW-���������5�ļ���r���Z*�j�?~	;v�@F�yid������MS�[ZƮ��U��M��ѽ�N��^yo�wA���&ɿ���������Tq��*�8݊�)p������
�\��/M��?^�F� @����}������|�-�/&�g�|��e� &�|Ի�����d:��A��Ͷy#�#�޽��2�6V��N���O�Cb7�אHh������I�벸T��J�ŕ�L�D�q�C@�?w�*�J�4X[���/������6M�K���Nx��),՗�+����$*�!�����q���%����Ó���}������?a�°�J]�MT��e�P����7�����x1���g^�)K�̪gCk���$t�e߈�ڱV/R�	�<��AEZ�m[�bTP^T�0BV�ꂄ8�8�c�+C8}�<��o���fn�7q��˸��y�������{���}x��H*%-Ww����L7E�L<�t�.݌I��$����)��<r�������7�zٯ�6Oc����o�x�J>'��ƾ#�a��?�4��\��H���Ф^��/g���?Ï_{��h�7}�����������A�K~�E8ة����G }/�h�2�!������.~J��<������|�o��k���!Iݦ��/%��"/��̈�fm�Cw���p&��-��˕���n}�F�3�}t���D{I��a�X���]�a�M�PD���?z���o}�ػg��w���[���
�/�Ti+ʙF)ƕ����x딄>�ů}�I��:�BTԊj��.0��J��w��ǆ9�N���$��^
#1!��}BG���n�"�BIv��7(���eTGrȫR��So!lw�g�f����p`��'�z����3����5���7�9�Bc��a��!l�4�a`��T53��~Ǫ_�E�F�$���K�]��E�O�O)C��iV1�����<+��ٲC�H��T��)�8#��<���lGX�FS��J��K�ސ�|��)?}�M���S�N�Kh�5���x����#�͡��o=o��2�ۼcL�X�A��OfE�V쌝i�xD�f>f��g��_Vɺs��['�x���u���M�ϲk�^7��*�eY�G��٫u+����	�<�!5��	�O����)u��ls:}�X�CNr���	a�h��x���%�~#�,x��a��7q��Y�k#�Z?���d3V��o~�ܒ����U�ɋZ5�rsI�$�X���a��܎�<wX���ڭ���KJ<�o��J�n�"�ހ^i ���2�j_�vOG7r�D$�ٿ�������k9�>	H�.d#lߴu���K��t�_%����YT�o�{���"׊��G����cQ���d`K�u�P���rmYU��,[�s#A^L���DǀR��'Ͽ��Bf�=,�/���ـ�;w
RڣZ�d�֚\�uWU�w�4�d]�:-,�ֵ��82�U�,�_����*D�3J܀����
S��&QS��f#��
O*�4��c7��秆½W�]���g|̖Tt���?�q���!d�Z����_�T�F�LsLڡ��gF��T�Xu?�����o�q6z�����?�L[��bt$����/3�D9���������?� �&��q����Y3�k�l�@�M����t�1��G(�WN���%<��aTWV�ܫoˢ��j}A	խ
��ahD�Q)���Ю���^ S�2�"&�J4�o.v�)TbS�$�=�d�O�i��_�����cfBi�zBW5E�z�s�ǋ�Û�/�vF���R����6㫟y�������ZC�l�(�I��*&	\)���ߑ��*�g�|ȪeY�)�)���ݺp�Bm�F\]�J��ױ���y�k7����x��W$$!N���fU��r���n��S��G%1�JHG��wZIڡ�=��1����o}d0�"L�;(��P��1"�\D�a�'/S��z�dݷ{>|b��	g�o�!���Ϸ�O�<<�#PO�=b�!���/�с�Ndt�T��!ˉ�p�Wy��O�1$�Z�v�:+�c��?֞
o�U�R>	��[�Zm�EK>O6���F�.w����}�ئ�N��$,k%��w�fsU���a"�ݔ��3WpJ���TFT�����l����
�,�ժzuc%��7�<�*L�%��C�sŒ����F"�7�A9����)�Vv��+���K��3?ŗ>�il����|^I'̷0�m+���hvJ�{ꁃ�������b7C�q�,^{�KDf�
� �q�u�I��5rn�A���T���l�&蔩�k��*f�suq��+�WQ�w�����q�(�5�ߨj�ًrh��%�(W����ڶ̝P���S�n$_b���J2�'q�V�Hs:�o~k��<���Q�#}X�cK�/��|�T��J�����t.n&����G�`4��FQ�kT'{G'�?.�]�α~[;2h�J�>?��=Θ�����HuU���<�R˿��_*e4BVI�� ��H�>t��r�\
��F=M@�A:/�&�Z�ɺ�+��������M
�M��K���q���
�s�
�B���q�,�ouk:͝<��R�I�L�EF�R6k���2:�Z���RҮeI%
?�y$nΊ�)�ܔ��<%87h�kx�yW��P��Y	�����ǤqN°� ��_Wgo
��Nf>��]9�pqa	o�u\�E�r�,�P�ÙǛ��w��!���@���g�Ssq������F����- �F�{��R�}R�H�u�jyc�v�W3R*��|]B��$�������+�8u�V��*U�*���/s4V�A9�B��C�+�"�mފZ-�����R���/~�^T���\iz1A���	\C6^`:=(gh��.���ҫ��uc��F"�BEw6��4����	^x��a�G��=,two�w�~]^�p�Z����n�V�N����ܑo��I%�v�;z�#�t����0�g�egk��q	Hz"6�qD{I(G��1��s���a̱*he¼�n���eb@��I�lP�OP�UP��øn��9R�U��,2p��+v���uS*�֦*�>��d�;�AT��B���B���{����R�"���3g�Y�p���c7��A~N�ҍ�.r��N�����_��<�9�w������K�HM�>�s�ǁJ�Q�)���� j�c�^���'}�!�1Y{Y��c��$YU�g��D�v[���n��g�z@�6l����hKt�3�ɏ�Ǳc��jd9m��)�i��m3���#�¾�{��s����պ.���jL�Wy��������Y'�B<W�{v߾�Hz7�S)��,�{��E�"=/$�a}a�����]�Y��q��"���.�`�<ٳ�x���s�6髽���c J�E�\f����U{�a(4~��:�u���z$b����R1�й"�.�l��^��͕,��9������H������Zd8���@m&a��CؾegN���޻�FoQHY<��"�I/Rɜ��]g�(?�+�9Q<g���\MLƉ������V�2�A��N:^2JX�m��J�5-'t�InuEY*��1���R��1��	���o\Y��o^G(�uuy��Ż7W�mZ��igDdv8�G�1�k'덈[LVMY�!Cʮ�!P&�l��ݪ-�ۻ���'��#�pr�c���� �'���}{vc�����}�G�5��atL��1���/`�έ���B����^}�m1��;ronm%�]�s=��ˀ�H�j���(������;@����n�I�{�`�88���)w�ܯa�*{6����a�����M�Dp�����M,_��ԁSL�}e�y�FD��]<Ǜ'�ՙ(*�jc|�>qɣ����)��� ����M���e��:��b<��!�޹=� �'���� �Ͼ��)q^����d�Ӗ0ef��O=�0���c��x?^x�]�-�����ţKX����vm���X�\�X�/��]e�I�����5<%�<v2��EE��T<0���57�І�sq�kv��[�ŧ����Y�:�ҙ\�F3Qi-&'���o/�@ӨĦ��0�k�	�Q13"\�*��br����f6�kL����.ߠ�30�Ȑ򇹲ܢ����|�G
��_�>�G°^x�u�~�4V%|ܿk�?�W�F��|���1�����޽��!�I�8}�<�C|�'ϣ+(�\��ε���OF���G���nC��C�>���w�;z���;�R���oCRq!c�{�گ����k|�ǹn|��>����d�F<�8�M~w�kw/H2S�'N�k���m�]�F�m��%�G"���@���o��J��?�6^����0��,p���S�������oXo���8w��Z	��l��%��c:�s=,5�p��%ٷ���}�wၓ'e��5�]]�O���X�6��,ѫBA.q\B����Hb�!��*����9��<q�wƹZ�ܒ�M��*��݊��6��������;����/��co�F�����ڲ���߉���ȑ�t���}������'1��8'�U5	��A���-�o��x�
qA#�&�R�!62y\��O>�'?��ܻ�^�������� ;�o�<��&��/O�a.��'��ż�[�L�q��
N����N�ŏ^z	�/_�
/��qh�n�L�êh�c	��F�oC|nb��_��� u�z=2��*���Zj��r�D9x�|�.����؅H�/s*H0d���{_������A|�A�HÇ3� �������b:�أzV1c2sp���FG�F�%)T��55.<��$�����ﻦUeu�j�X�����^u��"��;?Ŀ��U�����<��:J�K��A�SC7�Q*��ZųϽ�JFB��?���m�������ʍy,S����U�7C;�T���p��r�s��|�.�H^��8���nv�̥�4S=p��Q$# �3D����S����;6�@��XyA����_į���������+\�p�f��G��J�SM�jx��c��,cdb��8�;��HY�w|��Uo�������eȕQ4�FƠ�ҡ��l��ӣ(�!�0�gr�_���X�s�x�^{�]ؿ{�Nh�ǎ��v��5��?}O��X�6P'�b~)WD�*�:��ȾQL�f|
Rgt�N�"��:�'zG� I��|N��cp?i���#w'!��M�״5�Z���/v��}}��w�'�mw�G�`����p���y���v�]�qǱΈXiֺ�"�It��8R֌�۱�_��ѫ!��"��r����*��N��QKƉ�����<���6�wy~�$�����m٬-4���ʛ�Ʒ������zy�=u��[�0�>-��(H�o���*��'�U�Ud��\CQP�c]�$���	���|�C�<��sC����.�6��_����j1���wQ�{܇�N�)���F0��F��W����m��_l���M�Jy�Mu���_�6m�;����БèO���6�O��1��ӗŀL;m���?9�"�=�X�ꇯ���Ӯ�$"܉8��Rܩ%�X��h�-$��k9YC{���PVg�$�vK�D%�FUd⦢���9qo�u
/���kr�,���P�z�|b�tq�2�6�\����8#f�u4j�K�w��/�L��� /E��*&��J�Oy"k��!^����&�t��_q�^U&��$8��
X��{=��܅|���C^��A��=����jc�+GNH�c�q�b?��F�vQ�����^4�5��)~���u5`��[�2l�҉i�I�����
�#צ�2t8��=��%�K+:ؾm+v��.Ooif���.�xtt��QA'���i3Ih�N�6��L�	p��q�9��z�~�_�X��bWl���@�=-��FK˼Y��J�B8:M� ��c(/�ӏX|G��~]B-ph�:�.8'zæظi#��l�y��x��^y{$T��o~{�n�0���G�S�+�k���B7o��ۂʾ��sX��Ua�]�p��k*d���QȢr��6x����@��j9�JV�7�5��j�&�,��$�1Z�0��*�5���g*��c���9����~�ݟ�B������K��6:�l�p��\�&��Ǆ�=Lw8��D�n�x��`��q���2�?<fq;;p�ꖴ0G�6�F
�f�`E�1i��H\�3p�m��~�!��C�4����`i����m�{��Ġ���K����FLY��*c�>,�?�X�@lݾ���Zi�W�)y�+�ZF:�ǘFCvI&�ڦq��.�6�*
s��i�Vu�q.P<���P3���?�",isL���ۦ�m�%��nhq�_N6]A�ga�Su���r��O`�Aj�+�;��C�4�j,�y\�_L�w��%���T��-�M=�7O�Ə�Wo�ƹksJ��_����#c�-w�)���s���Y,���̹��r��j�JC�̌�:���$�6��q�[�n��-��4���M�m		sqQ�P��+��I�r#�2=&aX���m��4����S�|}ݰ�S%<x�LSͼ���������;�"�w	K�+Xk4T��!�cvv^�h �W���5��7c�(��8wn�G}n8�?�>-<14�M�h.�a����b�e�/�m<�<��[5=x	I�Bǋ��<�n$>i�Z����G���}�/�����a��W����DJ� "i���v�x�{�氦4�|�F$�P�V��|y0��V=ַS;�1�|���!��4���Fn�w������x���x��tA=���"\�6��s�����H�*�bv��/��@-T$ԙ�(�ОC�ee�Nk�����Z����q̯�s�[.�Ai���yϩ_J-]����͔ĝ��A���t`�k�x�BY�̰�P�u%�����߭��r.��R]Au�2K7Qڌ|����<������ު��j/������eS�����ddx�{&}�G�����d9��fn7U���)mXZ+FQ�������]��166��~���MrY���J��^7��ᇟ�yH[��ǧ����՚8� ��s���w���=�._��T��vsx�8 j�˫��
<b�!U@sk/9{�!�>��[�n�+]��>fD<���U�R���܃���)HQG?���Ŀ�^�O?��y�.�4�A��ű,�yz��K`�/1��ڝ\���K_�	���!��F�v�2G��?s���_~,�#���������ݘ�_�sϿ�c���ZMB�|��#��d�NMm����p��]زig�u��:s	'޿�F7DAC�R�!�v��`kN��)	�궶 i�(֜�����<��Q���D�c�"s��#eq2f���`��
��UL�����M�� �iiLW[(�{��3����ҼM����yb �_6ȦgbZ)���>�a9���X���R+#[j�37��2竒�R�{XZZ����Aӛ����46VD�8��m�n�X��X���E��"FF�΢26�����x�3O]H{�������u�.g�ǻHà0uj:�ş��L?�����.��y�t�����Ws�OM��J$N�A�85��!�ĭ�t��cC'����s|�!8��?T����%4�֏ф˅8�K;�^��u%%�Xky��d�~������ ��y�]��aՃ��C�_>v
��6�����'P�v041�-;g��a����<��I"p�����"�VVqmag�}�o���x���-۱$1}�84 P�.�տi[��tC͹�I��צa[��u�Z.��%�
`��TDQ�Hi�q�7o/��܁'�imdk	L�03%Fe���5L�m����8<�[�e�/-+zٰy+>�r��̏pk��U-���t4�����0}���J��/MZr���zL8:;$�#���Dk\�����7��,��� ��}ZQ}�z��s:_fyyAG��KE����jQP�y����SJ��^īo�C����g?�X[��C
/]hf���x䑢� ͵�a�~xá!�P;�>Yj�tUvM���7����ׁ��e�r/�#�~F@j>z��Zs=Ww6~�#���?�qў�N�lw]Ձ}���3��?aB�g���YZ���&Z��C=���N�S�h �1e��*�A��9{|bZWW��O��!��+����1>RV(Db.�0�����"���)����p]6�[�O��W���7Na�Mc�,���P)�ڨ���_���k��Ն<%�9�F*?�;����}-���~�--!���hw0R.���<N����y ÕQ<��_��E�յ���5d�����9x�(��VV[ZJ��PF��i<����Z����I�ȀI�E��T���:�16
��Eр2�ܒ�ŊVԑ��3b0�X^�d�S�������Lљ���^�p�Y����0�h�L��b�\�C:���%� �V�}@G�ˣ�H)��HY��i⾏v}%�Ϣ^�O�=X�����jd����ǣیI�7rF�C��*|?S�~9H=_J����$�u�$�������4P?/J�f�fK��_N:/�	xs�N���X��d�y��&�W��5[��őw��0m�i�ۄ� c=!�bbg��r��;7���������7k��<�=��o�gUf��F�$J 1QM�ZR�l46�6�2�g�mlLm�6��ZHQl�$H�(�P��+��w_#b��"�MUT��Ғ��̼7"��s?�~�xB"V�Z�3��?�J�^�[�M���{�ŻoJ�Rc�e}����ں�//gN=,�͎\�~C��yܕ+׮k̭!OPWV�Ӽ�렗#��',�!^�������#43s���m|$�;(��4��;��Hhba�3�7�H�em�,c��8\�����֭9��)AbC�b���⽭{,�! �۾R���j5������=9��LԃO8&����Q(y=�0��$�!)�a��N��t��ĵt#83���}P,%��$��~�2��Or���.̒š��"ڥ��>��7����1�����r0�U 3�����t��Ρ�5��v4*"��r��<���ka0����8��B�m�#:S!]�aM�,R�l�4��PQ+^�6G���a7Ьɽ�2Z8�<6�Dh	l�Z��s�i�M�ݼ��|	{h�a�Ԧ�Mm�'�s�{���?��O;�O�{���>K��6Ɉm������\6�dϐC��v�,���6M1v2�#Q� T,��4��Щ����6��P��1�`c�L.p�]36^ڽ�W��(�r���dT�`��M���_E7PY7AA����	0<[ݖ\������j�klI�s�+��\����6��d�&��hx^Q�혲6�Y-|X��(�0"g��k)���\w�C�k��
�?I)E�K�ř��X�T�|�TY���'/� 6������z��D���y����8,2���E�	�X�Q�*l6��RIk��Әer4%���Wv������艍]����
H�"��f����gSԐ��FAer��L�d2�p���$F�4�Jn�ZSTHH��!���o>чy|
^�Q�> ]�����O�Q9M�krH�%,Q5���Af����[RUTEc���:ᬢ�c.0 �g%^$�s��(h|���d��ԛE�>�_S��ѡsB��T���D���NOJj��  �t��o�@�yV�W�?��b��z3��<�uʅF�t亴N�Z�R
 U(H���͝J�i����%g��3�]{��}@/��7M9��ΘI?8��Lw���^���J^5a��PUY�}����+K����eI�0"
�Ơ��z�UY֯�S��LL64I}STv�C� ���D�L^H�A/ojn��]X�f�d	.�S��4f��Vv4r3B5���f� و.�H�^�T�PV����DO"J�$큗�*?@�C݈c�F�#*U6f3M�}�=m��D�S�/<J��I�RM�m~{����'ϛ���' ��bw��>�2�=�y�y�mو7ZR�0�/��>����F;8*< �M#TjM�P���̡ɞ�v�7��px�x�	���ˬ���ų䤗�j�	u�>�D�����c9�n�YY��ԛ�����rs�����]���,��d+�1��-�w
>d$�г���� _�=:�P8�k��@̑%��~J��߳��M��ZK�_bD�͛��N?y^�)�A�K�V�!I�3�5d�C>�Xe�S�kH�Tͼq,E��W�q̃	��!I�VifF#v9���H���k��Br G
��Hᓢ��T����|Z\Z��C��|('�y�$C�;��y�÷#���aW >�~��Oe$����bB�4T9C�q8���&�<��)��sC�Y��f1�#�u��DmE#�'����@��K����cn`xl�+obR���A^���\ ��f�tJ���S�1gCr\LG�s�!۞$��Z3�,q��O���^w8iKI�v�F||ؖ�"%�g�Q�gYQdQ�{��6�ӈ��=�|�M��PG�PH�@���ci0YhL���+FSV��B�³DI�����2P��bM\)�{�h�G�]4<�K�q���>Y�z���@fbl�8 <o�{����,�wM6����^ٺy�~d9��ȱ�p4>�3��yͥ5�E��D2�$�ڐ�ڧ��I�2?Y�ן{oR�K߳Y����x�r����/��>�ܑ��sj>�Z�$>j4fr��;�͎����V�S=|yiU�EE��I��,DV�Mά������D�#z� (I:�7�@S�8/��; ���1�t�?�P��7K��C��f������xc&>c�a+,`�;(Ёn���u�u��-ªG-#�S0���2���&�����s2�YyB������%PM�ړ� �{{m�+2�%6���<��Ru/���n#�d�Y2�v�Ċ�ZY�Dj��'e����$�\�DQU��ZEa��P��)P�V���Ʊ5�*�zoo)�2�����/Ԣ����|r�	i�N���۴��t�;��1�Ab���t��l�-���,iX3��{�[��R��*�q����8X�2u�|<a��R�`
�9��ꩁ�z�	�ӽ����{�◱�!�>�]�B����#���Q<�8=ځ-��5{nُ&���ւ9�%�uMzX�nW�`"�0MJu#tg�s%^{gK�$V��pV�5���Ϩ���֘�<�X���*���Vvh��.��^|V^�ڳ���(���$����5�gڤ�	ci�P7!�v�h�H�2х�S���<�ɬO�5���֛7��_�#���cY.��LVΖq(#I�j@j�]�&�x�f&��
�e(�\8&����z눚��i�/H(���| ��`nM�+0�b�!x漆��ؐa���Ag����JM=�7�ȏ^�(�]���	��y�T��y�8Gm�f����i���6�^��h���g�/��K���g���Ш)jS��H�8�h��t:�T���qj ��agNea�&����P��1�Rf�e���z������S�a��tZ�:�p��y���$�+�<��^�4J�W�=y�s���0�������Ǒ��H�g�Q�����,�aح�[Ĵ�B�tp�E�A��G���N�7Wn�_���˭����"�p��p��獃;Qޜ���@fOi
if�:�+w�./���	٬�
)u �ބ��1�F� ��Q����Q#┱s���\N�$x��3D��0���������S��Yt��\�PVwǷ^�=�?��� ]��=�÷�{
i�C�ġ�B!�G2&f�]�j]��^�i{	Cf������Fߣ����GQ� ��۔�fO���0�/ob�I��f��8�!V�0�;�/B��O�������F�@�VU3nȝ�6��0d1��d�C��r!9<��<$��	�e�X&����\�GΟ������]��C���k��H�eT�O�����K4��ܕR9O$�����O<&�e}�TVz�"+�3W���^��cUG�ԆN`dY��Z�W#�~|Y���A+�^|���E��a<t�ܺsO޹����|����0�ZӪ���Isػ̎��d<�O>$�G(kE��R*������3����Y�J���)��ո��O	���E�����#$R�(�Ʉ�Ld��W�,���\��suNEI4�I��������C���9{��f���Y~��"t���V�O7���8�o�q���Hՠ^�;s��H/ϵ.F�Z��{��H�Q�C2��(vڳ\ 7_�R�Qd%��ׄM]�e�!��+|"/~�k���_��ꚴ��)*9#W>���)䌙�z6�VT�[�M�1��*9����N�C,/W��s^�Bl1�ᱡk�P��[�&���=}^޸��4��P�1������F��~�(½Q�4����MH)�'!���q
Ǐ�[7�nR݊R_���
^H< ���`�����Ƚ�����;���eST�=H]Þ�;�XdM����U�c��Xu�'�q2~�#¥In'��;nD�]��^	�`��k(J��;�s	�'��{S�5�"�Bi$-�ױTt#Vd�t�`����ݼ6�Xd���j�J�l�v�®HI��y��3�')���wɍld��]�y(_7w�(�>������|�=���R�p������^��2^Q�b ��.�ڂ�$��a��L�j���H�x.�^��G<T�g$�,�2��h�KUω�)B|<�@��o$W�6 -����س�yCgİ��3�#!L��6z�����ݿޘ����g|�*+	�Ü�X)���*+����v���qu,�Xa���
ʞ�ͶĞ��4	�0�e
ک1J{�yW�����<gh���n�p�^�1��j�5&>����)�}ˁG==������sU�{��eqeQ7���A�)����}������m�?8���rC��#�9�ɨ�#U������Ԡ�{���$L�8� �B��8����P�Ǝ�Eutw��tJ\��kU�w?�&�r�R�	%�=��Z]"),Jo:R���b�qq=���6'���̐��bΞܐ�>zF��g$���@f0.ꁷ�R�g�}��J��#y���f�'8��d��-���\Ұi�p*�6z��W�Ұd�7�8r�	�i�ZV/����������=�&��zϏ+2�_���z.�#J��eIK}C��D/su��&Ns���3�d ;5�^�L���"�>�F�����/�?�rI��2�v��NZ�����ڦ�h�2/��	yE1C��Aj�ry5:��|����?K��Q$@t�_�Xޖ\l�Ɏr`oa��Yb��Yi�h<��d�q������V����}�#4�-$��dr�LP<v�/sFq�s���
���`�Ex��X�A
>7�Е�=g0�x�+�)g9�䑌#r��=���M9��$y�x5G�|��U��m��ۻ��C캶�B���jӈ,�gG�~����BjGc��`��Cʌ���7�����Ԁ�-ߠ� b� ���d)K�[�|��H\"'�v]f�}�<t	+If00-.T�5ؑ���������y�(��w$u�z-=xc�|��M��A��0��v�\(gO�����e�K�XN��B)�T2�>��f-x��8i9o���_�NGf �u��Y���l������W߽��"ǼՂB�B��F�/c���_`���o���k�zW�[[��ڑ����T�n�ȳ���ӏ������S�/*z���➹�ћ�l��1��;�)<��ø��;�ޓ�޸(��L��ql�C�Ŏ�G�\��U@���UC�gHaJ2uCE��?y��Ϛ�F%��#x7�"IGWx�Y��e�5s�ȷD���<�]�����f�g=��l�ø�ԡ����S�.}� �Z��f�+Ȉe�F�`���O�Aj�e�&W���xn���X�����l�;{�ۊ>;RW���_�\���|_��P���z����. ��1ܨ�'L����
d`J��0��H�ו_|J���I���*Qy^DbPZ�|���f$��O������f��2���P�����B=��LF4�k��uC�"�������/������r]QƂe{�P:j�J5T�F
�rRTșS$�S 'ݨ"3�������5ɴ=�^���d@��8��a�-w�n�����u$���s�K���K�YI��s��c0����燉�ʱ���ȶ"�D � �f��<�<pU�����S+)f/�b�ºA�{���J���.5y册Ʌ1t��/���r)�4%\!��Gz����w�h�5����X(�k�9͓���?u�	?�VB����`CVNM1ȼrڼp�o�R�ֿ�e�W3�绞7a��3eb��3^��y�f�Ze�L��eU>\3���hI����>n��h�*z3�3�n�۩���z��B/�\ְ�ڠ���D����.��+W����/HX��[����$T�L�an�r�K`��x@+�$���wvn�A�@�ZSS��8"r���N��gl&�<2��e�E���#��v� )2K�+�{�^_Y�����@ٶM�e{�k�&��x$�;�1D�9*!c�k�u�����U�u~l%�d��g��T�!ef ۈ$��+��p����0�iC��X�J0�|�L�0�mꟸl?ΆiT$�A�)ϒjı��iB�	�\���0�`b���bV��߂�� G�Kܐjܿ��&򭟋�RaX
�H��Phcja^f��D2ف䨦0�����B�U��|��`��U���IG@N-�/�+$���2�U|�����ؒ���i��t{l�T⒬�ZSq�(��X����$��5�h��\m��~b��<�$En)k�J+{e��s� �����
��$��{�%��]/���&r��Y9s�<7\I-8,^�y�ML��L(�S��3����, �@�P%/�HL���'�3�JY-j�Ÿ֔�ͅ���w��D�����sF0#ٹM�ɑ��U���[8�C���r B�H*��{n c
�QQ*ʃd"J�#Yh4���M8k��ׇ������&ti@8J��3����0�wg��g�>��2�0�K%i�6$_ɳ2h�L;�4	��m8 (���O�|f!;�c5@9�c�76#&��I����G��p&�>�)�hF#i�z/Ne\\Y:Ns6q�OӘ�skBb�\���yДv��?�H�m=FHS'�(�f1�>��7��`�h��"��@���Q���Y��'򚒟R�����p��4>���Ȁ������Z��^�N��K����4�X��|���׋H+6�S��3c"��s��r��N�<8�1�d�	�$fH�;���NO�1.��V�Ŏ2;�)�)�v��-�'���:lI�}�U�\�OX���-�-�-�>Ws<İ+E���x5��2��g�Q���:-E%B[�ЏQ��!�&PϑӅ�x�M�9 a��60z��m�S���=�5/�8:��>�\>g1O��j��n���_Scْ��]54	=4�`7%#u�j�P.�;���`8��n$;��k� $�JyYZY��}��D,��)��������0����PA���>�.�wy5��1��zeϊ�'$�e�A�F�"��F������'ZA��%m��|���xD�F_T���<��� E"&�0����ϡH�)�A�v�_cT�t�MG��J)i�S��(0�h�3⡗%��\�b���(��K0��0�����}F�z�\��I�ZJ`
C��Ϩ$���B�#�5�e���p3˞�}�HfT��_iÞE"���ͺ�I���;�S}.a��w��w&Ie�$�36 (n�o�[LD��N1�!����F��ĺ�|���ͥ�	ǘ����7dm�(���L��ͽr. ��*2�8���Q���s����1��Dks%�C}��G��V�m�$�����e�}	r~���#x�$dyK7enb���X���-!�\�x���+:A��?�Y\����[��=qb�o��_�.�|������n��:S5��}�����{J�Úl�8-�?ۖ���/˵��R�0�R�q6�����1+��p�h��2v��7�m�Y�9�������[!��]�a�Fq8l�G��j]��!r.�^�-��E�T�Hr��H{ԗJ^ @��BI:݁��i�F�+U�C�J`�5#3Y=���p/�$*A���L-�(�C
s�ʵ�vL��.ʨۓZ�H]�"�e!���i!�T�Hl>1�Z��h�ڏ��!\����k�.��z���T���y���I$�cE ��\�F<5��R����
8��!�����Ia�%��I��.���6$��ِ�&�oͅ�.�͹�*��3���L|��<[ i�Ą�A:i��B�.�ZƓ��'������U�� ����L����k>#�	'�!X*�4���AՒ[]fx1����	�'b���&1�����ܐ���=�!ĺ�`+���+�*֤?�K��4/�
y�C�Hdʕ@����T3�[C�K���(6q�4op$��<{&2�$�pN�g����/�㏝�7_����Mil�wWK2:�*��.�Q�r �z^COz�}9��$��9-����/��~��F�Y����J�~.����d���˜zz9�X�-�G���޲���p��ֽ{r�̦���OIU���C��
>DWn_-�^��$��:�[��2@�@��r�*�`Ĭp��@���%�	�2"n�`���mf:Dv7�ƎH �X��Zl�S1s`�>rR����W9Я�:��@V�)��YĎw��k�����/^}C>���!��S.0��t�&I��t�|l����M��!<ġ`$�1�ۇ:�"ā.	��V����>u��~o�����A������=��p���xi�As���y�h���+"��L�����4�Z�>1D�
y�ƒ���1���ߓ��}��o��SdQU/��M��9y���dq��裭^0bl�̈́�?դ���##[�~���^�/\�)S��r�"��&%����� 4JI|ôp6��iv̞[R�U.��u���[F��`MH�3��da��ņ��:Y_Z���7��ߓ�wn���1!��(k�R��O?�#ܣ>�^g��.�R�����Oeg��h����x�Y]]�܍��(��^��X�3���^�+D"�����=���5�ѩ�����/�W��|��e�~������A�cVm��f��z3(��t-�VÂ��F��Z�6=�bӳ`~��RQ�}d��(�ܸ{Ĝ�N�Dd��`�m[�Ǡ�F�$�<~NΪ��� 
r���x �B ?|V�yi��Cej�v_��Iy�'��i�n�c=1S�Ex�m����Y�� у:��	�X��0��Og�C:�أ��O�}='3�"�A+�����B�Yh�=�Y� �^����̈����f����&3L�,3qX/�Ř%_�۔gII��D6��;w�ȕ+��3����JO��3@u�د<����?�7l\���K�pG�I�Th�+`m�)�LV�ĵ�g�ƽ}������r���E7���P�/o��^�P�������\.�V|G�I\l��L�%^gq�e�;�����u9�ʳ�U�rf��]�L����N�r���nFׯ�)Y>�A���\�N���oT�� ���IB=lqa������cqt��ss�)���R9��	`����#5��N����b������A�-�S'�����q"e���A�*�ȄF�	]c:#\�GA�'7�/��;�F�±K������H�1�_�ѐ�X�(*��r����d��C����=���\��1Q�s�<!A�*�z8�5$u����~m4��VS�4"	-c=��E��#Y߃�@~ɳY�S�Q�H��L+��3`�#��\�LԱ�?����*���3G������%��J^�vHŘ��G���?��Lu����<�|A+-	z�����U<(�Q���/��ˈ@i�6���J7�HQ��P�9Ј�bxj�G��Y�����)�jC�mݖ���Փ��,����I��z�}�EU�'�4�^�	��4��Ԋ��P(�&.�[�h`:@�l��m^R��0�dkq��4��f��!,ϵ�ʩ�&$e���e������H�~�(��-YY_�7ԃ9"lFYb=�JA7c_�~OC�EL�����zJ�����e����D��ؐ�h0`���~��d���;_��x9n���D�[��5��tZ�+ �?�H[�T%��!	^H Q	��2��M5�zOmLҫ�_"�-�YN�M�n�}v6�XnO�3��z�؞�J��č�cz*G���@�]��Թ���i�����r��M98@S�D�L���R��nm��on��GzL.�������e�P��9�zcY:��U��'��L��c�k"�zM|����ڎ�T�d��%�))����(�vH�*���4̻����Pʃhv��k�G�@��!x��F�2�J�QqU������!�����AE�z1,?�0eF"q�)$őK�$����2gY&q1d�p���uwkG�+�٭{R�]h4��ʷ���,����z�Z�&ii�}������$)T뒿��l�e�2d�hܨ4P�xjg4x�m��� �ø�"X���Y�<�TKa�?v�����Y���j�w���z�]�v�=}n9��I)�Cw���t�#/T(�Fl�����oʫ���g{���]^DG�ݨ>�L��NE�-:�s�T�/v����'��Y�m�(��k�6dDN���H��/�bH�>��_b�Z�S�k����h8�fh��:�cȕ��k���L�ͩ�Ǥ�_I�񌦟�x�J���i�@��E%=6	P]�7�u9}�@:�{�V-V�8��i"�%LB�D���8~L������R��U#���פ��7�'�Cr&k�z/��z�R��\�~!8��a�1�.�JR�*Kab��F�P��кǏ����o��6��|��P8qQC:��֒���	5{�d7��xf4<���6�FčzZ�$�Dfބ�?73\BO"�K3u��8��$h���Pnܼ�FeA�
��ww�X��� ��L
�N���-_�wnߔ���(�͠�.�q.��q��L0a�1_;="�x�p �B���Y��1t�J�l#G|�d���<�u55l�Z�v�V���Ci�������=?fao�qv^q�Bj�r��g��vuc74+�������C���Z_Y��|��$���f��{���� %�+�(�9$���?,�9(l��m���4� ��-�xU$��Y�8;=�jUʊ�*�A\QC�rlS�z��nN�����,�e!1r��8�����5��s�%���LH|�}}}f�����b�Z���:���a��#�$������ϴ*�~��0ˋ�J�В�e)�")�uu�1��:���QD��4Q����*��p��_��¨�q0�A?{�{��<�,p��|��	�,�J�G��;���}/������]�c�H�	��3V]�o��@���;���>(����8,&�i�$���<$�O�PJ�<Hi��XBG5Br��i�ȗ��(�N��?��Q�o]�!��E9��(7m\֐f��Z�ٻۑξ�����ADu�Ng�^� k�k����e��I@>؄`��'�7��
�`˒+�BH���@A�*��N���j5�J���kþ3<N��XDܮaF1�%����X�{-Ɩ9������y#�v���GSV�/5Ec�|Y�f_�j��p��첁���
g����ݬ`�z�2QbJ$3ju�C<�M��¢�Ԕ��@k��L4$�!��T���= �c�Q`�!O�U�5C�`FX����6���X���6-�������@k�ͪ �@Ѓ3"{j4�d��K`|�����k/glpN���͠���?�ْ�܄(�����H.'!jl_=N��7࠰�9�d2������}��I�ސǾ��ܺ��J���G�ѐ�"����0��T��d3�7E�)s,T���F�:f��r����`<���� �����DÎ:��ԀC��1���:�r�I���jIlJ{�s�1���#���)��rY��9����g
�"� �0Cɜ����cڐ�h|��d(;Aa�w*�̅$i%Ɠt���X�i����X�8�zqr���7ˌ��ۡ�^�W9$�ug����n�T��E> �f�4j���BC4!��$E�/�\����y��\����v���q��z�S������N/d�X�ze%��K�X��<*�����@$��H�e�����Yȕ�+���5.G�7�=SG_�b=7����
�'y�Re2I�<ː$��Fꦆa�A)����ᄼ���ƟsQ�	4�IJ�����y�g�j(Z�m�#�Ѣ�jH�S�o��\��J���o��g�^����C��.����Eٯ���s��D���)�������c7|�*��%�(��h�"'��E�V��<�J������<!��.�����E�v��{.0�8P��O�al�	S}�p����̛�{4w��P"�h��Ƣ�H�#<G��ݘH�<�a2v��漢:�n�fOT94IBV�����P��/���s,��z��'s��X���Gno�����o��i� LW� 	�����	E��
�0��d�k�Px><��j"o1�L� �� ͱT3:�k�����n��Ѓ����D-z�ݔn~"��rB@�6�ΘL�v4��ٔѰ"}��[{;��4��Sʟ�[9ECΘ	
YY۔ZC7��:Ř��ϱ���,k��ژb2�Z��2�[1�T���5$�-�����s�{��IA�O:?��������cT��F6� ƆLS 6�\h7PoSг��go�),�����7(]� ��Qz������$yZ9����PN�!-�rW��I�b��F�7�"�K`Bv)��'��!F%!f̀�gQ(��B=����Y�8�ԛ�c"�+Uފm�!Ld�kj�~�ȍ�H^�[���{e�D��5�`�NI4ľa��젭����r�@N.\��HW�MEO��S���q,������1Y��?�ۓ����(�Y�iP�eΆD8�.����
�S꼆�v'��q������j��,�ȣv��5�(P����r�q��$AM�;y��Z���(�� ��_8W{�{$k��s���R�KDS������*1xA��o��,5ɻ���y �.,s�s�V�H�G��fh`+!�;�/�kJ'7�#��z�̎JP��%������^pW��z<`�`l��0|Z�`~d�ؤ�LE?YP�FúC5��!Z�!�Z���W��t.B5�?���ؐ�7x	#ES���`L��c�����s~QV)Y�՘��r��"Q@���.E;�d�^W�
1>�-����K�8xy=؋�VD��9(sSa�Ĥ$r���v�Ck�_@��4�\0Rگ$=���$k��/
��R�e �jRӧ{�z�67Vՠ�m>�ʂ�ؒ��\�OKb}0N3�$���*OV�ĉ���R���Pע\_�� �-��M&�q�5�wkG��+P5}~��1yf��Á+a�.�;���x���ז$��Q$����h�,g�"(FtC�A��}b?����rD���E��BM�{=:�%��u~�;��42����	z_EV��a7u(&�q�,d��6�_T�L��!���wM3�@��sg�0�n\��(��Ԡ@�({�t��J�f�]�[���
M�X��ת����1�`|�����W�Td	s����<��I<&�Ī?Ahe-����DlL�q1�q�����Wá�S *�F���\�XR��щtc���P�܉�%��1�0q�8 �%��
��8H�FٲVӍRDx05ä���gAcspPj�����5n}W%Z��WJ��D�T��#O�0���b�+�ش��
����/x��<CT�Fr ��Hp6B��++�z�Krb�$5�ǉ<�:4�Ұ�7rb��]�C֩�NV�ݭC)A�1�C/�tl��1T+�"������?�V�|w3p:h�/�(�i�V�J���ఔ0�S�5l��҆lnn��,Scf �=���N���L`0y�D����;]U�o���c���c��f2������X��� �E4<�A�H�B$���0,��6Fu�����؋4U�)9aPa����"%1ԛr/X���Y��q��/!`ʄa2���G��djW�H._�P��{O]lM�f��*Y-?`�"�;��r�#�5�A ��,5��3]�T^�χ[ ���' g	>1�Ej��	E�0�
jZQ�VO�{R]Z�J�?;h������@��9qSːC���2a�^���U�$��af�[�p���GN�F����y���EY^Z #�7�.�,��5Ae�G��>�LI﹦����fW�-hV���Y�5���`��T����}��R��W�Ͱa�=Ԛ:��|��#Ň�,ٓ<�gN���'O������Dd��X�cuO,�v*��wO!�5K��m($���h�����r��|7�۹'R�����A����Pt�^�sW>�vCήי�#�K�GŲ,�����YY^&��jZ�K��#X��"�����5�C�H���ߓ��e]љ�(����p&p|!xo&��P=��g�n�G��CY8~\^|�˲��1���ͻr�����U�r E<�Ø�rq)O�;�|��C{�/��e���l���EG��_q�h	{I���9#�^i�%Uw�����X8�"t	��U�89b@��Tbŷ,�!�m�#`gA�Q�ĭ8�,�f�AG��ꊜ?w����ĺ/�~���j��D+J�`��v�	��)&����w�p���T�m��ML�Tϥ�7��F,�Jf�Ñc�q"cN�˻r�%����mݦjp�V����{��| E[�m���U��y&�˨!L�,P�aCI�Jʸ�kCv�v{|��b��2|�,�����|�Nћ� �,��[���0��$nI����Į�Á�XXdKˁѶ�H�~
��~�(���2B�Q���&rOpQY01 �B�lM/ǜ��Q��#x�=�㒎�4�<0<S��C�Ք���\|�]9�o��Ʋ�ה��sE�9E��ג�ē�^�R=+%�������=���"&�ȲE	���{V����>���:�<j�R/�q�
�L��B{O�gHן�9/�=�!_�����6/*C���=ؑk7n�ۗ>��Ƣ�U*�GY�I�?����3����~8%�3�߸���cKy���}���w�0���F��x��,|����đ��t]��0W�1X����X4�e����b�H��!@
peuUΜ9�M��/��Z�Ƥ"�"x�06�Z�C��|zM.��k����	8��+��_�;���� ������V�(�>cM$!�\��j�s}K�3��� ��<bkE-�c�j(��Q��Q��Th]�M
�����WE���+w�ʩ���G<hm+|mSe��nc�����Pi���I�7�e��=5:w�dMBQm�R�L��B�يg�ϵ�zz8�17B�N�OU��~�>�_=I�T�# u��=�.�X=�N<�uˀ�T��>A�ƾjw�����
�fд�]�}gK�^?����V$�'�!A��s��Kaz�C
�S�dʡ]sZahJ]`��C���g��S_\eW�a�C�����"��2���tz#�ggh
ǜ@1eҾ�i��D���^�Y���Ж"�ruY�C����g��£���~*�?���0*8T�Z�{e3�� )�?to��sД�ʒ�X?)ul#�/��㲼yN��/:�r���W/���[�veW�8�<=T$���b�&=�[�J�H���8���ߤt�$.������r"a5�=��U�b�� Z8Ҁ�8���zW����=� W�B�\Dܘ�+�9��Ut�df4R��>�ؚ�P����	<�`8�v{@r��$�0|	:�0�*���8�#�T��G	���㭯���ʊ,,.qV�
c�I��A�Xd��TN�K,������S�:#sbJ���|H� ����H��أ�Sr�[�����ύ[[\��vK����/������>א
��6/.�Ɂ�ޱ�u��l�v*��G����ـ�����wde}S���o�'ׯ�/^{��Aq��"��+9u�ȍM{��"in�����7n�/�˥�ߐ�ww����tD{����wߕK�c�P�u@�x��)n�`����#o�jd ��XXaXE�\�z]^��+d�~��g�O!L$��D��jb��69}.�jA!�ax�u���=����E��'�~�Gm�������
@&ۻr��u�����G�ٵ�F<䜠/�W�Z
6�(67�����׉(�-���'y��wd��@>��*v=�Bژ1K�1yĺUbIKt�/T��V��G�/_C*K���qB�/��O>.�pN���<��l5w��W.�)����"�������!2@�:���Gy!=�w.�4!��5ϒ���s	f,��Ri��e1��_J�H���T���x/C�'?� �A_�;RٱH5��G������iCXN�Ȯz�˟^����j0�v�����{-A�U���l��3V��b� �I@mrW��FKw��(�B�0���YZݐ�7�����5��ӗ��~G���3��n�
���ʑ J|'�dm� �t�=7뗍پk5G��4�U=���lԓ��]]?F�}��Mݰ���'OLz yj6@HI��ν�1Q�\��D�d���WMM\�Oo�����A�'v]�|v�����|�M��aK�[� �g�6Q��V	sec�Ѿ�����/���-����)*�Q����u�ˍkץ��E�߁gT@�|}����t�9�d0�n���-���D5��O^���z�s�1D�*eKÈdIb=�@|�E�l �� �8S�S��(Q���I�٦�v�[/i����`g[�P�'�s��ܻy���s�3g�9J$*�O	F}{gOÉEY[)[#�k)�5]���`o�z��g؅F�Q��^@� �;q�Czh!/pZDI�������W^W�Hfv�!�OI���w���t�����{��C�g�|J޽������]9h��gH~a]r^��m2c���,�e���P�U&1����km�6��C"�A����I֍�6�#-^�3�4#4ͪ3I�F�.˹�aU#�(sxC��~���
Q//��A��g����>�8K�2'��cS�*R�y,��Y��������9ЃW�c�	�K"w���My��w�Kp�|���hjð,�m�N�飂�h�sÚ"����#*Cb�|z��Ï�ʇ��R�,�˲�� =D�ޡ }��&��c�|�g�UxA���D�����$���#�z,K%��-rB�u��w���PP�Ί�=1C�(�������g>�FBmlc�L���aO��@���@Nn�0$�,+��s�m^֖��X�IQN�rw̲-�YG������;]:%̭A8�$%�c�������؆�5k��Ø�(i��	J9�,B5�y�8�c�O�7�;�}뮌�-i(�[¨V̹����S��J�K��ES!�V���N�}E,�_&-}�@��LC �++%h�K��{Eщ�j3!e"���B�{��5��0,��;��A��Iz��q�(
�ٯ?�c��em�&�Ϝ��}�99y�<��s��ϲ%�Ν{�Ln�����l,�&�=9Z4��I�A����g�����Q$�C�2��v?˷1������ҝ.��٬���d�ĦD�^c�a蔶�[c���;�Bw2�1���Ã��t���	�[��,.���W��\. �D��1=��tq�h(}��c'�lwq �Qh	���#�2͜:X�P���M�8F�X�̸���L�)�Hj�b��w�-�AK=�z�.�h��9/'O�d\
O�#"h�h���ŷ��v�Mp���}i��7	HV*�lE[c�|���B�C{W¸�v0���!p�����tI�D���x�Q��p"�<���ވ��L�!�F;{��|��}W�|�e5f`��/��@�����壏?1N�zc\P��ӽ�P��P����Y��A��`?/�%rLf��2.'� ��"C�*;ccV���w���(a^�z3����1�#�v]lT�+_yV~�!2��hbV�5��>�,����hM�����\�$fEp�p-��@(�= &C� �Z��p�Ú+-@�F����޾�Z��"˖���p�9����jȡ=|3��s���k�^��� ����\���k�sB6Ϟ��~sY����e�<< �x.�Iu����zZdI�4;��,%+��<c��|�7N�����l�Fz �ss:RZ�oQW�Mɱ��r���6a	�_���;0eّ�i�u�H��ۓ�Q��jTy�D+ND�Ȧ��+_V��kWQ�T*)C=��vK��%��s��}O��7�*a���(P�BCb�b���WbB���ʡ�NE(�c��c�"3��
�F�>�O�z�����mYY[v2��M�S÷�X�p&'��H�o��%b�~P�hi<�����)�nD�^�R���?�Y�ʏ2#iG/�87���`2G�v�Y؈����šb2�ZFbL������/=.O>��\��}�����������ۊ��z8�,gϟא�1`!�4�0H׻��IT���}M>%��0o���N��D��X���/>�	s�4s;0((�B���h��!D��R$��G��xk�rY��g��ug	U$\SN�s�U�&�ڂ�][��4>�=\��^ts�rj�yM���B�{6�+�L #��!�WoH�is�:�0Pa���c}ط��ց��^��w��)��^8-ǎ��7e�2sޣ΋� �Ȍen�46&c�R� �C����6 G�f�	H�aD@������7��Δ���|H�eh��0vO-�"Fd+���t3�'�üY���������m�e]��~ވm�=�H`�%ҵ�O�r'�<-Pua��Sl���L:OMa=�EҚ��*�~h|�%W�X�xf���V'�,l�i&�O�*Md�;b�E��Ѩ�qd2I�yϝL�W6嗯��d�7��d;��'�]�D��{*�N�#����82�*�:����d�l0,��%�91�c�5�i�\�tVP��<Nl�v�!\�)"��r��$x��ј�C�B�����}�uc��{�ͷ8��hd-{^
�1<'������������� "�c���C��1�n� ��mdlk��pl��@2bRY<��HK�P#k��n�s����h�C��	E�0�01=�5��}Y[?��D�B}��`L��L��H���gXD�U��\��ikh���K*�s�%U�kv噲s���ͦ9:^�ˍ��t�ܑf{,�Ʋ�I*E�z ��g%�������3��8�)Ϸu��"?��7S6c�rfH,�с���dp�D����Ԗ�J{K$+Ŏ�<M|���\�\H�*iϘ}+��Vr��p#����BY���k��7���s��0�?F_����v<E&a�BC��lM�$��04�77�,����L��Dg�[ss�`���~��K�m�jc��4��HmTr�v�8
4b7o�$K��?�?����{?}�g䏄[o�߳rl>�~Ti��E*5��M|�`�T�
�ʬ�1���qwĵ%�vlZ�M�Z�5�'����\̙�=)��'<�8խث
��!sf�_��|�(���O�PD��+j`&	:5������(�4=�I��Y�^ �= �A�Wa�
_	�@y+I!�N��<��>WT���}��{R@8���ګd���\d.�K�A�e�hB�"�RS=t�<������;�-&��B���t�u��'W����9˵Rٌ��RU�#5��J�c;�D�yr���2E�g*��&M]���ט�碼����uoO._�S;Q�H��Ϟ5�n���(b��t1W�cJ;�Q=D��ݦ)����mA�:�gk�u
p����Ɂ3wi�G�~��'�W9���Kb/�sG�l�T��DHBvg܂$qeʹ���R��(3n6��U9�~�BY/Ѩ�j�!-�)�O9��G�"��@\O�K�"?0���eX~B�$bx��r�(��صk3CB���1�R�k�����A�ݏ�B}��4�c;�X��� zF8wm���<���,J'��`|𾼯tg���߸x����æD�D޾tI���]��t���x�,ˢ��mu�A�+<��5ޟ��v����dx�����Q�1q:�µ�\�!�	���3)��zӱ��ȱ��<|��U�b���H7`�ח{��r� d #5<����=O��U�0���5���B�z��	T���9t�`�*@^�}l��[�����7Z3�< ��b�
�@`r ���Y�-��o�'o��6�^�܀��_��g����M�y���{���p �Î�ߐZ�N_1T�ssu<�rwy��(��6XKQ>���ݝ�j<nʕOns�}ޯH�ϵ�Y�%5L�Y��P䣀j�		�P@��b��]�)���-�!��j��pnz.���d�4͋�D�8Ii�:*�I����%j�$ެ�;�l6oH�ȑ�P�����I�K��.�����t`�e�ۘ$!��������/0��I�{l#������i}	J�{eT4�E�CƔD��H�c�8�����o_���;�,�K\K:�GH��)��&�����,�,I�}@��vw('6��������E&!�z�Y)�*4ܗ>xO���h�z]�����z�
�Kn�j���z�<��l���mR�Q���T��3�̆JǬ�@��:������?����#�O�d[�4�p�P{գG�����ܡr�w �ޡ�@;F�B�V�Յ��NF4 �4(�5�ʩ�g�'�jZ�>7�b�ėa�#5��&�����"����F>!�~o�w�R;:��(;!"�y��ò��̽��
x.�O������O�s�DdPO4��H����,4��t�ݙ�~�1"$*NS����M�9����y~��^�D!n��ȕ�!��#@��U��"h�S$6����C��:*�Q��l��%y���ȣ�l�L�!ly6G�3/��,��s��|8�&E�#{/��nDʰ�NVd=%����Ϧ��}7���E��AoϑD^ ���5��=��B+��B�.6��t�`���YS����Ē�S]h�V!�<�aI��$q,������˜w�h�.d+��7e	��vm�'<�PF����?����Y�n� ��3���� � ߺs[�b`ܜH]�?B�#N����F���@�%��W6w�s��&�c�|�z���0\�`��k��R
�$����3ϩA|Bn^��^�]9P��܃^˳�=#O>�U����ƃh7�@���K��$F��k�c�'���b�*J�9y)RLz�F���P�s7�P��k�D3��qc�{�1����P�~�+����{qiQ�t�8@��_]�_�L>�zM�gAC�,.���px��۟)B���Ɔ��]D}��)��qݡ����*�Y`�CR���:�"�9�-c�w2%��4������:��0:	�ZC��cmO���Pf���	N��g/��h��qA�L�==�i�L����K:-��0K7#���␆��G+pFB�8"i<���"�L��ƑS�ƂZ���>�LO8��n�D��M/'%A"�^��1��BS�2kX�3�9ȁ��lȒSr�����@�9��Nxk��j�ﲢ����f�Da���5y��4��.}@:3ʠE��=��<�̓Y0���xm�ön�z�&A?σ�Y��6x�	��pBٿ��+̐ 7��':l�1$�V-1� :=�t��)sMK�zW�� �YXZ�J�*�A�eU���g ��-�̡Qȹ�j�0bR���1�7��1m�Kek��:���r ��2u�G�0��	x!s����-�*��S7�����;w��?���Dx"%�>�u�<M���TE9���}oK`[��4jȍ������ Ka �� v��8żsF5��T!ۓ�^U���O=,�>��l߹&?��?ȭ{;�+2�n�"�膼�îT
��^�р���ga:)���X�����`CG�g0�V�}΂I0���j�����͐`�98c:�i�d�x��evi������o0��U
6x�Ù�3��` �!�=�D���M��}��`�z>�u���Aݥä�ʚ��b|��#n{���eyV��ѧ�n��,���7@�ҍR)G����yA����j0��|U���wM��KlB�S�ٔ���1�	�����/�#q�R޸9w�����Z 
A�&2����t}ܚ��"����W)BP/X��Vh�?�U>��������}YY[��g7�܅�d��)4��>��Cy���N"9gt|�;�z�c+�dOAU7��y4/8#/�cpJAc��D� ��@f(�n���ĥņ�r6��n����K�[hjE�X cp|m]:�C�s���S��8vL�|�i����Λ��\_iH���l�G�#h��5�@"q:"	��1�R�%��Q�GϞ�'��ޗ����+�k?*�<{F^����o>�K_S#W����kp K岬_������xIC�U�?���[>��-�b}6o�Ag�Q�3�给?ޠ��)���M��<V�R���a��o�T��#s-�����>��^�����9�>aD0z�}�T/�������5đ�D��!QJ����Av	<��ھF�&ݡz����}f�1�	@����;��I
1f��.9�W��6C;���Mn�=�j� kKu&��0� �%~Y�7o�O_~YΜxH�M�*�|Ί�{���ի}��˜�����G�7��&���,7겥z�NI����T2�W��¥q��ߋ8
Rx|W�3Nn��Q*Z�h�!B��&�Q��И��O�=nI�嵑ܺy[�="L0Z�=��W�� ק��y4�Ɋ�/���\�lK.�ئq����l�:��d���s�Y(f�;m&T=�SC$�Ua���S��}�lݻ)wo��C�% *�2�����⥗^�Sj m���`q}?�*�{�m��V��4Q���z�7�$��u�s�z�ays���ѣ^Xq�G܀6���U���T.�۔����FΟ��0p0n��Wk�<��G���M��������,���n�o���?/�<��,6t/�mȽ�6�$�"5t���>Ef)��/Fb��_���=�|.1��9&2^sxi.�$� B�<h��� &�l�Еx�Ī6�k�I3��Hˤ�*�1³�ЯI�y��1�`�n�.�_$��C�c)rRy�1�p��M�[.%��1vh�׈�
��Р�������ի�8�.+��dKck��efL��%C!�!%V�e�I��S��컛7�D<���99�\���}�]���=����~>�g{�ζz�YY��vI�]�"�����oɆ�;��O��2�<�*��(�!���5��?���ˎ�������X���'�o�E-�ix
J���U��o��������/�Ǘ��z��c,�z�',in�oȗ���,�/QJ�V��H|����l��׾�U��%�|�2�m�X���V!W)�7�����~O��'׷~,�(����q�Xx��A�BD�L���/�<	�U�Ԡ�5D�η^��O�[o$�s��`X<�YW�C���[֌�[`��007uoݺɊ
P�X������+������~\�{�Y9�{�׿|]�6�U��f��$�.�Br���P���C�g��}�����6�-��'��Cj@*>��L�>��ʱ�'��հ�!�{}��k��~�����AQ&��hD�t�#��B���yv��.�l�e:��(�|.�d�8�5a��I'�oꞳ�����7IZF��AO��0CJ�� �seaA�ß��z�c������.1���2�|�$E����E�l\@�➤�� f�/�IMҊAm?����?��O�/��|�?����.(`��N��d¤����gy�x�^�>=2${L=޿��?�zA�}(���W�f\h���:�y\���Kr��y5(&�׎3���6qϞ=#?��dg�q��xPʳ_���G䅯>#�~_.rY^����P�o>�h,EP_�uM�	�ͼoݏ>z^�H��b].���"�}��� (�ר3����<�'���_{�����s���|W�]�����S�|�ӫ�N,Շ�y;g� @￝�����9}R�?�%%]��T�gl_\7����. ��$��9�k�u��]�9��<�,�ְ�ʢ:�id2���{���]^-�&BL:R��t�@�\��6��{;r��5��ݕ�����q�rlmI
H|�[��
�'�?1���L���g]�S�*�{���G?�g���^�3��������p�A�����+�#��k�;^����@�z��5��\���c9���ciE6���/q��лIS!p�񜽘1V�����zЃ�3�y�\���-g�y�%b=׊-΢9#��-Ʉ�����?<��#�?��T�ܾqU~��m)T�#��t3դ!`LiGi/2H�D7F50��n^P�4����)�����!L�����g������c��m��?�1"626[J�K��������c6C%�x �miqA�4�.z#�<��^�]5�%e7����zJ�����?�	�4_|��5���Uy��9P��?�)�MC9�MxBбseH-�eU��=��vj�C���A�6?B�-��A1b��/��}��Y��}�na��!Q
4�dcK���]�W^���>|kG�����K_��z�G卷.�J�8ż�z�j�&'ϝ��!Jx�$M������;�f�;z}P�OL<<g�q .t#_}
�J9��c��%ʅ�V���TY�M0�\Ϥ8�dKV"b�xN���ݭ-�è��a<��E� 4����}�k�[���t;+�Y,�����"ӂ�v[�F�R�����ɝ��ewg_Vj�3���~N�C�1��w>���gr���> ��%����=�~���J��\2��vt1���1�=e�.�9��\b4m��/0!Wc�%Ӳ���(���i26֥�'m� 'h�kR�z�{G�i����~[�8pH��5>�[��|����h%��('6�S��a8���=.cE5��L�}�Dy�:�3�	ih����B/=�)9�B*��Xȓ^�x�lM�ޣ�m��dKv�����Ǖ��o�m�v �0�c8�4!M�!)B��_�'�2b^FA��1 � ��}��[��̭�}k�����M��F���f�e����ߐ���O�ރ��]ln��h]|���N���?�����p���'?����)Q����O��DH(�B� X��ZLB�C{&k�+`�s�����*|Q�[T(�A �ń��Ź�F�8������������%�d}�c��_�B��B����<~�����?H��H1(I�9� ����Y�J" ^���l���q���2*�E�6Ѩ��q��xt�00�~+YO�(�����:�.M������fXP|&m�M��:*����d%t]�i���$8╃�тvg4�w��i�����s�vk�5�����/�ݟ�i����_}"�����w����_~*�S�6���$�`��"gEN.�q�"*�� ���x�N%'���k�ʵB��\(D$"D�tIϥ����L�|n�tn�X�p�b���9�B��1$�;�|c&i��)=D�(PC�!�F�=�)�T�t(�+'a�6����4��Os�~(�IZ<k�h�aQK�;�W�~(}W�[k(Gϕg싨��G�Â�/� <�61�1`p��pu6�[�-�'r��O�?�տ���C��1[��&W �-S
��&M�<Ee/�fQ*ζɥ@'9�'S�iC���h�̢#�x,��ˋ���
��YRG�C$���`Hp �7uJ��>|F���dS6�`��z�v~ ?��ì���~��$x6)�ؼe�I�on�U��V �� ւ��4�`C'�e$�hV�#U!�>��wkpN౧@\c��y�?hhU�j�߃��x+h�2*3ɦ�N����I��^�*��-�#�I�[�p([�63�X�U��/�� ��>�4���A�ֶlo�ewsB����$<��[����QР�O��?�_��`�تY��XWmR�'O	��ze��N��>����R�3�&J�a��:��G!DJ�ozŐ���oC�8F�O�)]�H���聘 Ҹ
�������B{��h���7$�m���)7�,��J֧����FM�mb���Q7Fh��%�$]��%�f�p�AZp�(@h �ղ�
��I2𿵚W�F�����>}�q"(�K�� }���\�gI�K�$A��܎���7�ƞ1� lN.��#�ld�8��D����ɻ�~G��?Z�$I}� ����ft�07 �����Bd%�
��c�TxHE�N
�i$��ӥ�+�����f�	��R�UT����*_��NZ�O��f�ǃ�C���\߾�{'G�'�����<�H�-X�$�B,)X���K�􆫣���΂���@���dH� �$��@ ���{Mn��di����q9��$����;�tN�8��I N�z[KV�x3=�����b@�)0x^�S��K/j�z	[�꽳��(u%(*����{�#�� ӣ#y��X���My��[ɭܕ����%��b��7^���_���'�|����
��|r�|���6��h[��X�p]��$�� X�Z7�����yE�D�% �]$Eq�V�كL�(�m�a��F�Kǒ���.�"Sd��j̒�/�t�a�b;I�t�z��m���K�Q=M.��Nr�p��	1)��8m�dVn��&�M�3��ߓ/~�QB'r��մ��� ��m-�xI����t��8�V3z !��D��Ը���B�t�r^�TIx 06N�a��(��y��[i!-�zzN��ǘ3���5'��6�]ߐ������ӻO�Nc=��K�Vg�jAX5�������SA�`m/̼����(6A#.�ݬ�/��	��76��G�$���6�f����4��b��w�K2 ��,)��Ϗ�p&�������I��D���µ<�}��{��wn@jM���x�_���T�T9�.nE۱�E�H("�!~���W^��$����W����:Al����D�O=JB=Y�W���S�k��3��e��DE1i4��6�]B�Jk|���c�gj�g`G�\�o}�+ɚKJ�p)�n�Ic�2p�cS�k_�۷�0��&m��{a�s]���L���������,�-Vʯ׍\tT^�Qr�^���I�	z
Q�2#;8-D�ޏk�	�LGjo�Ҕ.��k�,A'4�ߐ�-4j�dH�e!��1��#y���gIK mz�+W�˓#��[W���;I����IMn4OB>�֊��i��h����L�k�K�������٢���C��ψ*P�l�	�,�W�hq���w�0lL�)["�"�r8�Q.�ͧ������?��z$����u�H�c{k��L��븾�"5?y, �G+�\��<���,��.�=�G�d���j�p,�?а不��X�2P��4%��X�x��X�	�2L�U\��pmSF�-�L���A8ޒ���
	�Cdkkm��xD_�0\�a�dM�r�����-�G̖��r=i�Q�����O�T<)�qհ|�Z�1B�e�cB�q����uPA�E�� L�4��l��kZ]5�;o�Iᰵ�M������x�x}[�ӿ�nޔ6=��8Y G����.���N�=��z��=oB�
�F�5ڏ�8@��;�c���C�`oM&i�7�yE6; lQ���T�x���1���w
���d�o&<�dĔx��D��G�+N-Ni�����٠� 4,����kZ�7��D�H�UϱZ�#�� ��8 R��x�2w�0���F$ҫh�(
��k �Fw�N{c ��	���>�h�}���$3d �t���z�������$ �[ ��Il� �����`�"Ia��#�=�ntE�۷�	�!Zʮ-!�F �&��#pb$�S7ɵ
��H���Q��SKca6HŘI���iH%�h7>�h�э�j��<>�#��� Y�5i�f<�ە�����u�eC��EZx'�_x��~�y��:�0͋)xM�6ٕ��M��m%7�ads���7S����t�S�l4���JZ����2�ǒ[3�b%�'u���:�L�Ϟ��d<FˋV�]g�x��Wʣ��1?I���L���$ 5<U@�'@.�3�����)�_B	WWQ�T��2��-��#������>��/�|�he����d��e
T �.U��F���7���jV����#d���s����s�.I¸��QZ�A�{h�Ť 6Ztz2o�o��}yp��E��;�1�zP�9��~�={̬xK���8H����8D�DZ7����_=W~�!�#߹3P�w����N1a͓ )RM\�&�5��P�`3�vR�p��*m��"�`ck��tm��E�a6�������&�|$��ƅ>W���Z`��@t���CNK��ʅ)���#6����b���iq�<F�j�\	`�Bl���>"�bӆF�m�XP�#�����!52�:s���!��;9�k�7��&!u����,��S���I8����g��܀��~�p;9>�;�R�@���������;�>xx�)�v 7>�ʳdN����m�ɖ]u�.Ay�o���ߺAiuV@�*��
d�ƃ����u�:N�����82{�1Yg�)���u4��O�?V�(?��g�����������[��\_<L��Bc	��<�}�*g�G���e�A�j{{�ZEu��>��~r�ޗ�צI�մ���}-��Ԡ\`�_����&�q_�ɷx��_�1Ƞ��<|�����I1�u"c����ϒ������z����)��|��'D��� E =~!N��k>}FNZy��-�	�[(@ ��91�.�X�]'gĩ��|/0_ڴ`�=�x��\�����>%P�6��/iz��g��
���379lF�],D�c�&үSj>�WMTKŨ	X���b�Eam(gi�<�ݤAP/��'����D� &r��^ܗ�����!��o�y6�(D�t�5ضK+��=��o�ڪ�}�+�9H��iի�X1��:4������ɕy��{(���O����'?7��h��nڔKֿ,�I�M�=xS��"==���m�J.�a�BO����J��n�p���(�e��П̬U��Q�~�i}�;ٟ%�O"��n)xQ�������DV��&�����)���<bh�����s���L`kr|��Ё1�����e��!��d��U��K�7��W�\��ׯs�P�<L.��'�dd��;�W�\]O���~�L�?��m����I����S��Odzt�Fk7nߑ+�o1V�J����r7&E��ڪY��uok��f��Q�RHo>�=��&Y����Jy��,�x�KLe(~@��!�~�,XR�BH�\�d��\T���/:�
 ��ts_�[��}��f�72 M�W����$ä�)�����6!��6v���Ce�V�5�M�����m�7���"5Vh�2��9#���b-���%�����L ��ѓ�dlh�ᰣ~He�?H�As��AZ�vkI !#���S����y��m����g7�iy|x��ںY��݂!��v��2&;H��F@t��;��k���%+�.~��������˽/>�t+-�o}�]��7ޥ+�l�,ϒ����/�h��&y�ؕ~��MV\r���L-��ɰYQdH��I�)�Oݩv���P�祲��]�|���̓��4��͔�JB`0옥a����79NH�
����:�*��ޓg���`.�d��EO<�o������$m���I����K���ꜵDTB!�'n]�~P9�Y�q�@	<���=�A����o��Ύ	�Gv��_Ɋ@�����m�ؾ"{�'��ɡ��ݐaz��ڀ��_j���N]��X� �C�l@��"���+��0��Z�*$�L�DoN���Ȥ˵�j�q�r�iŊcS�5E��A!�aq����!["�+�G�.���M��,X0Qal4v��\��{���Lr�Ղ!IM���r�\����#��o�o���l�\�_�f�ף��Is�W��	�\h�=M�
��dil$-ؐ�����p}s=�z�i�����20N���Um��pl��~�n*��sԿؐY�T�t3ψ���Ez��$�L�6�j@��{w�H�o"�o�d/^�7 G�t�����Myr�D~������(�����҆LL�q����D1@�5e���Fr���ϗ�-I��>��˵ D#��H5�&b�� ���;��7ohe5{'�zQA�&Ћ6�qI �� 9����L��d���i��'I�nm�Px��ڛIq`���5Q����T��D�Q��#�ay<{���06o���J��{#�v~�������K����d)��s�s"�RwS>��)i�K}~��<�;��׮�p�l������efN�V�_� �d�D��&;��V�e� ��5U�b��'��bM�����,�o���D(�Ҝb>�%b7a���ҙ^��2�R�&>BӨq�`3�4E]dƥ兎O��[��PD�����i�(5�P�K����D�%�mm]���>�gU��Wek�(�!'V�F��Me���	s�A�Ǥ��%�i�γ�c��F�*C�"���cJ�c"b䉞��ڥ.�s�E���0}  �{�,�d�nonʫ��.�n��!�����R`BCw�_��y��N�o��E�����-����73I�5���9f�%,������Qc�����Z�,h-��)��u�(�@�s3	<1|�f�����ׯ_c�@�CY��
M�~5�H5,\���(	�({�- q3�� ع�.4K����YJ\ C<��ilU�w(UY��ln�o0�7�VϤ�6 :�(ysXPhO��K|�"�K������O��Ӄ�ژM�'isY҂\)��Y�Ӫe�4T2��I5����=#j�/�����S��Y��W;'�Bx��њ�a]r���%B�P(Jd���U�Ȥ����b�~0R"�\��x��f���_���i)@l��e1p�r{����ӊQ����4�01��_H��c0	����+���ҿ_����on���1{��ɭ�ձO����Zf�`}@��^ٖ��S����vgk���Z���v'���g�xK���
Bm/����d�M�0�i�����^��v�*%<����T�v�|�+o0����9x-y���̀|�ٕ��^���@~���t����ՂsO&k��A���F�?��1?�3�g�q�О���E����$A�3���[�ӛi̙MH�r��˜=�=C�	�jh�GP�;����da��R\
,�YzX�
�ҳ-�u��B|nB���nW���NE��?6�ez|�I�	��!����U�s 𻖬9@�ge�v�E���	�f;)��O��G�����#2s^ ����1^'7Gkni҆,�͠��YfD�=���ViAY	>`�J�KŬ�L��Y�L�*P*.]����S�^.`=7t��V�ǎ�B��� e̖H]�,�4�u�Y��4ȸ@;,+�6��.A� hƑ�>�/�,��@.*�\4͇,�Yݢ� ��^��N� ��A s}���~�%ٙ������$��z��C!z���#����� -�{�����}n�A=a�4�k�R,���q���sU�6&ZV�<!Z�;�����?��ț�_IV�6Ba�`��E!��+�ʝ;���$Һ�3��+��bL$C�^m��	�I����p\ �֘���]r[��4]�.gE<�4<#[U�j�˹�^�X�2o�gx)��&�3�ጅiY�e�hO�����&��<N�����Odcs���v�]���93S�O@)����iF�ٌ^�.��(l��x��W�~���m̅�G���&G_h�Z��B|�7��?x��!���Z=���?�ϧ�@ ��h4�.��n��q�8Z�-=�hq��$$7�@g5"��Z|�j�F �kϿq��-�"nqx�LVZj�-x�Z��<��I�ٲ���'�E���Q����G4��1@�ǉ�Ĝ��ҀL���e:�������҄��͝-d**JO�-���3�q��('���O��{�D4�����gd�n�ܗg_ܕ��3[;�o��7�H������}�����%&i։��N��ĳ�6�!�u�z�h6r�E���F]c4��\Ƚ�W|$����r��!�0�!F��[o�:�`_6�vi�Bp�YZ,8iG�e2��r��K���ߐ�_�O�����ь���1�`&	��}bUֻ�79���G:o00�X��E#�����n�W�x��֧"�D�N��7wv��s�����4��d	^�@죕��b<;���R���wrt��?cZ{�r| {�5�j��*�� ߊ�|"�� ����_�o��b^�~C^�����r�N&̜a�j����N��e�k�_k����j3��&	���6�ǹ[�6ԉ6q�ƿA�����F�c��zl*��]�,!��2[N6E�Bli�Kn��u������#�h���8%D���H���"�0]�O�ݱPD5�5�@R��hۚJٿ:�d��G�zsm�5��'����v���	�����H��ε$"�	����~B ��i�noK��������ג�I���մ�^�W��}z��3�L�|�qZC�b2X	�OD�3�2�RjC�!�������tF�
\��tF�]� L`�[ߒ[�_b����l)5�X|'��$��6ە�7�w�!�z��|�o�����L(Ъ����A!&���f3�p.Z:��C3u��SOVi!fIxO��> ?�;��{?�_��Az���^�&�~�u�������>譛7d{�fڌIa�b�x�2>�x�[�b����4p���k��P��b<ţ��>}�1�����(��	���B���d+��g��'IP4ɚE�&��;��쨸>��,��Jֆr�(��YGuc_Ԍu��$'�*˘�K��ٽ�]8�`��p�@���{�����Bz���g3�)����(�K�θ\ԓh͝�ٙl(���NXоi4u,0'ժ/�lH�2���9�:0#/cK_�k�E�^m �7m�L"9I�E�D>�/��l%s��K�Zlh�A2?��y��\�u�,e��,))w�o���^Z����|U���MZ�pz��
����9Ψ��ə$�b�V�x)Sz��k�H��M����@ �$B�n�`y�ܱg���ɿQ�u/m60��ߵ��� rr��;ț９|��i1+#*��C�w;�
�XX��"zD��t��@�)�$Ǧ�-PF��D�t}}B٥��@m	��g���H�=�~����j����P;A�{��MR��6�ƄZcݑ�ƴ2��}�B�;���u�n��)ފ���%W��ٱ��'(����'Z�[G���w������&A���?NK��͛�Yvd���'����iZ�#���;��g�8&D
���E�X*�ʸ�<=F�R8�1++B��}/.d	F�0�{i����E�N?2��or�ԹX�X�٘�6C��R���.�s���j���cZi��q���.4"�"��hѲ6�
�l�wt{��%��� N�u�d}L��/ܓ�O��,Y$���=y��>��>@�c�.s��%"��$��	6[W�
�C`pڪ�AęQ�d���V��꟱�0�&X(@چN;��Y���5Q�|�4FX����w�Ҽw�AZ�ω�}���K�~��.�I �t�<�?�_&��G��Q�f��`���@�|���IV�IZР,�0-���ꒄF�H��y0׵3ف���XΫ�$+nB��\�}�i�hOh�n���0��TK��ϵ�J�7��0�g��=	r5�r�~�mV4M��L�E2e��m
��ʜ�Q�C������`��3O�>�����/ɷ��rp�@�6����PM���=�O>���*�i������7nȵ�����ؐ��|)Y�Q����W��d��Ut��ע���r6!�g	��xbC�8X������?\�����[���v�#H(	�<Vv�3���]� �{}t]�>�]��`������M5	��v�Wa,��)�0m��ר�����v���Dp����?�9�{�q���d���t1�b�������%���d8^����D"�# M���@����is>�/�~F�����ƍ+t�<8��+ZLM�>��F���¥�>ԦT ���q-���r����*`1���X�� ��@���YQpK�I����w�ӻ����&+�e��������v�_W+0L9<�g�?ON�����m�	}Qhfi]��/��B���yZ#�$ Gr�ۄ������%��"�Bc%,qVK�J��W�NqF��rڀ`�{P��E�Y��9PP�%�vp#Z�p�A=���^h��?��?�7��M���a�%kn,IPǴ���1�B�`����@�f-=�����K�N�}����T��׷���˒����fu���l�X��4�~��E��OLÀi�#C�%��Y���E�k��-����Fv^U��?o� �6P &���'OX�8��s�7�|T�m3M�y��A=3�a !�1��G~�^C�2��akJ��l�h���H���]�;�JXo�ʿ�o��l_�����p���ޑq���d������Ri= q����E�^����ޖ?>|����k����iwD�6k묦a����uƢ`p���.�Ty宏Gg��Q���Pu�|�(Wn^�?��{��G_�����"�	4w�y��`��-Xf��e�Ɉ���#���[o��_��S�4�w���ҀbU�{jY�US������ĂŠ�(�n.IH��lu,o}�U����K;�BjFNA��Z
g
��'���֐l�'P�ӓ9[z<x~�ε!�fA�2cUn�s�/Zl��4*+w�Z�;�2}��Vl\v���L�{����hMn�p�[��Q @\uOpw�Y� E=d�����h�m�� �ɒf	�޸�����S9H�݂�N�
�~ӕY ��t��T���Le8��<��T��Jbw��ٓ���H���.�r-�������N��.�
����	-���%��s�ڵ@�>�?D�=��r'X�?TY�-:D�Tz1���bDX#�7��	�_2�����J���e}̝�ސ�_}���Y �	�����4��6���@��Rg4�a�OȌVW:y(�{�t�u(��8ʺ�}-j�,����p:�NC����q(���>9$Q�,�Np��p��0�)U�h��}.���w����Iq��V)��	"�.�]�n�ul���I�'�š�@[�Pp
#*K���';��'��?���#���0���E㦬�A�SB��q*��~����_|����T������C�O�i���M�W��^CUY3ॡFG#m?��?9V���;���M���w�O���"�1W�U��t��:#bNJg�Y��Ĝ=c�1*���=����8-�	) �\�7�ܐ-\�4��xM�N��A�Hz�� �̤&I�m�U��<F�q����\.T\C�;����-����B�^PѠAB�S皰�2C�fw��qQ-~$���7��m��d?n�Ty�5����am�]qwѿ��f�~�,�[��мƞ�9��z(��h�ю$t5I����ieg�8֞D���-��j&#���J�n.�=9���+���������;i�F%�� ����ot�-�,�R��>���H�xz�ޚ�ڸ=���,�FQܤ[�G���_|��H-k(P����+܁l("�Ч��J� 3�س��4�R��_}$���w���������f�ju���P�����]d��X��G��/�.��(��
��%�G�.�h��"��/�_����w��Ӥ�L����C�=:���X�V�ٚI�3��/�����;�����Ҵ%�+� �'oGh�yC��j31����a�4�5��?��}=Mr?��~�)��f��u\��,8S)��;H����3�ݑGI������?�h�BF#8�����{��<��3���A0B�M��8M���;���G�9�}vG��&���8� M���t��}_�;`&,#2w��UeB���ov�*Hأ� Kr�B`���co1fe�'�ң��H�)Sm�1a�{1X�"-�y�e,�*d�L���y=Zj�=��G�ɳ��|~�_ɭ+;�[�66��x/�����rrX�)�!D����=�cT�v��@�'�+G�3
B ����<�����rp��ݐEM�w��f�yQm��g�Z�N��e�b,>��S�˿�w��*�āb$3�:�Y�z�wK���%A�X5��h��xsc-=�!3 ��[C��������|q�|��C9������9gɝ�J�b%�:-�Y�P@c�:Y9��䞂�Z#_IΔ'q��e����>���7Q0�n�	���O�M97�S0�!��4f���l8#]��YA��Yw;q�S%�����d�|���i�����҅���Ek-~
뜭:�3O��z�\fi.�~�Y**��X,&,j�#��8On� �/�"?wn��5���	��+�b$Wu� �}Ԙ`Vqc��!��W��A��k��^=<[��[�K4�~M�D�����KJHK�$ª� �D�p]�u'?����d��O���V��	�X����)Jy�/z҂� mAhsmgC�$���<�;9Y�V�al�:G���w��&i|0�7V'����Ȁ>EK\��.^�C�
>H�������w��.5N�1'�w�,�I�(о�ɚ��Y<&Fk���-Ԭ�D?^�@޿��s�Cݨ�p�Phup�"�����-Բ�΍���X_l��� D����ׄ�����2�'�\��P.W-��iCW��e�vd�G@����60H�e��qRD��Z�L�u���k�x���8�&�����q���әb\��d8I�c��Б<{z �W���.�ɺ@*˗�(*��ް�?z��DE�����"iY�#*,��z��t���~J~��9�Y��/O��,�����J<���V0��W��8�����ښp��r�^�wNҬqb�O Z�F������\�Y2)QG��};�Mu4Ofs�|k�;���%'Y_`# {�f����'� ϒVK? nH��0?��`������&i�LC
#ϸG�%�5��ik�w��4��G�����(-�}y���i��:��#pzV�	���@��2$p�������!�v�̆Ԍ-yMr���+Ě�ȇ��Z��]� ��U��d���n-X��z���n�I$�C��	æ���QZ�Sg�k*-D�Vc)~�oă�ѐ���Z$��,|�5H7\�6�ev%mx�;<ͥ[ī=EJ��ح.j�&����g�D���7�s"��4�Y<("E�e����Ҽ��A3�֜���� :��{�j�z0܅����MΝA׃'%~7Eݧ����R�rS2�|���m����E&��O��  (��0o�ֺ �'�j��G�7XY��4�V`��i�A>><�u�����$��Gl���(�{�&Y,SGN}��Gd��L���H�A���=����M>-�#�]Ѭ:x��F�.J��ec�l}=k�P�F��u9�ٌ�}^�tacB #
"T��������!d���.�G����>�-�_�}D[�56��E�
nJ��dۺx�L����n�f�G��]�T�7[I�9.&ĪJ��,�k���z,U��4���l_FM	AC7�J�a#m���*���3����E�:�)זJd��>0�%���U�n���V1>xv�� 4�il��:!�h���,���)O풬b��:@ac͡.����r�X-��L��;8|���d�d�+�gB<�c�A��$�'z�Z����p���6���i��@�)�2AԿ�ų?άnک��V�4�B���:��j	�m�XS�E���Z4�'c�, �0�AQGsHХ9q���c��z˹ç�hj�1쎥d��� x�h�P���������;-@�7�Z+C�F-b!��7��L�#g� Q"�ӵL��1]5 ��Pt�Ԇ�N�p(��«{K*�#���4Q�HqI> 7��!#S���7n��A[Z���d,l��(8E���a�qi�#�Ӗ
� �F�[S�F�dT���n8X*��-��n2�(a�@n*1�|����n�XX�z�D�`Ӄ5�����kT� [��W��h2T��]�O:�ks�����p*��*E��X��������"?p�ndS���h��	�'!>��^��; Y�����Kb\�A���v�){��,3v
���F���Hr#m]�H?�mk��$�0Z]�t�3}*5aBR��j�S#��[Q�<m\ڦo5]�`tf�h/Q�9P�$�A�ըB�~<-��M���ͼ���ʴIg�(4,Q� A���%�5b�o�̕h9,�� s>���a(l�AK�[��qait�No i�x�����j��{a��Rv�X��c���{�,9^,�K�$� ڮ��1|D�>0r�;�6�ƍ^F`kg��5x�C��Q�G��\Y�d��
�P�U4>CW��jX��?��U�����BH�/��P舵�l���T�0� �o
��FW�l��{ms{�2~%jYW�fT���X�s�,@��\d�L�P�eyT�O�����
���a�T�_�Y"���LFo��A�����ȩ�Z9�Iwq��ML�)���-�HnRg�V+�'�VDp*h)�&�K��\DM�ڍ�,����5FEP�n
� z�e�x�&y�tuo���bN�h�F%��P/
s>�L^d�B�u�8��,���D��ٲD����'ax��i��iX;ΜO�DI��y��:�ZAq�7�C�>3gQ�����f1��)�%I�=��ړ,�-:D 1`lXp3�*,z �%؊Vk��/>��B��kC�ө��>�n#�ՆM�Q#��aM<m�yBQg��L��k��uN����_ݕQl���7�7g�.:�͌�2���]�X}�	�ڂ���q���Qc���0���L����~����F���ؘТqpo�AM�i����g�]��R�#��U��Z7y�[xj�`��hB�;J{ذ��B���:D�Ќ���9��".�u]X$�K��H�k���cF��rU?��$6��p	����4N�i`�q���J��F]͊e�Q���Si�ݻ��Ѳ~x���w�d6^��eaM�KU�XlXƈ���v�F��~B�"�	K���I��
	Z6� ��c���G!Jq��Y���z�'<|���Z�ε�!I:Z Al�슲��x� ;�!����Yxt6&�h
�����e��+�Gs��� ���U@\c��[ö�U��$�K������ʘe���rY�8i�7�|S>z<���=R�]���|����t�Kq���¡��|Ն�̝��Xl��u�\Hl�^'�E4�u�ZW�5qm徽Mhv3ĴcP��?z/��ͮ+j�(
	��QT��s�@o�$D(<��5��":�ut�6~&G�%Xe��3 �����i�F9�UgD���gf)�gC?���*��.Wخx�ȗ0�G�Z�G-�S�H�zA��ƱHBE�Ѳ�Yt�<��w�=�z�s@WD+�ҕ�7���iP�X�uEV��P�!yi��<���^��|����ƀ�ސ���O�����oΕ����Y�a�^y���e��d�g ��T�^e!rz��P���i���_�<�:�p)g����c��qτX���>�5-��^�� �+�_�ǅ_��[E��`���G�2(F2^�`f��,�lN��oe��`�j	���E���"�D4���?�*�2&�$������C .X4���t���\����B���A�wZy�����.�sh����%R�C��!"b�-�r���H�YXh^���5���.��XҚ��Q4X�FX���������{�ߤ}�!�\Ro�����+�.v2c��it�ʀ�V!�M�{�|��Z��`�G�+6���A|4��Z��jj���%�T��,Q� @��ǭ�&��S  ��IDATU��:�j�]�K�?�C�Qh7�qɱ�O��b$_��4~��<z�(oh�x74y.���W��+�eǹ���--I���#k����E���Y̦0) ��0�y�n��	��G=w�B�D�e�G� Mi�Z6q����L�*�J3$�7���M���8=��N��
 Sq�.ph�9�I�-5P�Z�Z�QH��'�f$'@Y-w�����5�3�E!ԅ<���^boU�-��bL�cAC���sk��:�׀Oŉ�m���	���� �E�9�s����ig�����`�$Y�dJ���:Y�����R[��|�����:%�;=?��ώ����������#���u/W����JܢRN����?rBDS���׼֍�lP���Z`U���b�!y�2�?��'�}&��<�0ZϚ�����u���ć짪0�*�`�����_B�9��4Y�+��8J�֙�ͿVK"h
Z��Y\��l:G�>�HQT���U���M�zo���ؐ�����:�qt����Zn��-���d&'?�I�����P�d���Ɇl�^'�E@N���U�٬��8}�rI	,93�,���]jR�8bq��	`��/��
���n���;��x�'l��)�Nǜ��V��Kt��J�*��-+����W��Q��
M�Z� .�����55��M�h;Z�v��8�g@x<���ũWwv�FI�[c>]�1�j���*��QYh5�4��v�]��� ���ޛЕK�r����%�S�n��z� s��ﹰD��]O��Hf��|ʠ�̀A��<j����wKM�h�J�n|F�$�¤D���s�Lޕ�"�Y码׎��5 ���,	����%�����LK��H[Gӗ�Nt�5^j��Z�k�0N�?R���Z���
�k�/1-�#�k"'�%EJM�k���d5,��1��6��O�`Z�HX����]Pn�'q��+ƴ��;ƭ֌����i����5��Q� �M�P\a�7ufqw����8�bL�����D�kU᱔�g�`6���3�L\]d��p������W�q+W�oL�"͕��5-A5��h�C�us���h�^-������S���j�Cq
D�����I��!�ݫ�)]�� 0��i��k�:����K��e� �\��5��$
�,���O���BX�
��X0�5xE�����
V��$�FB��j`5���E�6yX����D��X��%p�EGq���)�=\:����g�w�ͱ�A,8�k�6C�WO�J����.�/)�ٛ���'�,\S��)�x�f���t:�6�͐ܲ�8d�$��X��QI���հL�6�7�6�+В�R�t���}Coj���~Nک��fĺ�E'��0�c&ˢ�i�Co�v��������x8�V�K+��q�����q�̜Y�}�^Ǜ��?�����t7ʭ�΅PO܃�� I��ёL��
ņu��S���t4��j�E�Y�oAj͂�b�x)]�8�P!X`㪖�HJo�C��B*�Rp�����ۙ/r�J<��O�ߔ��1�R����O�b�?XD���s��GJu��#�����n�I �j�sK7e,��S΁=�I�`���o���K#�`�ݙ�q0h`�@h��|������=�*�r�t���X�D��ɍ����X�53�iR���B/Ht \Q)�@t���;��aL��Ex\����<j�/��<|�������9��SY%��Mv3zs�Arj��wU��������碍W�����w��&ls9}�{��}g��@AXu�����tFX��/�3�G�E��:.��n�\��j|�2w��v�2�= )�������B�NB9�h�%� +{� :�єF��H)-�=���h���]������ e�IV$�i ��'�ُ}�~�Ǹ*��HI>��a+�Y���s4����q���%�$��w����ם=3���-��H�4��1R��$�mֆ4����d� �u���ߊ��`�ȧC���%c-=��0����hT��!V�z��`���߇�}n���󿁦��8u�$C��4Ɉ����~˥m�oK���B�����h�(f�Y1�k��L�M�8�Ј�8��fr��[Ϯ�����nh�xh0ot�f:�D��Oɺ��� �i4�E��
tҹ�"Q� n�S��P��K͑�]����ɺO{E��H���<�jgm$} Ƃ�L��>,���>�/2�NI��y�v��Z�4�,�;�R�%?}ii��ʃ�Zz�J9�����y�����τ�k����|���Ih�֨���0�6�ZEZk����Ђ6�O���&|Y3Uՙ;d��-�%�
��Q�HX��:�^w�a?tѪEQZw�<)�׺�cLh�T�p���R�b��?�9�=��NY��&�%6�M�k���agԿ��:F����n��`�%E6}$���esޑƀn`�i�Q9�q�:��|QE�����4C+ú��Q]Xڋ]a�(� |�V��]-G!J>G^e��*Q��H�.��9*!+K	hF�̨ت`ʠb��.���E��j郕��������1J��!���s�j��:��֒����<����T_X$�/1�m�7umxE��bId�o��m���k���T�`3A;�᐀
+pP^�ۆn���PBo��%u}uF�и��;`�E\�ڂ)ݒs�+�|q���G��V�\����&�p�N�υ{����U���.AQ9{a� .Ȁ;B�Р�ZS�EK֫[1_**��&� >N:7ji�N��V�p]����x�>h|����P�璍�Q���6�Y��YUZ�f0�ScvQi��!,��B!����G1!��ރ��V?\�I��a>R,&<������;��(��uV ���KLC]�i������~g�Z�?sv@��JW�tG���3�tcV��6޾�rc�v���B�F�Q�,�8��(8��qe"�U��Y!��z�.f���Z���j�d,��7ʹ����q��2rj}���@k��"�l��R8�������Ӗ�Q���꼔�`�L�Y��*�o6��=�g�zn��T�i�"x90��,z����$\P�'��~f�X����P /n��h�h���{��o#���){I/���	�`��\��،�%|	�s�s�����;w��|��ʴ8]�BYe�w���-C�CE?�*����	c�@�M�k����:�wڢ���, -�����r��**��QN�kyh��>!�S���em��K��b�!��p���5{/*wF�T7�8��5t�S��N��I�Ѳ���֞3�h��\�ªf6Ԯ	VR�y�v���uc���P�1H.T>�X\`��2��m�W�_.�L�d��π�F��-�mqN�a?*�8;o��� ��4�����!��d�mo�ຆ�e�JAr�5�p2!������k��Q��ҍ%*��A4�,�ް�6n�������D
���f�z��tnl�i�ؐ�O�� ��	����s�1��7Q�D�/	���(a��A������e��5�>��1�T;��1O?�1�2P�Oy�
��v��O(��z8��~^]ڒ_u�V��%I��LiO����w�GA�*6`V ~Y@��.ϕ� �@�d�q���-ϋǱ����E�������S��[?�}�P��$���v߄ޘ�J!�{����~p�h�cA���>����DK�QڄD� x_S�A[>tJ�>����E��e�� H X|Q'#���V�>��{��4k�Z���͑ݙh�H�u!B8�iXҘ��/��/s�nB��䡪.�M��n��Ϧ��d"��\5��㼳0`���X|Ƅ���T�q:jwi�!b��TN�����=��Dnfٝ{U����ք�Z��]޸�ų�.�{g@1">�9}_��g��7��F���H�D�?fW2���O�B�?�?w���J�\��+	��b^i��V�N�_��n�)�ME^�Q"MrcZs��/�Au��)M�����S��m�VS��B⤠��������*����h.z��V�����˃�Μ?/P��3�W{ _|x�ɵ��*T��A%s�J���9JMt�i<O)g�X �f��V��K�4E���pwfp
��<��}��)H�U��0UY�
���Ī���Q�������.]�q+B����^�ٞ��
���X��\���ߞ3�;^6�&xO�H��qs�9x]��$�J�T,0?k�������p��|�EWx�(, ]�;�=���J*��)�/N�s�~H�G����'���"PLQ�[����c����P��˚��,�3�+�Ƣ�ͅ?�/�l���j(S��9���"��5}L?4;o�3Q�����s�V#�U�k{<KT3�	<�\��%I�..�[�����k��/�����譒�~�y�S]�	/۔t.ދ�W^QΟ�'����x��\�^���/�sԵ	�,(���e]ED*�9����ԃαU^h0���6d�)����+�ᾭ�
`�h-�:5P,��NA5,�DM׌�������T�v�����5C��E`U�Ȓ$��͋Q���w�zG�����my��?F��}d���</7J�S��k�S.�;�!�L��r?Y�PP����ɡ��Ore1\cZ�ܞ�+K��L�!�	�d�Ų���Ȳ�㫂H�	��2��\.���9g�.�ѷ�y��������G� ���%��=�M%dE� W%�s�v�_l1ڹ��H_�Mk���R@?#��m�m��neb��Җ�3>���8H�8�j��Ap�`�� �	�h��k�X�hdS�O�nݝ�^<�����1��S9/��0G�=� =v������yy*�3�fc��2�!V��7t�	, i�$�����\�?(牣#s�^l�e�S:ت%3Þ�Ssn���)p��VGc�U��ܔ-��:i�	M���@���X�V�H�`��}�.7Z�����ĹNV�����xJ������\9k&��\h&�N�Ez%�)��8���6C��Kp��Y,�NZ���'n�d�c��D�{�P����4'k�^��gU���U��K���q�>�i�����C%��,د�+��3@��t��	-�8;��[�\��F�&�A(HE�c��%��&�@ɞZ�JWڷ�̫$�
�J?6RB�m�W�s:�m���~�
�h &�Qkl];8H]�ac@zzJw�m.ъ}�h?�����m�}��2s3(WH�*^D��# �n[C�EV��X�Ҳn�Y#�@�5#����\삕�?�l써E�y�Ue�RT0 ��bJ�O���=d�q�LNh��C	�V�J9�����ʷr�y�_m(��jy)�5#��^m��惿
+��\D�ꖅ�3��H�v�]t�V�*���WM�����&]Y�c�bn�����/\(.me�eB)C�}ܖ鞆C�ȭu?D����|ƃ��u��Z3�i�k�ԭf3����lrH�N	�$�,>�h�����0��	�����bQ�W	��qM�� �Y��-ə9�T]�l6z���v��k��E����mBUY!Vg����������iת�=�,-{=���-�ޏ-��p�:_��������S(7�ʐ��SBf�!d&qH\��UR�<���P)r}^��	<��K� ���E�ը�w\6ưdZ��2��P>N���5�o��箷d�9�Y���V3[��F\�ֶ��јc
y\�!N�+Dָ䲐h�b]�d��[�Z�F�˓ci�OH�TW*����]�(�����	�;��K��s�W_���Q+�5�d�ދB�X.��mK����O��B�h`�܎(+�x������|у����(�2���>�KN�AWŢ�M��E��]h���:E9+I�,����	.��}a��k���"3|�V����5o�3R?ǤÄ�VIsJ���(�~��b6�<�?�3����&�%G��N�7���K�=)1])(��%9��b�N���,�BnA�/���oZ�AQ���E:2�T��V�9���.LL�cq�AT��o���"��l��>Ԉ�Ī̵I���o/�@�W�I� ?��{��D�: >�(��1!���L����R�d�4V+M�*CvŦ�Q�d�m�߶0�X6�z���;K��,D�7�n���[��eGY��jά]� ߂�K��BHm1 Q�&R��dWI(�9����ѻ (�@j��,(<&�+\��r&��]Y��p6��x�;+}����9{t]��V����
��f���YW���������Z/]��	C�����'�۪*��$tm�ڀ�X�I:TuJ�������۾&�k8fQ��H�>�����i�-Hy���>�@�o�4kK�f�P�����9�6T2��(���.lJ�X�?������ꋂa��sNq����C�\��7�oA�KD"�����RSy�+�^_�;���̌a�_N]�G�3]�Vo32��º��/��N�7�[+��&��Z�h����U�ϝ9Bi����~3\l���VU�	����E{��D�R��0��
��B��ɊЋ���=h�u{����'d@��ja� ��G"h�^� �J]X��"�"��KT���޺��s5Yk�|��\�����ǥ��>��X���u�T�Zq�,�X�X��`3��Lȥ��/s��K�U�V/"9vR�Z���\�/>�Y�������alh�Z�v:�^���"���9���[12(.� ���<{M�8( Dd�j�ι*��_���p+\��Qy��wZ9n�,�2��z�h�Z�E_�e�����WC�]�vn��ɭ�rs��&�@)Agy�܍����J�2EF'��8\��#�Ҿj�g�̤�4�+���@�G�\���E�X�M2amv��k� M���� ��F�e�^���[�7I�����o]�ݭucۀA��cfc�PS-C'�T�'�z���(�i���%X8�� >a�yN�ά/��؅�������"񲅾���V��;}�+珽ֶ��o�xHj;YY�k�Rߗ�$B��	�m�a��W���#��Ԥ}:��6�d����6Cl.b��6f[�Qd#������j��]��TM�Xz�a��E���;hW�tb~�W�*�3���y����6�e->���g�S#_�,�j�(�}ɞ���dF�b���3c`��49[��遆TH�*���Bq�.�/"ň���{��M�eu�W�9�
�l(��{{ϒ�ڐ���s�C��_jh���k��!�N���1��bZ�����+�8��*D�
��Xd�6�,�Eς�8ț�!�=�g�[i���<Dq7e6�<��K�-�2�fs�+.�gS'�м���;t�K8K���Y$v!���Rr\�ES�Ύ�7���.���kRH��5���؆r��yB��z�.V6�kɂ;��=[��U�k�5W����s�u�7'�t���j�(3zA��'����Z�|��`�&�рY������BLk��OYkT9������C1fzy2���a�=�KY��y ���Is9Hm8�6�R�M<bۉ��:���2I�Ͽg�l/�R>��|Ъ*X� �ƾ�'9N	��;��{5_�"\��҅��۪S7�eЪ9�ou7�%���Z���+��ml���.@(����9��(� �l�[+,�P�ga���˯�㠕�0u��o���5W��B�1���dIx���7�ͫ�lZ��[�N3l�n��d,=����E��q�B8��]+���V���<hA1���^���*��9��Q����;����ވ$����zV���	�i�G��_�0�v�h��'f.�4G �BF&j��ƌmY��D�5����Y�3����������ݯbo�,�N��EP��}g�g�h���dM��N?[}팬�Ϲ�|�2�q��#�ub`4*���.̦�H�����יs�R��d������Yr����;�w�먫�X�7�+6⪮��b��KEk�5Z �w���t| |TZO�Sɡ2�T�UE���[�!�rs���V���9JS�8���Յ�6��DV�DV��)X�|�E�����q��7w�ܾe��*�׋��[s.H�,%�!jY¸�\�����Z,ͲQ��,�E[�����ʍ7~��9 .�쪈ZG�=H���/�ca�=�{<ēA<8<<b�C�N۪%RTZzem]�_"^g�	�&T����mW��.��=V��T-4
�r� ��~�ɚȵm�"�Ԋ<��6��]rɪ&���YX�H�}<E/)�j��4�`�b̴[ҪV�A�1�):@t9e-��\(�Oj:������o�!�G+�3S�+�����1[%x��Q
򢹻	�+���Y!"�!������R�%xW��v�/:{���<VA}��eN�,�KB¢t�f$Y Í�@��i��rGϬd�Q��q��[+�}/]C���>e2fWǪͣbs�@AM�V�iZ<�Nu&;��6�5�E4�K6�+p�Q6I�I�'�{$��Ͱh7Q�p8���],�<X�	����E��t�j��L�����2Y�NX�]�:7�5�r,��vL<�f�����m����S�����4�8�4Т�oz,�|�-c�@��Hy��z�tTLϵ�uA���C�ߩ�W(ϭy��s�.��S�8}�����LzvO\�X����1jXv���x���v��]�����*l�T<�*'-���#����31'�9m�gA���K:��������wt������7�� q�?�["�έ�qox��^y�SD��JN�9U|e,P�ӿTL�H��N����ݼĩ�ӑ�ػ7A��I0>�D����j��E��������@.�B!�V��%"��8;�JxJr�DX��Nx&IBX��5���uX�����e��fQC!�\��B9I��[[��9��]A-Jh�9�{��'�9����8/�ń6j�x��Y��_9�*i��eW�����ܲ��>f���U�m�r��̾䑸pJaa�E�M�iKjik0���Cp�1��i���� 2Ցk����N
�M�cM͈]pS1��1{p �w��)fΖR���BE�*���"9���(ܙ�I�^�xN=	gF[%�Չ`�_(�l%w�V'?�R؅�U��������_��Q0�\w\���̦�r:�
��UB�ОDbd�L,J�����B%��s�i���Oª��K)�~m�k�&e�b�~-�r�F�!�@m�&5�>Oѫ��������%�6K~k���(�=W�K�<ԛ���O�-6��N�����-�9�\��h�J�j����%�N$8�yG��5��/�-U\f����'��ٚ3�p�x7�P���u���y� �AHG���v�%��Sg4�Xc��C[XW]��.���Z����w�|�c�C��]�Lmhщ��&���\I9 d�-ڇ�����2�Ї���4@���n��7�o���7��7�%_�������2_˒>z�jK�����b�j5�E��=x��áJ�)�j�Lym��l�di.X�P����b��7pMHx[3P��[,Od�Tl.���)�4��Y���<о�s.��bD�1��4E���[��;Y�cA ��VfӖ1�V���Bx�`��������*���Y����LcA7AyK6&�:����h����7c���A6�۪��ܦ4k ��� !<��D�ʃ�$Q��x�Uicu����4��$㎽�W$o4�d�:�j���(�q^�@������Z�sk&�W&p��6fW�Xg�A�2v+j���!��x�sA.m,���Ż�g�\^*.:8���?��P��Ҩΰf�B�@�h���܌�IZ�x�f��DkX�݀h�ᨑ�dْ�~���[��}�W
����|C7I�)S�ER� /��N�M��g��d�տ�/xW�	o��7����K�ݰ%�|LZG�u�?�󂟔���7ؾ��2t/�c���Q���,]�(�hI���;�ɩ�^���j�E�o}�!kI��җ����a�]H�bX�"J��R�Ǎ�#Z��[yAo����m[��T��P���j���HWk���v.�t��'ٞ,�h��}�c�B�k��f�s�@,�	`��	�$@4�[L	���
H���2�sQd9ހ�e~�xqp�[#v�-����f��u������;`�v���w[T�F)\kw�]*'\fAh\.��47��@��9���I���y�K5��,GB�Ψ�b�D_˻3 f�[/��%�Jc.��f��#ѽ+� �X�i�"�~�;n����̏J�"�G�W���<1���X�a�3�$s{.�ٕ�}a�1�C
@UY�4��>5��\o�:�RD-4�ULo&�<��z1�0L-ӎ�Ρ��QGR,~mOa����ϋ1Aq\��(힤���#iɂK� e�"���Đ��4	9NR-�d��s�MV�ޏ�Nj�',v�����l]��$�V@:�$����.'�������O�X��PX8M��;�̄ �\[�LNh�,8���ѺF�6�M�[ђ�u�X�d�V��a�7�U��J䪾��TZ���e��X-��X�������\<d�VI�^F���t�*��uW���І��q57�@���F^Q��{6�����[�d��j�eG���2WY�=��b���j޶I�1��5!E@y��x5�yvEk�����Լ�ٹk4栦�vy�B�-��M4�v�jD�㛙Дp���Vb�ڑ���f0�A�T�h �5t���s���@o������iÌ��VX	R��Ҋ�2�H�f5���ϧ���V(�|��6-Y�5�R�ӈ����Kw�`�@N��5�6��tFA�ʝr��U��/)?��Om�F��N茊���ME+	A�7�\�?������.]��O�%Kx�Ͻ��-y�����ǿ���?~!����Щ}���.�ٯ���\�ސ�ͱ<}��\��=�;��F�r��H���i�j͓[���Xc(l��+��:k��;ѧ���iY����L�E��@'���E�T�ō�X�,��H�,ٚ������R���$�����k�6�LX��-Ux�v���ߵ�/�EGy9�g:�',P��h`<(��p�*m*��ʾ̡34w�:��W)���e���݂��L<���|_��мf2�XL!�'��bW	��,X�(��.oT$�7�l0邠���cl�P��\�m�Nf�ښ���ḱ�Vћ��=<i7��ɳdi(Y�Ӵ́�ɤ-��@X0m�F�$9$����� Ҭ�bJ���ۯɟ��?��^}]޽/�>a@����+���m�u�|�;����bz��e�Cy��Lъ����J�~���}S��?����y�衼u�UZ!����!����|�ʦ|������G��Z��}��o7a?D�']������ܹ}]�6���)�cE,�x��Y+��$�窌��<���ВD���Y*[�Fp�3Ŀ�}����k��+s�α����f��79�����,�G�������mi��G0)beE�*�dw�۬���7s����U��2!/~/j�M�,�� )~�["��moM�^ۚ�y��y!�w;*��T#���V�I��f�鵕�,:ˑ��0[ o��d��rnXƲ�Db�Ù�}��\V��U��j�=��*�5`����Ớ �t�����G�(��Ib
������<��[��o3	��� �09w��@�w��M�������Gw�$+`��4��T��aZR֪1o\ߕw�����ٕq;��t�G�'2^����y�k������_�뻛����zN^,�Lh�\��#���X���;��{?�Q��Wn\���Ci�P|��-�A��W�"�����{�8���8fE5�g~H�\� A�|v�'o�v[����粽5���'���sA�t0�Y�m7n�$���C����J�k&���F������?|M�Eex�p��m�q<��;�|�4]e��̈́H�����@+w)B�U� 1��eƅ�X ���J��V�I��Fî1	|C�bC����ɲ�˻���ګW4��q�HQrH1C㱤�����#��ǌc;f�W�b' 4z﮽���n�s2�{_5 ZC��(TWի�����2O�<�v��ԽX3ʾ�p�؊�$n�*�ıE
-_UJ�����܋,ۖ������GZ?tbqsw3�,@w�j��\8]���V��0����L�p|��O����'���]X.i�f�ҍ�2���b{�\�`�α�8���qڀ=���/������忖|����#YL��Q7�����m��Ơ����%���UJݒ���ɃT=z������2o��1�S�{ggC�I=�Si�������P������ f'61t���F70|������T&өl����8��v_���i�Z%�ޏx.��l��e���W�B���7d9?��i*�.����8��������y����;o �~~(����A�$�`@r;E�lT�Ad��Ϯ|���ٍ^�_����zd��l�1c���T��
^ts����XB��2֥{4�k8����<!a�Q��¡�@$������3d����;��풱'B"��H����	��lF�:�A� ְ{m�>���@助�v'��O�9��:낋a3Q���e���+_�FPk8uJQ]�vY��T wȖL�!6�TBj�0_p�\���@O��Y��mI99fvj��q3R��V���^�+��ݖ�zW��-�-5`�����ŷ�O����G?}Op�+��c�Đ:e&פ(s�'u�ׂD�@�j7���'r>��h�{���'A���,�`5Uf�U<k��%+?7*-=�K�a[=�W_M>x�I`��#�����x�9}���j�����X
�$P���hA�Q��}��{����D�9�x����������� u�����1���r��P�6z�E���;.�֏U8������h���WE�!|	��������� FR�J�n��]�֩Bz����ֻg���ƙ��ũ��3�� i�3�U�����rq���<��[�F�ڳj�ƀ:��`�5B@�	�0������z� ��� W��$z�N�,�Է�TpĽ�Ҋһ�m�o]zìH1<�e���K�{��\���s^Ü�s�^\3�@#y@L��,��V���4q��Jl��1���g+Zm��0`�o��۾� !��L p���n�1�A���C�256l� ӡv{kK���893f�nԶ��b.7n�R�aK�����D�7�am���xnx�M�ꚾ$�PlW�¬���Pd0`�UY:|���^+с��Z��=�cC	;�U0O�.���~�}M0���C��o�X�շgDoϚZ����U�vP��V�%��D��K]�`)��@b1]�W��B[�&,�6߁�㵗<�z;7]�܀�zX����x|�%X�/��W�BbUӰu��<�BA�n$�e��B1���H�y�Lꂍ�5�5�Ԟ����dLC"�0����38;,/&m��ϣ��ۉh؈^P]�ٹz_���H��$?��)�U|M�1�`�����n��p)���K2�UB�6��i	�m�v�3*x�6����7���T|Kܳ�ڃ��V9���>�c�*l0g��B�w�"R7 ��ũG�O�5��,��崭h�.��JTz9.����qk��!�A�e�i+@��%�0�������==��|��}O?���s�ۿB�m>��J��-�F���Xy�d'@�BߟTf��V���7nJK7!��:Ls��So�Ÿ�\M��aA�Y���Ռ�j��"���'�AWC�)��,�v�F|�!��tB� R�\cJ*��`n
/�C���cZ�ím��1�s���ֈ�� �OO�w�+��p�R2�kl�<op�5�g]�l}c��r_U�]�З����lT_m`|�����RY(��Ts^f ����ɖs]ӥ�� ����腰��B���d�J�9竹�.�%=Ӄ�.��=T�0'�`&�~�M�R�-���5��8�OCv)`^�T)��B��D�+�-]�%�ӻh�x~�{l���l*� �WY��]<1�CR����ĕ�H$C\ofM�A��y�S` }��f,H/�.�6���b�P����)so�:�3�gf��	�MK��3�9ˌ� ��x��魓wxx@0rck�d��n�v�/K��o��Ύz<�L'\��r�F���A`�w��A�\L	���t�1`2wvwh@�n��g�8d$�=5�̅Q�r�3J����I���k�5O��A}�l<>���C[ȕ�o�Ӊ� LcƻpU7F��e��5^�d��K#qz<�s��j4q��^G���ct>��חr���t�b�ᕠ2����>�(�³�+~�5�ʏ諭O��W�eu���%��t�H��!��<����\�c5��'�A�B:�錯VF�,�[Ww���kC677����eBSo��o��)��ڵk���^kSǿ��;����3�����(�C��߆�\�'�~���"?����Ϗ�|�0`�5cq脾G�]g8��]�a�ڤ|�}�'6�@]p�b��֤4��"m�Cb���Մ�z��#F
�$�\�UT���S��^d�66?O�li� .!�*}�X���#���yɢ.�Q�ׯ
Z�(:�py|��{����@^y�%���eS��N ��N,1���f�鍾���jc��#IX��y$�51��*��@7ۖ����{,�*ɤM_�$B��K��Ȟ8N���}�v����қ�e0�(O���1�I�B0S�<����ϑ5�IB�q�sqt~!�㩾�56��v�$SO��А�؍>�o~M^x�ey��'j�ے0/7S�UE�$	��3�a�Ț����6�'���lߗ^,	�ma��K��;}���_�/^�wvpp���=�^�y���`�a�DC���ǻ����9�Z�� ^�X���b���kF_f3H)����!LO����1�IS�{�^qMez�]y��֍k�w?|_���!����n��afd�?�մV9�����=������d�XW�f�P�Q�q_x�:�����6�.Wn;w�ƃ�S�e�7�H7�&���,�jV��r'�� ������e�*zj���2�x��✧fG7B%�F�wv��2X�����K�L�юY��z:��Wa}ud:i�Ǻ�V7�ti���T#rH���&= ��
�/��$�~;�.6P�A�:'�cY�ԃ�w���u9x|Lp�J��b��m�Xmz�N��J,��	v6����9�Þlo�d|2����n���T��75��ס^*Q[z�-+��q���"�y#k{~�T����4$�)������Zjh�ߥ�.dɡv5:������������ -���%bG�Ox ��~1:s4��k�������f}RL�o`�v��}���w׮��`��D�`�G� ��HB!�y�pG����=�L�n����$<���F#�η���wO���<9���ˉ���}o��.] `��� �$�nEJ9��
����9nR�V�GQm`b�k����?�2P���v+��-�|��]�����p���nb�,�*�`��� �4T�b���v��⑸UP���瞗7^�!��'^Fwq!O�d0\�+��&���C===y"g�gruGv��dyZꂘ�a,L�M��t.'G'2ׯ��Qtx'<Q�usW�%��^�B�#B'lT��!y�x�8���OEט<x�X��L6Gb7��{4x�nϼ�����s�"O�G�">���� �L��gཐ������ÍM���Bc?�A���{j�g�yE��R�"~f��4nҊ|//NG8dj_8����
�/�ݳ^��￺�����p��e�F$?b����V,F{����?���Z�O���+����G���7��^�!C�̻ہ{3Yh�no֊a8�������4��B�Z�*�pV�x�q������N$�YfZ).҅�{����zS�� @��� [�z��d����[r���ޟ����V��xق�0��ù�G<,��}8Oİ�N���\8����	��L�������|iEs�)���4�W���z_�VD�w��"�$���1
��r����g ���Ȓ-�ӧ�*Hق�}�`OSs�:�D���������H7��;��+[�]�{�<~�Tz��|�e\�����\�R����E�vGr�aB�.?6�|�$?�R���.w"�v_�x�U��?>�d������=����L.��7�%��Y�����T<�r2l�-��^�gÞʆ���<�Mzv$[W�j�d�˃�cI{W�:�EvDھ���t��l��}��.������<}r$�ի�ɽ���~!;�����t���u���S5��=�~�'��u/��9����-���n(,��s}����_o�}�i��q���4��ʄ�+������.�0ʢR�)T��0����	tPo�t�~����5��zb�F��4��Չ����X��Z�d�Ȉ����jN�����sޣ�������������{����]S35 ���ƀ�r����?����� �C/�뵏�X��l��FG�]]�s5R�.ψ&`q�P����?c��;��_�p����ŀ�ZO�r~�%f�sl��y(k.�@y����Y<T�d0��&%�냲��t# �!,���1��I�[]
�±r�m�愊��(*h�B�m.hI�EA�h�.V�{�t�n�+ן��a[�u3��λ��@���+;~ ����!O�.ZSj��#{�81���Ñ�̵�
��<<8���'r��_�A�T~����s/���,=�;w�˽�����^E����Ăᔅ]�$��zzݶz
'��;o���~�O���8!r��Ky����D|���c��i�$���H� ,�v\��CTxrq!�ݓ��{O�;o�-��ױ9�_���v��|�/�\��0�3�>sJ�2�d,�Z$"�/�Uh}�e��ӱ
�T~��=
 ���5f����bT��ȍIZY5o�8y��"�|"��Ɇ���������o���HG�j�fӵ�B6P���ɗ3���G�	x��.u���P���K���&�h���lt6��LF\��ZVj\6�"aP$��+� n8hm������W�m�ޟ����h5d��"y8�=�0x��q�xc�PHvVO����	�P�u���R5v�Z�<��T�kЈ�e:9C����6���]�V�CkY��'�OȀ4u8B���?E�l��	̫G���/A	G������w�.������'�h|��B'fB�U�t�<|����_x^G��H	`uA����5B�>�������ge����P.�{989& ����FK�йn<�Ɔ;�	��� 	&���� ��Y���c���wd� �����w��n�\L�r��=������#(=��t5�����sltn�2GȰܽ��̦�)�dz1���'d�=y$?��� ����ʄ�0���ܞs����K��]+i|�/Yg��N�/�X�u�y��T5h�|��(HT�֍J;$+2q*:���BsTŢ�����S���侎Ǣ�'�����<@�Zq��֬�hU����5�23TF�=������E"��c�_�a�	��}$���.�V5�%�f�XE:j�pm5���^t������^�=0G 6*+W��W4G�5s��W��y�`5�H0Q �*3#t�E�j�(,��c���TL#�Ԥ��j�@9��3wW{B
"-ެ�i%j�-tI��������e����9�D��L�^�~Gc�U��l C��X�� C���~b���Sr7N�&�vv���\������c� �����jDl�M=�˦��{j�P���x6|;�k��n�8�Q���C^���	Z����'�� ����H;�'����ڕ�4.������?����~�u��8t����Ɲ�x�Mf��mC��]HN�������/_��W���w��]���1XN��'��r�;Wec��l�z��VoI�V5��1�!��������x� ����ɚyF��=����j�L��d?I�t�H�5�T����|J� ����2dnx������@*^ ��n~՚g�q/tZ����i�H;�D6>8P�)1��2�bz�5�v2	�y6sO�d�hscC^{�5��/e�{���BAK$8�P�
LE�>6R���\ϗ
�����u�=�	��`ղ���{��oX��Q����H9��(�E((I�ER���e��>��C>�V1$��Ay�K�q�,�%�6G�������O
u�Oe0�ˆn@@m��ݝ-��K���\'�?�ご���F�e��yXl$�1�H�Х�"O���H���ߗ�����!=}go��x�}zGo�-W��`�g�&FE��%<I~=���{ �����^��sE����}5S5\��ssPԗ��HLV`�H�=8��0{R�V�0E�q=>:�Q���p��ck�y���ń��.֥z'[��#�=Rci�rAk��ځJ?��6&� ����F�2��B���]�k���`1�ة	��2�:YW$��ꜙ��`���5"U�i�c�)V|�j��_�\И,)�����E�	
F&��o�ހ����ْ�C6�=��cS o��<S��!Sc�{���^{��}���H�4 �e�5�B^��+kV�}H�5�"���Q6cf����Sj	}�
�)���D���W^2]��o,��$�IRO:,^�<#��k6�.	��p
�Q06kI���Θ��� ���ƈO��v;��ݐ7�x�v՝�Tc2U�)^uO�Nd�����:��4t�,�a�T�;��c�A'�	��_~I^x����׮r|��{��G����G���k0��LN)� Z�^|��z�)
�tL�~�����%����ǧ�SeD����S����:'�y+7��zc3��V;%���B��7�&���0�3�ں��F�9m�F��O>���[���mdS�٧ GɅo��0���X�`S�䊅�q
�����3�-�b5Y�yaMֵ�Q���lb?���1�9�+݈q�ύO��``j(W�q݂Hɲ|�dH�C ��揈T�x{7�J\+$�=_4,_�	zqa	Ub�P�K:��&"Y4��6�W�k�s�]�Rў-�F�4U�9A_�H`DX�7���0,f{F�?�!A��ȝ�U58\�@��@�I�F ���T!�]Q�$�(N��ĥ����IУ�W��ļ��K��҇<U���1}��a�솾�݄��7e{�/�j�)��рt��UƓ���oi�dUnG7�2_��a(0�iD 6a��Jӂ�py�1�67��8x�T_?fQ�s�n�7��m5Vr����'���� �\e��[��`�"O��Ԩ$����ݝ}y���hl�R���6�ko�)��r��#��X�p44�Z^KCx{Sc0j�!K�o~g's�g^�y��(Nʾz/���\���<��A����Tv��2T/��+xq~,�����tt9�"�����Vq��>���~7Lm.�ኄB�hC�ڀ{s�~ŪV(��V�z��#�i�VA�)0�>Y�2�������a�B�=1J�y�X7x�"�-�J�֥�5@�϶��,\�
z�5�(�Dh�����P,]H:D�]Ы@�hK�����_W�V�AzɉV���i7Yn(C�>�5�h!:4#��K��&
��䐴���٬.��0�9��*�c�&k,��T��4L&
�b V�����%,��+Q���h�Ό��~'6� ��d[fe)Č��!�\�\O�a��� be�����5z�VxcsC.N�ը���� ����m�t!���Y�a`T'����;���@�h>Yrm�t2���P�_�1��������ƐyL��U�����fC}-�2�ax
B@��� 7eK�5���ʮ�7����L[]o4�aᑬ�!~N�J�1s�'^��dk�
��50j8�狙�Ȯ�4Qړ�!���Pi��/�d���"��b���[_�B��t�٩���_m�����{՞�MV�Z
����ic�KCtS�#�����}���8���<]�V����u2v��8�C\P�}z&]��'3�t��v"�\[�ѱE�mk�̤����k��i�u���t1���sl�v����cѹ]�i�����:&�S�����52Tٷ{�O�zo��yǺ�H2�S2]9F��9�L�s���3�І��=���]s�n�������4>�ō<d#�x������XZ���WIl�����EN��̋�2hЏ���+��h�i�PE�&�[��r��ТB��O[7,$#ә|���V%/�pS7Ր�N���G�)C,��l!�Ʉ,V�����I��/�Z��J7J����L��P@�ܟƩ �D��jD���3�����x����[@�$6�l���U�]F�����G���D>�}[����������d��yt|��Z���Ic�01����9S�X$�^	F�p" p��`D]�{��ӰkD\�q�&/���)P����+�k��(���W$�������	��*U^v��Q�{VYN/1!���K����Se�����%Hi����F�XY����~�%u�GjD�Qkr}K�ݓ�O��'8X�ˋc��J�񵗌ގ�^yN�zy���<�͛Wc� `ɋ��{��s�I[>|�T�H�ѵ���	��tL�kJ9;=�Ou-UkD�2 �^ K������)��-��z�
�ϒJ-���rD�1��P	�5O%	)�M���$$e+WY�T"���
�3�x�jqARcHЊ���*zC_UV���Cz��[}u+�Vr��~&�G�򴛒S���d� ��1��R=u�/�rqv!�;{����+��c`���kh{d���0&���!:)jU)S��XÌ�^kK�k�2=��<�ANn��CKb��������H��B7���!��!]�T��P�+�+<�6X�^��4^P�u�R/���==��.
��j�m�-/��60L�-��C]�zH(5'�do�`m*#�q�..�;�#�Fk߅5$KW��LR���1;;5�� ����e/�牿40ֱ������i.���7���)��L�䊆�����(��>�`��1ӹ�W�����WiC���%,1� �\��o�ɓ|lj�8t��x�E��o~K��ޒ����+����R�eVl[L�&�8p�ݒ�9����#�Ԍ  3����c�m������ܫ3VI8~��	�[�-S���R�)5]<�S����1���?���ڍ�YS��0�	i �S�e��[�x���ru�!�	M������a�2	���K�{Ĩ�y3��Y=��19>�)��Үn��D�� ����위��PC��9W��:0�E^2�B�D��~.��Ǻɺrrz,GGr�｡n&��:��S��^Q��xA �L�L^2;0�(�cs�{�v<>g��su�>|LC�Ҙ���'r��s�\9��)Bz�*�Fh3Q'5�b��>��#f�@�@;�\Л��£��F�B��vbW�
F�i��H�;�"5X��G��uI���vP���rޔ�`�OԶ*�*�eczԵ���iY626�{ ����K�R�V�ݼ.���o�� ����������m�>;�w�<~��%�n\��g&íM9�Áa��-��<�������w!�z�������7�_�Q���\����5i'��D��<M]_-�w�w��J_ٿbr�����/MKRO�%�a��<�27"4V����t]����M�чm���E�X\:>rIiB\��⑍��gKģ���P�������5f�*/�3 5��Tq��Hm�?��&�W�*O-��y'&t��	��B7�'��M ����H��<T��HO�S�NƬy�Ot���
σ��*g��;�>�jiM�uw����cu��s�o��|px���i����\�j�@8�s�����Fa��� EqdH̦�|v�cz/()�)���|�;U�
�(��>���ZW����dLZP��ۄ��%Iwf���#u�;��1�,Ԩ?x��.���O���i�X�42���2:R����"v��w����@�go��la����a�l�5�қ��m-�V��<�'��݂���]'孂2Xے	p�uL���z�)7<9B[#U�@�_����7�O���1bC��}���5;�V"�޻���ס����Ǳ{m������\q���2�Q����Z8S��t)�b&+�6��Ӏ]�ϔ��NYzFջQ�ß�>� �v9�V	�ƥ6"�A 6*�bӎ��ji� �R����I"oTd�Q�s�>,[�A�e�܃�,��4aX�Rvi�
�L�Ue�Ž��/��9	t�R�CJٺ�Yo�7 5C;��N���e��\�Sn���<�x���k8��?��$� ���X3H��p��C��� ���wpp���\��w�t���DO��|%��}�W�	�����ӧ�@�ƨ2��h����c��=}z@c/���r*�����e�
F���ٙ��`�N)Q ��@���%�u��� �ұ?�{:W���e4�uFs���7����Ks}�F���@l��%�J��uA���<���r�����o�-Z!����,�"��W�ˮ�{�3OPh�75��D=�)���YA�L�/�"k��
�Mz�n�2x��0{<��q!Ý!C�b��+�Ꙟq����{�̆sKnD�@��ަ�w��: BX��o��)U�V����e�-��𹀘��@	�G�
Y��<+	^ILL^�h8�Au)�ۀ_1���/	���V��s�>�`*�P$y�G ��P�tH` v�g�F�ܷ��@�gr��5&@"r�sd��)�~&U�)�c��P���\ 3��!������sxt(�����*�$Ps�<��n3�V[��|Q3#���ݼ1�U.h�"_@(p�瑊�$���E�R���la�ݤ�qBX�&�s�~��4n�k-����{��2���3O+�o���sc�ٝ;�ӓsv0�:23 ����+�{1�sD�\C��#2d�!�}>�Z
]��2[s����EZT��w� !T8�&�U홮m�K�����P\�K���W�fkx��nȕ��e��dH4U�X-q�@
6 �?Z�˘�L�a6�p��{�#쳃�>�\�],&jp�v�:jNP��3�z!!U�l�u\�������t;�N-��H�e����cj��>��|���I���:����a��Y�7�'ry��.nݺ�:�F�H�S���4�o����Z��=Tz�ZmD���OXc]|@��2?=y����U꓋���2�\9N ��n�g,�ce.���m:��j�땐�Jw0 �9@�8A1�%vz�qԍ��4Ġ�ĘgKhӷ�� �����������2�����u3��8N��n�Fl�{r���k�֓K]I����Aڵ*�$��/r;�����ݝM�u,>��>�dvnD}���m��������!��A��;����xx���M�s�HQoC�p���BzK����y�����:/]99�ٻ�D���ʻ���`�&r~<����6������;�fsS⟫!�����/��zeS�}����S��\�X�e�������%�G���8(�zT�HK7��˺'�zۈ�Ʉ��:�E �;�)0=Z�<^�w�[������*�+���K�������4���mQQm:���H=�Ao��i��!9��Id����?�@��' �5t���Cd���z�(��A��ij���mW�O�3��A3�d�q𦫹'�փ������-�D�kO�����ކT���t}&DЩ먿Ib���}=\W�P�}���B�@òJz�� ���\>,�B1F��aMm����(sl�0D��3�2��N��(�Xc��NL�j��t�F�\i}�`(��S*H1^>����<&�R#ۀ�VԫD���X6G}
�t3 ����k{{\L�.6��Ӝ�kI%�=���n�Y��^�	������,���1�9ρN�2>��x�Olh+����,�}�IUjGÎ���ȍ�{j�F���w�s�&Չ�w��y�i���S��X@M��Skoi.�39h�K�~Io ��z^��o���#��T*駲��'O�-/��3ֱ����M�ߏ�uq�lƶ&�P�Y���H��̾��Ɵ͛8��lj�Q�\�5��d�ʺ��װй��fy-�;`	��Lu�"�
f�"Υ��[���&�Ҍԛ�ѹ=?���cq�A���Ï>փW�_�ٟ��w��=_��Q��MP�S� HX�daC��W�a0Q[v6��"Q4���	c5��H��ӣ#9S�pU��pVZ<k&�[$�!<=>��g����p��EFN���a�j- ^	(_�D���'�N�����*H��/�&Kmo,JZ���gFF�|��.�(�&�S5eܖ���:�<����Z�/�I99:〷[h�=���;���[j���i�cx��8n˝����g��P1je��(����;�#�
/ (���El}��u�y�:IA �6�h!<k�1i����f�s�FF�zU��dfIv�S���\�[�ݢ����1j���\��ȾA�Z�<ťI8�Yx
I���"'2��s�5ܐ��NO�S7���NH������ӇO����c�ك�m�0�Hq0p쏃ua�Mj	a �s���C!gIm<�_�0��P$D�%C��+�a �R��ȦRW�K���	8�N��NO~p���!m��a������G*�gB-��Tz�o�.0��?�T������d��!f��tf(P�㉳�5��&�LI�:έ�{HB �	o���	�*�j���Q<=?��Oo�#�y&S�b����P�
\]��H���L�(�;��w|��IH�H���vƍ��.5�V�:�e�`��*�{a�.ȽU����Tw�Ԅ�p�38)��¡��R�Ϳ`@�y�����/��d��E�z�	��'O�P�0�f�7�uiDԿ�kkU����#�;S����*xb�
ϰ�9�����U�~|��	l���mJ1�G�C�7���̦���^��׎�#"WcG� /y��6� ᎎ�>�"[�ۺ֗��`AE������\2{�1��3�%u�j-Ą�:�ế�+7�ސc��	��΍h�7�)�?�G�or�!6����D�fm�
�+���RՁ��4��3�S�VWڵ��UXS�E�Q�KJ��c�����q(RsԼ�2	
�p���[�1�;�Z���Ŭ�*�S�z����~t�T�Ùlm��n�n�K�jw��v-5�����f�j��	���Z��j�^���or�V�L���ِ�&J6�$����53
���$�j��sd:��a�a��0 �=�����:�Z�F�o��p�٧Ea���* sUr��s"�[J�!֭��n�o~�(��6�^��i���k��h��/1/v?��L8�L)7�E�H'����G83��u9�S]7c��[:I�^G7�Bz�ϖ�n�q(Lj������ӦRO���쁎�>N�J�:S�sd�w[߻�k=%(�T���YUˈ1a�fb�8�T�BJpgwW.�N$�ˋO��[=�v4�ؒ���\xR�e�p���[h��x���ϛ�#�A�붇L�B̌�z ||��]��*�us[OЅ�'f� }zF���.L�>��q�i�ҼYF��@)�%֯60�AdJ����N+��gVjQ���`�e����'u{�V�V�Tph��85~8Qeu+l^�v�Q���T�g���)�V��R�����?�BU\T���5�#�ʕ�:�)۔>xpH�,���C��{C��SNd��԰?��&�,�|��d��[#���c՟'-<����l�4)�Ĵ��X�"����ac@���D��j&�9_jD.oY8��^���=�"��ڻ�9�e�g�N�K�+]9`F�i��R�O}�^��b!�ڭ�)e�JX�V.Y�VeW'n. ��`S�^ݕݽ-��U�`��+<4����uy���(���}��\,��}$^��
O�@�J6 ���)�[���H x�M;� ��I�;�W_���ZN4�)C��M���LP��a󠶞b�Ȼ����:��X���n��'ަ���
]P''\�C���lB���`���q�a��w����v�	�jT�B>��ї�_I?:�"V�������G?�Gyrp!�܌
�26%i3�7�\�HH�_�cF s��wa�"�V�X���@p�2�dI\�p�i�B+z��t*nhX� !���Rh'�:1ۅR̢�2=T7oo��O����Hf;&3����F�V�n]� 1�&�������3ti��j<�{�]��׿֍<a-B�+�{�!LD^
��ԴFڦxvzzLwggO^~�u�IҺ*��\�.��{��nI�� �A)��#�`@d�	���T�m�1s�.;6ʗ�3���X��-p�(J��)�kC�=da�ggĮ^�s��q�P%i7x�il���Za"7e�h�%+7�4f�MA������+/�+/=�%�P]��_xN6t�����?z��b���5��w�@O++�C*��(�_9i; L(h� B`(P>鵨��9�	�Ű� gOO|d7��}(�ɜ1/����0v����uH[��;�6�Kڢ+��V����FuF���'��7��M���59��x2F��z  ��	��c��;�
a�����矓������M)\4T���'^Gv��J��&Ô�����u�qk_�����<�w[�N����4"�k���Ƙ��'Ʌ�?eX{-}iD�A�]$�Kљ�BL޲~0p
�FdmG�+n|l>(�Wj��j@#5�S���8#m�Ș.E[!F�r��{3�����b<�����koW�5g�Y��Z5�
�4$A0��'?�����[4�(���Q/P�W^yYn޸N��>8�@.L� ���ɍ�7u��c�r_(dޖu��轶"�Y�U�@"}����߈�`o���x�}�[,��RQ�I��~M��Դw�z:��Ɓ��5N�X�X�Ƣ+X˒ކx����e@��1x-&&��YL*I���� '%c1�x(�lBlnY ���!���'Pz=H�[�����_�Wr]>2%h�=S� FX)N��)��y�����L�d����`�$�~�+`sN����v�4$�899��w�T���/����ʵ[$A}~ck��������z��I�@5v2����|G�G|*����إ��Vcv�'+9����KƼ?ؒW����==��ɦ���]�\�1��4����;��ҞF5�đ�6;��F�������02�vwo��_�w2=����#�zIg�~EZ
�Yv1e���+[lV�T�p��� Tc��Ŭ{ӰȋS���
�+?%-��|OEl	� �Xo��DɌ�t:�ٲ��� �ykQ��P`׃a	[@$y�:�X�у�����v[�v�/���Gġ@w����~On\�*�޽-?��P/�j���zg�/�^�µ�U�7oܤ�%�t�`�bm@I�U�ۗw�����yG��ǲ�3`}����u�����>��} �ŵȺ�;DX�u���Ii�Uy
��.�^�B��
3���!\��Q���3��3tQ���-u�'�U j���2̶tЫ��45 .km1@�����/M--��5�³H�9��̍����g%�XĦ�w�������Dr!7���n�xy*�Y!5nn�h�Z�c�P�xE�]P�a��9�z|�M��c��N=}�X=z����o���lv�d��k��+��'���a
��Ŕ4e�vX��P�q������������~W^�u���}�'tG]b�>��#���~.���w�]#=F�d�K�}[M*�r:ַ����G��/?��g/��ɹ\������`�����r��Sz5W�^#����|��j*ӉU���*�
ӖI���n�Q֫�����7t�uI�`(l�5�GY���Y��?��Pb�LL�5[�3�qQ���,�B���E2KV.p�V�l{6]��vL�ъ�����~�S�.�68X' F�Y������P�ل���#�`�i<�~K���O���'���=��}�v}�]���ߓ����/~A����7���y���TC.����Ԣ��F5u�F����7].�QSFFk�;�6�y)�Q�^�i�����0]t�*������gMG3[��&�XoX��BR�4�_�;�d�j�=��I9�R^��������=E��Z�؈�I�{8?���Ō�C�j�t�?<��E˭wղ��a���qe&o���N�۬{��A֣����ӓ3.,����@Ճ7�Qƿ�����������vv�<zz(�|��.�����ȅ�����;�����L�^�fx*�������$*���M��7��?�Gy����L����L����f�����jhX:І�����-�����{B/�T!w�<���ۿ�Ax��7��?<<��!��<:↤fn��LSF�J�2`�i� �mQ�U�5s�Yͨ�.-0	ں�sX��� �D��MD�}��8
�(()�T�ȳduF��|�Z�R+�A�*�X��vb�Kfmj��С��Y�|����x�!;�̰��Z_��WRY{����g�� R���'���z���{M��	����?�^C�D����>�rY2� ��I�&<�p[��Ъ5�2�k�R9�!�5	�V?�
�B�x�_ʶ�i���#�����0NG썋+i&��d�����4X"V��1S՞K0>�'�<۳VmQ?\�I\��Z����'�u��Bx��G���f3����#��c=	n�b6'������x��������UƢa��v"�|I� eW�O)�8y�򖘠/T����g�62���_�-�|�k��F�j���V<�Yv�
�2��b��Ԕ��+����a�uu_��$���?W/������a/��v�5
t�v,f�N<�(��JҲ��~(�o������ ��>Ɵ~�)+�������6��v��#�	̊)��=��ʳn�]c��>ˑq��f/���!���B�3\�2|u$�X%�v�H���gUm�h�v	�f��"��������9X�9`\1В8�����L�gk�uM��.+wwv�5� >6�����9����l�9��Z����X�T����c2�a��s�P����{���/�50���
_a�2�vH�0�EK+C�/�l�X�E��(�l㎿I��u:Im���~� �����\�|U^J��&�wł����׳P	-���4������,�<
��[J�����ء�%�����^i��X�/0��ّ����T'JS��;Ӱڠh����C�GXg1����Y�b��ƉS�?����y�ih�����=8:(�B�&��X����-�:�fm5J�h8�P؅ЀD�ed���0�w�w�S�t����Y�M����/�&×��,��z�f|O�B�J5*��5Ss~i����L�d;���귃�*P^c�N(}-���ӛO�0+!�%P��R���FW��27���u�������jZ�`���IůbSa�],t��	�ǆR�J��;�h�e�0Z��z(}��&�+���k�Ê�������nB"�� ��?����O	 �i��u]�zR�f+/�[�Q��-.�Ա�~�g�0��б�kp8Gs���Jz~��C�*������� E�ѻ�>`Lf���w��9s�1xE�[c�d�����l��y���3�w���t�0��?A1���FnD�E(0��I�L�X����m0R$AUK�ȸh�����Y���Qi~VC!q�vI������O��_��� ����|+�C��T��T���e	�@"�˒�YPb "Ҁ(���cfZLR�Ҽ4�a�@<���j������bނ��_Y�7ǖ���E�~��
�S��*s�o!�x	�H���v�:UJ�W�j�=J������a�2Wqڶ�p�f��R�Z�	Ұ)�����z�,V��t=��)i�:*������[��Fɀx����
�F�μyȰ�.���y&ۇg�$���6"�VS��Z�p=�k��:V���1�3��	�S��� @b����G(�0H�GV�,�Rks��|_"}��|��D�)s|�T�l1�'O�Lk�3*w7F#�#�6%�Tm��兆§Σi�Q��;�|�Z�O>�\�^�J�e	,�p.PѴ~�̑խ������α�.����1k~���|-JT98��U<0�9
�DMV$��xJQ�CmL�̶��8� �H��$j<���)V�K�%ӂ��/j^~����~��{������"d��:�N�%;�E��W��f��-��\c����	��B����#A�5u���e�`�`��ҭ��j��	�B�ަ\�F�*Vl�P�G��6�8"a�D�<s�����+����c��p�%�����"������I��		��BR���
�v3�k�b�Fj��`$-���u�!ڃ
W�	(�Ě��=^���!�P��6e1[uO^��5Ϟ{{�Mյ�[m_�K�H�V��2���ڞ�!�6�T
a���Po#؎�Ƙ�K�2����)J�5���r^S!��,-�2	���q�bzP磎����(m�Ľۤ�#�����P��v���K�l2c������̡��c��Ϸ?�LC���,���k�-�b���e��d-;�F#��^��y�Lle�}���m�~�:��<kш�#����XZÿ3]�hw����#n({���.Ц�m��M�'8E��U��Q�ކ�h�OHʜ�-��iWRl@L^a}= �R[]�r�
�&��Lb5Fn�0<*�g� �@]	�%�u.��ۥ����^�S3�]�H<�2�f1t1GҌ����/qjv8,]A��\xW?�B�����a���1Y�%,�N�@m{��객i���B�\��p�FIcW��^{�gF���<�kӐY3���SK��m��Lk�{&Ћ�
X�{F�4N����[�~���*������&�ԗ��Y�� ���뒾�#
Q��ؠ���R��c4mt�V�56˃1dY@�8Y�d�6�p�A
��E���V9�|��==ՋyE��V��+�fsf/���M(a� �Q��c��lI�7�M�!�rNl	��-b�=nY�D��T��}K�!�Pw�Ƚ�JJ�,;t>�z�t<#���ɚ���_�2�XA�\�%����%K`>�l�Zt�&6e��Ctم2�����[��������ro�9��gm8jL$rɜi4ˀ��(5�y�J���g��:�Ûd6.���8R�-�gCn�75�
�	/g:394I�j9�t�v].�J�|��Vi�Qb��*W\cqZ���ϋ�\0&��3Kݚ@K�1.�y�%	'v�����K�سM�^{��*��E���Mײa ��K)�:|��ٴ:��ie+X+kC�5N��s��c�;P�M���{��4�H�E�����<4X��PIם���uJK�P�?���bкA)�:�}ш4mC��u��4�M��������c�ǖ*�1F��tf�"?����<7�.7���8�3�{��<=8R��企�T���5�;��t#�I+�y���7 #H���Mb�0��D`p`8V�v<�^��#j��sz|,c��f[�2�Ѱ����u�E��J����aN1� ~q�$���t�2x��)5�:�����do0�"M$��D\$�^6q(35��S]Q���O����*�	��`Ǹn��<�ɯ��*�S(�o����51��98����ţfQ�O�Q-���Z��tR�Cq�/�wD�$�7��ݥ�`N��%a�FcD����/^��QmD��i���.7s���?�fM�I��Xm�~���{����#@`�[?O0Hh- �]]z�����[6�M���ӿXg��i�P�0�J.?����U��Ū��1 =p�l�&fK�.�x @��2[��� �a
�V"�t�"�r�ʶt��F��Eb'v�Lo�-j�"}������s���cڦH�� bD�ʾ0`�"��~A���]�N�v�a�������ǬNo�}z�K��eb;�HL'�/TXgJxhm}�S��\���5@5�)I���Ű0�'KZ��4�YCY���r!u!�3��h�o�0?�io��.��h�l(ZAĠ��Zơ0� ��5��
�y�k'o��%���` �&m������ ��5�ć�j0,Mf+tlJ���6"�#�7ϗ�k4�[���<+F�����d�Bf���5ø�iUj�p����[H=;��+�M-M�'[H�p�1�ڒ���Z{"����Ð/�F��믱#�,1%��T���mFB���އ�]��X�.�;��wX�K䩁�^@�	����{|o`AS�,��rxv��X�u��t���7���H��@���}�re�X��mİ� T �B��0S����)��W�5�q���e����Nj��<����ӄ�(���[ְ%�6I7� �bu)��2t��зƠb�ya|�E+�`����4���gP��:(��|TU]g���K,�GK0XK��%�
/4T7nD�<�7&�{z
EK�g"��\'6�"�ک�	��i�p�G~��y�����-�f���b��Epϛ�oͷB��V� ��L�N�9}Y��J#i+��·��f��j��at��*r�*��ĳ�q�P42����F��������Ge�`��yT5>pmL�KB`/�OcMC��eq܄�b�~��K	�c��������:]B����g�Ƕz<=�OY�2�X�4��S� ��*����=z)�nn���ߒ5*��HmP�!�es�%c�Y�ܘ����o`P`������!�oLj<#�z#�g�,�/:qg -41�KH��D�0�/f� Dv� ߉5���yj�5�.Q�V+���3!U��ik�P*YK���ŗN����PՉ�Ph�02�A�FI���JH��BP̦�NC 63E-A-�m�*�&�a�VI��C����%0��-���k�a$�wV�tH��1J�MmB�g���	�������7j�U/�K��i�N�{
�����>qsX�@�C�d|��^�C[�4��2��d%������W��Y�F��OU�exv��{�n�i��v,��H�Ł\x���ԒY��=s��Yo�n����ځ`��m`T6���,�?��\.&SV3S�!CU��U�0�}�W_}Y^{�5���m��6�h^f:��|-<;������P��6O���Yq@*<�XG=���;r6�˧w�d1m�D��mds���!�i2�t�sҕ5XS ��ô�r��⇘,�#p?`�"e������I�J�x��$��S�H(�5 뫀��;��{�
k;��EdIhG!b�$ �D����[D4 �C�aY-�)��!���DdV?�͂Ǟ	�B�qn����u�c=T��n�u	װ��w��@Uc��Jճ��x*��	�d ������;��K��1�S(�����7cbƮ��B43*�3m��ō�� ��tg�ۉ��(ч�-�66ʽ�x6w��:��s�b�Կ�D�
I[�ME�O��<R��ܫ�ip��&��=It��\\�f�x-�5�7� <�lZj��g��h���8-4�ؖWՀ\�q��<bH��c�q�a����lnm�����2��0,�&`�^PW3mH��f%�h{O�A!O��Z8TY"�$Od�@�=2Y�2�"�];��;K��mj�i�0 k��6�f�:)����]7"5xʬDI�U�L�E�TQ=�~:ZW:��z�"~.�k�����4``Hd��W-�#s(��ͣO6,��`C�7֠���%?��>�V,�P�Z"#�D4���=\�\똃�Ԩ8���/�$i���,�aX�&mN�{��c����F.�s�Q0R�@e� �����M�^���e�՞q]�r�����	��3�P�/�XZ+
���cZZ_f��@�b�ݽ����ܣ��0��u�G�g�kϲ6�a��U=/�T�V+�le "B��I�G"~��v��g�H<�\ �)`�j�뵱�Q��D��c��K��:�-�r�B�Ԁʼ8�� ��]��/\���������H��7Hu�֍�Ql��U�;�"x'.�a�L�]����=�q�� m��8`,�`�}�X4�����T����Krx����=9�щ;QAO`�V�f:a^}(�-�3bz3�NҰ�|)J��y֧����T/Ġ�J�͔GsZ3���\�UT�������Bz �u[>�&��I�b�������&���������z�d��Y�r9��l�gO�0F_<����uO#�6�]�qO(��mүa�B���T�^��3����G.{W��,�,�a�^��I�_���#@o����B��j0#/''�n2fF���4|�wh��ʵC�'&އH<�ag��#�NA�Jc���qCJU<,q��)��J+�;�u]������%톶
ByKP�vJ1o�n�N���zK^��a��tZ�;�!��^ p�q�۹��!�5_!�a��=.
)������ʖ%��zX熙�����F�	�2��`:;���!�#�B�3��z0CG��O���D��d���;ﾧϟ�~�8uqL?�-A@��R�<"D0"��~);S����7�+g�sX������g��1,��'��xU C|�W��FDc4�7��d�M��ޛ�ı1�W�2,�hD����ܛ�E�#pլuL���?�h2/i4=��6�zxAi�	�9��:����ZQr����=�g�$Nw�쁬gv���^Ƴ�nH,�m�V��=4d}\��ח^������ ��C=�����'���4" ��3.�8Y�|k�	 4�-�Z������P��:��\ Bd�2!��N��n����O�)��b61�\d)�����)|K���Ǉ� �En29����
���� *�,��,�RA]�и^�'َU_�������%�}���;?���пݰBХ�&��;Ò����g�f�����w���Lv����g�����b�x���2m�����uHR��-���`Db�l���2�Ce_Ð4�h��&p�G�Nv��@u�P�`%б�����"e��ٛ���t���ƚ���f�`�~�u�V��gO���r�m}q�1�����X8\����\"�F"<��5���P���a!N�E2w��������h���: �>�5�7+�M�v���p ��jRϪ���+Ӿ�gl�0���(6�$�t��F��F`�Ks��閥�1�y�Q`Sۜ^�gwۡnOv��E�)��4�~�S,�Ge�&cu��w�Dv0^/�GdK��gԁm�X��v�����E���������\�ڥL� @�9�6��P;�T �C�>��sn<�d�`��>��T�5V�}�? �ô�/iH�,EH�|�p ����,u���x���N��N�h  �.I� ���Ҹ��R�Bi@��3�&���[���u�4a�7�$�?��ڔ�u C|K	;(2���Y��·��(2OL'� �+��6�������5��hVW�<U���Z�%˽+��S���C5<�@	�1|��=OI����/Yg�s�e�#-���%53����2�'���d��g�	ռ�!��C�f�I}`���.���ִLW��_�b�ڵ��^�ցg�İ��`���W�5�8�_���g\V�q
�O����(�������`�n%a6�q�2�{F8��/�dn��!�����q��Ww I�pX�(���l%]��t�V��Z����$5e�t  �V-�!|���ﰞ���
�I���:��������v���1��E�e$2�dE�젯,k�ÀL���$�0����|��l_ד�����*k��
)�|� ������e�#��Ӭr��� d��kn�scig��R�{I)c�5D�ו��6S���Q��,˚8���7iU��z@��p
�R�l�M�&{�� *)�uXR�^A0:�`v�2T���aCwp׍DC�<?��6��L�����k�gXӋY�\�Y�?�q�y%V/�rz4؈M��|�֊���P���	_�0lb�҉|E��UU�X5 �H��nB�K�MA���6Ff7���y�,^փ�٫E����] !!����<��x&��������S���X�����n���cy����8��83��tl�<�F>�B�`,�3�A~`6[�H� �+99�ç�r�ѱܻwϚ]�=�����}Gh��4v"],�3+�=�g�#��l�0�Ӳ41$����*mm~�e�/"�4b��p$g�I�xɲ$��p, 7�����X2�*M"pS��3.8���p�,ͅ�d �:���bQ�{I���tŚQ���U�6�y�}�}s$��Xf(.��K�H�a���X���%�gtV|����.	<���H�I�>Iy� �!ӳ��Z��k�TQ�:;S��eCy�:�`��2���.�Q���� �X�J�S׋�� �q5��D���4Q	�c������k9�zMu�:��ƞ���K\Ka#����A�d�����Һ�1ti�.	�*)��:��ʝ;d�E�7��Y�.O�Ń�W��.J5�R5l`���_�*�Z�z�U�MC���ú,�*�K�*�q���i,����y�U�����ߑ͝�rr��WbM�#�4g����-r�U3�!4��XI*��Vl~<�f�!��01�>��u`�*,fE����M�Zt���l��?�ϩ�QVBPq�%/B�'0Mi٪�UZ8jı�ZVV�c��+J�]��d�<�8dhT�5��դ2U�(�C<�z�wb��j�ѡ�kU��,3iүnR�Ro`|�	А�j�E�5 5���f��9\#r��ِ!4�͙�H�b3:,�b̈́Э����ó����4I�Y����PЀE�%�*x0�׬�Ӈ�;Jj����َf&&Jk��u�,meY����;��5I��jH��2��K�[�8���%�v�؈ ���{ߐ����X^}�y�\AN��3u���L ����Փ�$��9��]4aϱaڔ*(s��У9�<�X(Q���������ѷ9�8P�32̰��JOT�B�s��,	��Lg�u��E�9{���(Y�]�y[����]�A8$+'�Q�����/lӃ˄�~Τ4�E��(�&�_Z��-�'EF�d�b$���t/�%�#�U��� h���2c���hcQ��"�L^�_�>�z��W���5����M��+I����:�I�,F��uAs���T�����+!��c4��)��NGl��و�
���Ijb�ե�4�Э�7Ne�\���t�~V�xE�mµ��eշ�٘�|{φ@f[7��#Y7B��O;��Q���D_L	�n@���6׊xSM�Z�Y8�kO#r��:E�����'^Ǵ9���H�ִ*����C�Ex�#WMXK3�s���Q���ZP4�ړ_����mʂJ�9%%$s���}n��֖��BUhƎ��xOJ�"��竂�et'�zL뢙4t�t�V�ႡIľ9��k� ��+=\!�D=��1%�d,�Rx���J�s����=��?�����c5f��1�tƱ�y U�Ӑn[�'��T9�jD���&����aE�O@�*|^[QT����BM��%������%�q&YU׾�l�6h4<A� �I��ٙII�1;g�9���{vٙ�G;Zid(:�"E "AB �u��������/Lf��� G#]��s�T�����/�u�
!�������o���D.�Pq�y!	o�R�ɍ��a@��
Y8'
S�[[�L�$�dE)�,z5���5KP�)i��l��W�޶���ܥŴ��+��by)g���qQ�Y]X����!/�c�Q=��py-IWÊet=ٵ42�����D,�r�%euR������aK��-\��k��#��~rf�ણ����i������� ՕE��*�u
�:'�-�� �bcʘ_0���9���=��}r�N���������Po�I��M������a�;�5�	����ϩ��K��9MBȱΚ�]::=���XG�y0:wn�K����E7]�,cY$�$�m$�W!�Og4q#��z��D/�Sf�vT��Pok�I��E�C��8�!5��m���@_��>$����$���x�6�}bവ��"�85v���pm8�kĕ�g�'bRd (��Y�GGG\C#z�n��dG�F��0���bѓ�Q��1���
N�w������Ņ�NXI\�}gEp[����Y�ǹ��L�7y�+��E"��F3�"=V3"V{"�e���~("�7��e��d��u�7�w 2��
�H�Y%J��D�H��6b�#�w����W�6���ً�=
�Fi��ټ�Q��
�o���$]��~O�9�y����;���������9
몠������>����O���fKQ�cOw9���ء�`0fg�9Z���x¼�gl�-,��,&��n�>&s��~>>�y�p�����撀�$��Ӣ\��g�I�C���k�n�G�?�1��������xm�i;���I����+Z"Ms�(c�"Ή���(ɼM�YB1|v�ob\�]�k� `��Z�Ft=�B8�bOF^Dj�HC K��� ���h��1އ[F�+&�Z���[W��Nc�CU����U��w��'�Q��<���:3&�*�7\�l���򦷱\�i �W�F]���,I�R�#Z6J��L���o��Ĉv�@ڜw��x]�m3��Ez���x*�������i�Ë��Rr����C���ĥ�Vv����77
:ق�E�S' ��MT�V�8��$���o��YC_��g�˟�8]�]������S���|�ΕY�Q�l�1B�2l�Έ&��R,��yM!�xY�8Sv(N~T�b�@�t,*��#�!6Y.���JFUx/�}�PpWi�Vd�fٜ����C&f^���S#?3�t�Jha\��Bw\6�o���I������u$������Z�n�IV�8����	�C2-�c��)��B�@,�F�R@��ܠ����!g��/���Q��8W+��Lw�.W*��S�Ԩ
w� ��h�2j��5؈������d5!F��PB��0Ԛ�Ā��o5둊�gH�X^�4E4:y(`�E�|C�9ll���\���<�"��i�{]��݋��H�&q(�f�ϗ1����ik����X�!mx���y���p��4σ"��i4�2O�
��3��YI�Β� ��W����_��y�&����~�7�駆a#u�d����q9M�m�^/I{�.��]6~�$K�/[*R"�g�dtt��Q1��y/�X���H����~	n���F*KT6≘�p��Cv���-p;Z���\,�p3���5SDb��xu�ueF[�";���/2�b����-� ��O�\a������=s��'�c v���"���*ɋDv��^��&wZ-lS����=PG#d��B���Ι\��0(ux?���ǩ����y��(��+l�Q%��n����2va ��Ս��FQ����r�y2�.� y����u�4@�/�@�����7�i	~��ҕ�i!=�s��~S�{]��H�
N)�4�����5�q��+2�[�*'�t��~�#��?į�D��D�:��+m�{�N��O���૖��_{����o���(wR�6[6����#�A>U��O��,��-8W=n@͇Zm�����2�=�!�y�v� G5�dɿ�Ğ��j�h�ءSp9B����R���CޢZ�mH%8��+t_�I#�b�*C�����.�f�0/�P��9��78��+�����=R��d.EA
jɉd�?\��7�Ⱥ�c=W�JD�9������ .�?�9��_�|rN|�b���Y��&y�4��2��{g�3���I<���,#�a��š�S�h��K0˝\�U�&?��=�ZnpB�٥�ޚ�|1[cF�6��S����:�tm�P����K�U�Q6f��Pdqd��`!��͜5��2q |L�6ދD�]� WW3���輘q��S)���2@��Tŵ��d̹�s�)�h2�?���ӷ~�:�?��vx�>W����:]�*�Vk�H:���wٳ�M���<��7y�9�
���I�	|hY��O�\&�G�=��h��=z�eC�:�RQ+.��b�90�^���xt�V����V!���ymdQ�W��e�i�XHY7�>h�
���#���H6s�^�'��R��K�N��/9�+W��n$MP	FH;kaB����Ϩiw{�C `"U��ٔ{�^��!e��}�-��@:���%n|�F9P�>f�3�;��H�j�Be5�w�_D&T�?.n�xڧ�'Yb���R&I��lS�Ml�k'�@0��^Kϵ.c^ûd� N�S�V6��)>w5\Y[3'7.V����37�V����2۳(���r���O� '��bC���J��A��ƞe��W;w��h�糖N�K�/���cc]�E��cܑ����N�����t�=���8y��S�W�:� � #f�
� 4�"<��+�F���+�|f�r��V(bQqFx����Ъt���V�	yR�^�x�I��{�@r�б�����cWJ�ƅ
[#b� �<�,���mE٬�>�|Qh�3�p�6��[,LN6j�E�Vw��m!��[�r��ݤ��S����Pw9�I��=���n\��M��߻G�<��p�Z���sz�g�@?|��p3���q���� s�sQXϽl�a����"�U�a�[ţ��e�ZҊ���I�AI��d��fBji�,�z�#��譧{sn�y{-eO7cja$Ј�Hnz������k-;S�ɋ���/���%��'2ɇ{�(吖��q��>dl���hy~L�>gF��1����p��`�J� �Yx�_R�������������|�8���h��5�:+����Yoeޔ�O��D���Wf,�`�xO0=K�K8A"� å������=�a��
=�.x�q�5vI�ap^]����s�6�?��ҥ�?�Q������$]�aIQz5��FkKI��1�C�XHE��q�^�ܼH����tBמ{�����ҿ��/Q�^������`�!�ڽz�ۗ�s��W._墥��������L��4�#m��^Ғ�;Kyq��)M�_��?l�%�!���a��{�BN�|��Y�*�r���ɵ��0�#>b�X[��c�ow��=�V�kU�Ѹd��X��H���T�3ll�GY�04A+��{r}��+�ԫ�Q/���=t�!W�B�p�ӥ���L��,i3�QT�����аZ�go������m���`#<��:�-i<�p}	%㹮�5�Z* ̵)�ڙV4s�C���C.?�|��SF�Jj�^�d��l.�����'BX�d4%������\=��7�X.���:��Ȭe��!"�YBS\f5��.�ڀn�ۣo~�{tyg�>��4����_ܤ�������{�y������[�z��-��)����'t2��x�ȅ��1��¤\��d}ccr+�ٛ��vuV�h��<"��gU+Jgl�bc�e�e0�3�W�F(�>�^s��{"�ڲ�q|��jV��<��˺���%��*�c�Z�2�b��?D>�����r?x�و�ͼ������~��ŗ^�Ͻ�)f[��_}����ߧ��5h���$�����
A�K��N�������M���|�~��ѭ����O���(����8E�����),�r�/\*Z�*nt7D�Q���=��e�}��`��l�hq}�;����
���?���<x'l/k#"�J�,�*�����'����Y����{�m�=����j��$�E&�/�:���(:�3B
����_gի�_�k�=N�����W_�/﹔Y@\Oo�s�񂪃>>�y(
�H�.��$F�;��-���EOĦ�iR1���)�X�|��fXLY3�eAm�$����!Ʈ��b��G=�A����x�g��ǯ�*�u���5�R}g!mS'̬����}��|N�+��Xo��^�:�^�Lol�K/~����O�'��N;�@ꏶ�\ߦ��}���>�=`u���z%*��ɪ���=����������l��m��k���Wߠ7~y���Q��A���fQ��q�Kb7���� �'u���`nH��xif����qf��(��4��#��$=�Ll�e���o��'� 0 ,���y���$o�)W�"`�bsu�jOU��	�̈́>���w���[�0t2K
�D&˰I�k���go�l�-z�'�'o�F�����!Ɣ�z/\Q��F�,[�q8)��h,�����G.H����u:�
\f��5UHi$�\��0nkVh9�lD�֊0+��H����f�L���uZ�v+w��@f%4s+�����=����k2$�f�h.�
��#@�zՀ$ό�j���n�3f���Z���P����;��o|���W~�v6;a-����]���շnҭ��;�Ă��Y�X<u��y�|\/pn�=�o߻G���]	�ƨO_���^x������Fg��X�Uj�f��y�
��d,,D�1 P�1�n�Y��JdE���E#be� 6�E:�.��N�R��R��d"͠�L�h�.t��1����k��̈pڷL��F��\Ѹ<>�C}s6w�
[���Pg�Q0���\�!DY�{?�	�~���9��tN�`w��Ω\���/r���5���e�-ǰPU7U
��Z8%�6�!���p�]��	.�Ri�������d�l���2@&U�<�3�$_j~��o.nR|_�Ǆ��̖�EճBbk��Կ�q�F�C�mİ8�b�{X�Ģ��)b�g�Z�60 y
��3ڠ��QcT~�i��)������Z���o�3�����[m�M�m��J�*�f&x�[}����:����9B��޻7��_�~��[��w��~X�%�"F�\r�eڔ�_��H7�����x���������z��'����٣/��<������?~��.��pm�\.4�W�-�o��U�����5�Z�]˞�A ���ڦp7�N�`{����ep�Ay�T54\PE�!���x���C���J�ݼ�P�g=�V�� ��sGj��`4��6R��"��+_I���[\��DTP�[�M���T~��v�E��`BZ�(�50`�4
q�f�E�p�k�W�q	�+��;�pi��/�{���h��I��'�wvB��C��n��p]*��$ ��I�p)r�a��k:,�pC�hu�����C�@S��i�L�E��ִU��;��LWɒ������¤1ݻET��E��d4˞���}/�=�F��`~�T��5Zf(y^"O��������$"�M%�Ie�~�j�:�v���`K����tRA���r</ޕ:���:̭h�p�9�H�EA+�dX��٧��o}�EZߐ
�w����_H�}�t�hΓu����I��0|j��a��3��N[��߽N�s9�������T��o+x�����޻7�N0Ph��:δ�7"��rn��B��"jDmcp�7>7 �^ V-c� �N���sY������h#�B����q/E@W=h�4 �N������@�o�2�J�v�W%�j���V�� y\`�dFa|>��Y�lݰle+���:D�ԮB�Xk0&hT铟���/~�v{!tY쳇����g���ɱ�n��	��yp1ߤ�_�1���T����3�5nZ4���4�z�9{=��X�f�_�$�*�\q�WNҜҮ!;�x.��U�d\
��r��*�Y��ϔͤӻiŶ*p�Jr�,;��qJ����2��<��$�^M�Q�'3��'��:��
�a��lb��b0P��)�6xY��H���`�1���+L��HQY�� �k׮�h�u�#:<:���������W�x���0�G}��0��l�ܰ�Ѹ
'j<��p���������e��rB�?q�6�=��o�޾y����_S�T*�#Z2o$.�.0~�T<�c���p���ůL�0,ɧ�3������1�$B�ŏNz-����i��֍�{�ȉ˄6��2�'����D���т�s��tY��a�F�Lb���P�Wb�#�ZL���+Y��t�B�w
qy�@c�w��
n'���L&�������'���.�9^g^�b��!���N��O��K[��/1�.��.9hg��H:�u�3�d�6��?��5�����yc �ո1�=��.!��7�YL
0m6ـ�c���D\����1�0R2��@ڌ�"�4� 'CE�(�i��9��j
M(�{��E����/��I�"Zҁ���{��
�	�U.�S���=��-��>���2�ׅ5c<GS�p@u;C��s��=z�o��:���p��g0�R��˛�ua��t�A�BD˹x�F�y�]�+?����t�ɫ�'���<�{����Z<V�C.��y̘�j�n1"1�ױ��y1�����{.�� ݭ02y��Y��&�M���j+^����^�Jo8���Uv�!X�&��e��5�@�ͩ=ǚ:����lT�W)�%�m��a�@��lm0�����鷿�iz|�����,h0���2>���M�[[��t��>�����O�@���X����L�r����A@	�Cݞ�����;��j�H�D�@S�N�U`3��HD��Y���7��gmb�PDɪ�o�^d���"z
�K��>������x$��������j��\�{5IG5��V�#ۓ��A�� 쎨��q�37�l�!�$�k��!����Ua���i°L&cft�.�PW�Ya���|0W���I;� �)Á��9�&ܓ�}:���c��4�ηlT��׋z	㽳B:��K�49��(���aZ��Ĉ��y���|D-ݪ�J�6y�UJ2�O>�'�ȫPg������$���U�EU�K����FD�K�4�,]@�Ŋ�ի �2{�ċ�����)��lL���*�z���]�8q&-��>x"�S�������F]��I�z�)N�}巾LܹO��:��X�#m�.cQDˉ�O4#�c6O3��n53m�)I���_	Ad'�����-��d��RVY�n�r
N�*5��^�U8"%����&JY[\9�5U���M4o�Rx��*�fQ$cd��UCqq���c��;�����!�æ�CIs�?�UaN���4�8$���Y��u9k���R�_8Y�@�gs}�����&5N��-~�bz��o�*\�f��������{�����WwY�k��{�CضIgsI����A�z��y�AG!څ�0�Y��qr���#�%�*��VC�gs�o�=�:ƌ��]:�7t*�%�i��d��>fD
cW��&�Q��X�ԝ 1z}|�Ec���'�E�_��F�pN�ܞ5��x1YR��?��w��3Z�u�.:--�g4>ڣN�8{o����3W��ֿ��{��=q��?�$�|�'|=��)W��l�Y��F�g�����J_����nj\2`��B��^7�y"�#���Tm�{���JJ�B�]�D�_���p�B�8���Ǟ��� Ҝ�r���VUf0t+�\�a ������4�r+�M�^"��#�m�m�>��U/�l|�\�K�L
35���e�x>:�i����9���y��c�����]��?����O��oݥ��.�`�
�,�� ����?���J�����	=��I����7��/�����^y�'���~A�E�� �TYm#J��m|�0!�t�`9�_�P_W�U�`ٛ����LF�5���Elq��*Yu���G�M�X����pu$ȉ!��!d�w��3${�`"��K���gV3�g�"�^s�e�U���zNi.GD�)������р�f��&�)}c :0��ԯ�9����Q�\�%�4ǼI��K!����d���(sGb�6�s�2�B����R(��%�,;��C��|d"�Ln�4��Oh�T~e��lߤ Lv1x|z�}o��Vb$�Gj��L�(�5t�w��:[�����/��o��Gqa�K+�벐S���yr8q�?�w:����7Jv"?���_Y8<��[�Oo�9��?v�����|���	��O�E�{g�����=W��g�b����,�����.m\������/}:�=1����/�����۴��pY���UډX(j���]p�ty���:�a>�Z����,����ͫ'�8V���A�%�XQ�^e�*gd�S�3�NP�=轋}C��.ַ����,�C�iP�*ңZ&��85��x�8V�؉]p�~�K�����)Gf՜��,En~9�*���<q���q�p5���.�s��)�l��h����f��ˆ�|���\gO�����^{��1L ��"�YV��Ԉ�]���ֺq���5�k,�a!N���
x�rn�eN��"�ڦ�~3^��@3*f�%�H�*�,I�V�Y#셚J��)o��RA�2���Wz�T~bJ8���bo�Kf"��W�6lH��]*�Xh�)?�}m鵫Ɍs�V���I��pB��[������ͯ��Z0��3�}���K�޹�&�5�J�a����v�0X�ؠ�{����F��퍵����_�ݫ����IS��ں�����n�ٴ1��"���ڄ����<�V5�Mv!�q�Ur	��e+��n�� ��Ar��5��h�bk�‹a���T��ݮ�A_�ׂ�@����5���^��b�j4�
�x/��J�7�jIBk��%��8�j��B]a.��2K��lk�[�"�Q���_���¯�����f&��pI۳�l��������v4����h���O~J��W�p?x+��yx��oh6�}R4�o�ؤib|��F�@� diûH�y�%��M������d�}w�������^G~}�Z)|D�WF���	��ߧkNu�n埔�볱2��"�@�d�0��J�W8�pjz����╸��+Wo7�� }��f~,%z>[�_�ͫa�{��׾J7�n�3�'�~�^���1B��f> e��!��/�Y��X�j�BA�����o�E/��}��/���8<�O�tL����G�����%�uˎ� ��GV��qE��;�Y�SP�=`Q�8�Ph������R
-@Z�H�灤i�x�j�;�uao�,%:66���g��FR��6"^�p7���Zѿ��[�[<7�x�UX��x����e��E��bj��fð����]�~��]ۤ��錅NZ�h;T+_w��eD\=
����)���W鯾�]�����]�Z=��E�t�a���ֆ]�%Y�Ȕm��,�DN^�r�%mȜs��3]/�(�gA�	��6��;k/$�4�����q����k+�Q�j
y��4���S�m퍜�C`d�N!$,gڢ�V��(�����̘�>ZCYsE4"�p6���3
�+}�_�&���c����s��ÚZ@�O�[�Cb�t��W��:x6a�A�}t��������~�}�{��9G� |����{Z�^5����P5���,�.�I~���B�7�+���<M�πV��̀&�L��
k@�k݊�i���`K����_b�Ga��֋�(��t���������%��t1Y�"�qaZ6i�Ȑ�B� R��Ս~I�7ࢥwnݥ��?���'o�	 24���
���������}:=9��wn�O�z�w��<�B<cy>�!�L2Zͭ +u��D{�+<yf@�{�r6V�>e����|4nI۵̺�%|�l�fW\|o�<�50�p���<��]c�S
y[���-5�wȍ���_F���� ;d&T��\|C;hd%Oħ���x�/��X�7��C�����K���4N==�����U��X�
R�>x!�����ݿJ{�{t|6��ܥ�~�:��ӟ��8l��;B��>�qˉ���vև��S7��ߥ��S*ú,�A�͖����Q�� i����iN��XV�,�T�%�c�\y�BT��.��E��V�eڥ ����a���K��g�a��ߢ_�>��dJ�J*�g�k8hy`U֍h�2ƥ�1;u�����N�@-��Ր��e�4N�.��w'�?�� @�Y���X��J��~�a�$b�tI�,(j'�lIgc!m�&�1\ߠ�
ֵ�E}ԚR����.T�~��h�V��b�=ߏ�.�(d�9�����MRP��Ό���:��ȭV
��~W�k�Xh�Nk�*nZ~ z2|��QL��'	`�y�i|�ݰ�kD����H��ʙk��+} >f�]46��QC�Ի����)��v����	W�����'���-��!�ze�>����c�x�.�\b��<����^�:���}����O�����{��=g�	�m?~U5aBC�5Z�P��x��}�1�_��Ч>�<}�o�K��o/��{A�����C�.���Y��q���֯�(m��8V�ظD0.V�	xƜ5^f&��U������|������g���Z�w��
�����;'�����c*+���YF�0<@;�ww�é�D�8d�+D�h��c��R�g��L)Td�a%�\�=:�!v��W�Χ���5<�T$�f����rnL�ձ�'��\9�B�*��>A2��J�qje��|���8>�}����d")zo��̠��$ã��y����V��GjM�'�ȩ �u��O炇�(�j_���������t��{�ߓ��8�k���L���]6�)���f�����K�V<g ���v��km_�*��M� �������x9�;�ܣw�D��F�aC �5]��ބ����ӏ_�)��3�-��9�Afe�����4���$�~��M_��hwsD��6�vJ��������6 /KQC/q���Ş	�KX$����
0�4���亼z�b@���MM̼�����Stus�N�@��:}�����u�?9fIEn �
8�)}	�Ű"J���P��O$-XA�%��N������b\/٘6�5�hˀ���%�:�j�R����(`!�΃�N[H#�n;�5 ���SM�o��ɂ�J�1��e�,K���Nj����X�^)�}� �&bZ��ةa �B��'t~>K4f�H����y�,��<L.�d�A�f��y��ǅ������Xp�Fk~t���g�#�������q�/�H��t]銈�H�!)OD�~�V��+�J�Q�PR��՘4$��K���;�V� ZL�����V�9*G{�4>����.j:;�-~wt��O��6�]�P4"I�� �gL��|�zC�P�����C��ޢO~���7ޠ����.��7Y�⠒�q�RƁ�8��(HD6f�i~uYNn+����Z,x��s��.S�#�v�������=�7�,��	����!���?7��ExE�מW&�����e?xb�f�Sj#.�����"�+��f|��{�i^3��x�$O���[��:9��ـ�_i˲tU!��_0w�"��M�\�S{��e���q�_��x&��Re�)��U���d��i��p�X������jhd������'l��b����\���D S�@- V���W�)�B5�L�m��" ��kO��Ġ�p���9V�)������)��,����c�c[J)�!8�Y�p��z@�j���^׈LZޯ�8�04�8��QiM���~��u:��Կ��ަ�0��r�@#�+FՐ��\j�194V�����qE���lZ(Ѵ!<���9u*��e�s��Y�Jxe$K��	��.�"�x9��L��hn>�B+*��7 �z;�
iƙ��l�_��M$�z\�ɶ0���g�;�Y�^x�#N��P�ѫ�D1�õ�i�BЮ��1��q��e[ѢvxK��i��E�_6�K�
w�%6�U�<����������D9��qa��撚+�7j�Ե��5��I�>k�e^�` ���t�@\%��1>HYZ��!��=�;hb�P�Ŋku7�F���Xm�3��^x�M��9�}�F��N�<(=���	ج�;����<��Ec8��l���D�%z��XE��1/f5#�/�Ƈ��XY��2l^��F!�8��X�(4�ޡ�S��a�ͦ�UFk[����^
��ŌF��!"�EdƭR\�E�4�}_�R��ڳ��q��q82I���ڐz�Snč��-
-h��W��G�gR����}���<>>����`PwWG�a��*�cCѐ����l�͌
m�\�\GK��dC��'nyc6>�u�(��Է�
]�>����q�L����"Y-cb6E.H0&��l�	6#���&@LRI #�XO<�B�mx(x=����&n�Bó�LD��Ȉ�C��Ƃ�a�pGZD@��GVƗ~��QUm���]\+��$0�V�l�V���2��^�9ƵjX|���-J
t&%64Nc�������}�̥d�Fa�p:�\�N�=����
���W+}�̬9/���m�-r�L�/k�8�����n��߿G�Gt�ޘ�y�>�X%}��RZHZ��h��Ҩ�b)�k�'����ݿ/\��VF�F�#�&��uBO1�,��^���b�O���Cf@�]؇qV<	�J���n~d]F�[�iXLT-^��3�J�t��&��XO�h�&�'��B�hg�</�v��F��t�nޤ9���ӱk3����]3o��_D/nu�3\,c���s�<�[y���;)������R�G<r����=���@M�����8�Cs����Z��a����?��$�fYJ ^���I�;t�҈>������]σWR��ҍ���yƪ��MD��i��K��p�����{�o��S	m�52�!�x��t����ݦ���g�:5��0Z�UQ,K��5LR=[� nݚ�t�������y���X���d3�V���bѢ<����\llS���?�#����-k�������N(�m��xR�N�^�t����'�1��=lxi[�%�[��ad&ґ�5���]iY�Z �e2r�$��OF�/���ϸ&�M���D:��<՝���4�)�ᾸY�Z��Dʾ�M[��ĀY��E�U���~�wz.|�#�Pq~Wo�m�b8��,-i�f�����:ŧP1<!F��4��҃`*0=枻.]��8]��t�fttzD��^jd.�k�a^���U�V�����r��y��h��m5`\ *8E���p�C�S�dXj���Ȳ��x�����e��ᦅ�����Gx=�����N�#
�|fD����&vb%�v�[�K��鴌g���0�L�!6I�)�E1���c��999��2)����\R7$�1Mܰ�B&��2����/���#�yq���c!�t�T����FGF�/)a���,^ �\��B4k�M���+V��.z"���@51����Iް�
�����8��G=�џ��0��j1��H$Of�U�F^[�]2�|9���V"���P���b�خ��:��@&;�T��s���c�%xt�������
��7�w5`ή��pr!%�>a���(�_`�)X�Yb�����Tc�k�Pu�$ÖN��F���&$lO�6"� ��P����pq}t��%f�E�PÑx�Cp�&�,�	�s.�ᤧ'���x���X��>�A�!Z��|ߴ�� M�	wnnlr��`��ftR\l�ㄬKz��QȽ��~e#Y�E��n�^�II,6.�ů��D��&����	����.����i���m�q3#W�+���]��,�m�Q����F�$����"�k(�>.>ge�u�Rv�ɘ�;d���.�8��7������s�	�l����r��6�YD��&k�l�kg������h��P	�iUG�JYЛ+pk��@^kT�Ʋx�= ��W,f�^��(��G��f���������#} ��ߑ�Z���]���ƽ����͜e���&�(bP<--�X/sI@�0�Εj|L�+Y�8IN3%�5Y'y�`q���������� ���e����b�|��g���UAtk]�:�>��- �\�ăm�ż�R�<!��x8�b`�͗��	�C@�*����u��9fK�m�w+���K2Jјz�"(3R&�$؊q���0-��q�)�撱Lr��tx��TP�Z��܃ }��f�����ɚ�uw�v��|ڮ9��)�qJ$�`�e�f��`�Lk��������so&	2?������%*y�t��v��2@*j�������`��lQ3k{�	蛴Œ�� ��&c�T@Eh��s��bX��n�=<����3I��,�wT2��ի�f[B�3�z$�
s Oq�,��Q��e�����a���9�C��^�,0�����G�K�Iо37Q���z<������`���>�ǐ���pET�Q��	j� �>m��Vx�y'1TP���Qٔ	�M(�w�Ng�@�sʯ'��V�6��6��I��c �U�pխ�Q��y�_7a�J�Z�?��<t~4� ��¦�Ùw�/Y������>��8�AV�ߒ�!�g�f��|��]Ht��t���L k�|�6[�O�O���}Z��D1pj���K;�K�[�X��	���u���Z(ч7�D1�,�>��`�1|:3���'4Fk�:`!f��:��`��$�8Ÿ�zo�`�*x~�X�sQ��,$8#h U�!z
_k���[�a`z�rU�pF,[��gT�B�~ED�����W3-�<�R;�\��c��!��geՈe8E���O,c��p�>��L�H]��4l�,����ݸ�A1r�`���D��ނ�$ѣ�C�kW��"N���/44qErJ��Fu<M�D��e��_�}��3Y��ʇ�yA>���2��X#��y<�����V�{�cQ�گzɞ6T�DHpC��M�E��	�[�?`u:����6�D�|X�&s��]�L�JJl�ӢY"�h��?��]p���gg�!,	F���C�!���9gR` ��`}��ȉ�(ɄIk�J$m��4���xp����K/"4�'��1���Ԃ����8����lA<����Ur�`�6ܳ��O�@	+Z>�aA	Pj�Ҽ���m�у��}_h_���r��C�B)yS�/mf0\�ތa`�4��z��kdMXk���_yL��7�Y��騘�b.y`י��^4ZYh��Ϸ��p���ȼ���!�,+���U��}"�p2omm1q�e-` �bֺE(3���{4Z�!qhr(�ƇQ+�h w�dx`�F�O\�����qCH�v.k!<���l:��w>���wY��k�{Uy <�F��!%��e$����&�ts�3?r�YH���(��e� �������/p�A	�����#w}�����p��L�а�_uY8�l|K�2�li��.���.����K�I��<��$f�G=�aj�O�F����S\=��q)��wEd��7zNi`������E�(y��=�I��hOm�yx�������}DH�ꚱ�2�������{קy"��J-���qT5SʇaC�D�C��K��wz��Dj��~��}Z�Q�ӏ%
&̍zttțt�W�ΗrU�xa���t:�%!Hz���������M��N8�׸3Bd��f��ŵ��sq�\ؼ�}*������;���z�pTx��;�E�=���ǰ� UGgis��#i^�/և=�yp�?*N'.�_Մ��Pܦh{�S��p���8�(�#�4'|$�PKyg#�r.�e)Ӈ=���*V�^�
��j�6�y�ހ��tɫ��:{����y �����̓�R��r9�>ǌ�}6�e3Ut�3����O6N)���@��/�|cV������oL0Y�0���&����	��4x�3�
�!		�L�,��z���m��?أ��6G��������!������"L��9��1�u;�� �/��s�{�ƍ�����^	sT�.�^%��TN>O�N ��4y�?[���@mߢ�I�$�x"�֨v�Z�Zྸ�ĲjG�� �M��	�� �l����b�0r�U��N���ՔvM��D�]Q9�3����6��@�ч�F/�ï,��$���"@�ՋIx�.��)T���Ix�5��%��#T�8.K�,����8�е;��ga�o�&��K!����dg�ov���,�~J�f��V����Z5�N�.�}��Fx�Э�uC&��7���͜L���"af�]���+b�g�R�u����8и�l�(-h��$�w�B=_�|I���/,]n���ݵ~��1UM8h]?��w���A٩��^U�������/�:3R��������'�wz6E�B6i)d��܇��j�m9�J���A0��!�`��^�B���"9Q��[�
��؋�FLJ�;b�ns�2��C�l���s�,�t,�S���FiU/B$Uk�B�2����C�8g�Rh�����k�,IU�+�Q�sZ6n�{���{�y�+��|�Vx��nq���F���L�m�i�Ni�S
ջHi�G.׀�CdU�w��H��Z�1�.P�[x�aʨ��`'y+�R ']��ȃ���S\:�i#8m���pG���� ���$�q��}�_��.�,��q��ɫ���D%4DP��͗Q��k�=�_��d��sU�BVkA�`D;"4���%�B�M�͜�T�Sqx��TɆ8���o���j��<��W�r r �����k���*>��N��>�B�r��C>��4���}��AH�u�oi���*b��~�e`�Tހ�9�,����A��p^ٺB�!�1����W�����ŏ�@g�gtit�N.ݧ����˅h���1_lx����� ���l��^xt{%gX�7�'�2<;�#���`��K�y�Z�Pf|&�
�)�ct,�.�L8GpL����7�
�nYKV�,�z'M��a_t�� ����6Z�k72V�μ��ŇՅ�S�OY"ߚ-�	����Z<�W].���MW\O_���WPˢ���������I,���
�@���Y
��ZQIQ��^�ȹ�`r��E}oDō�h$es}��V��=o�!N��ȧ��n1y�|�`\+Nc�&Fc8�3C���^���sY�z���/��E	=�P���!��M��x,�K}%,M��l@<�f5b0�!�N��̟�G�[�?�K]�j+��!�w���cv齤�!���g����vĒ�v;�5'�p!�W+>(�d>l�s:8:�J�^o�iY>p˖Ō��/M}^������M뿌.s�l4��0ce�貱XF���s�t��ɢ�3�h�Y�!�T���
��V��l�4�+�����&ɁXT���P�>��$�>���׍�Te�mE����|2����Z���4還��6�n5M��;p�,��q()	-s#���-���X�U�r巵Јs��-�宥��藠�G#�[	��+��ٚ8�-�b�t8�Y�d�N��ˆitaz�̋���]4�v���H;�2!��C"���s�+�R���}����1���Ma���C<��B<G��T<HzBkf�mT�߫2����ۃ2	�u��SHK�56օ����K\��
�ŭhع�N����X]zx�K�$��l����D��|��;Ⱥ����#&�?��*M�^)s�@���ݢX��1�C�(��Y���[�s�ӚC
x.k��?�v���`bv��σ��`�|G^Wϩ��2���#��FXl�Vď\��= �)�V��d5q�"_�Ǚw�И+�]�L�K���Lc�5�W%����b���#e�m��`!��%c�@��8W��Ӹ^��4n����3g:�h��d^+g;�~i3*n|��YM���������l��P���j1u���Dúr��{�ݗ��.d���+��SZ+����S�G���к��0�GLÊ���s�ƛz]��何p�E��ß�z]P�,#���+ס!�yi}��B�gRYE��B�di\����ߛ����G���S�t�u��g'�Z{5N�YK�4l��%w���d>z!��Y[�Ǯ?N�;;4?�q��T�����ܹâBhI���[t�`��]�F�.����enu�d�U�Ё�P)�5Rx���h<�Ss:cc�a�|�=��A�>A�ذ`��u�h9k�B�z2���L�,:р�}j�/�'i�Q�$P�qX5"$'��	4l1�~qY|w@��S�}�Y��YH�-إ�x>� 6�Ʀ+{$�4�R��[)�����^��u/އy@֌8�G�n�/9_�d٪���3�{����4s���`��M&Ѱ
K^�.)�@�6�_���FF\l1��\�%������ ��aq�F=�} �o��`l�4头=]��+�D�M���4�|*�n�9��`�"���x�-���AX��bS�"޿xd�ȺY�V��0�M粣��<kp��}/�Wi1aqT�J�Z�ҙmv(xm� a��G�I3�d�g��L��H��$Z�����U�'�c�y�&���7x�^�J/��}�ӟb��?9���c4�1��kpS�̘��i���OOؓ�z�J�B����yC߹w�����#�A\��NM�اJoQ�o�t��,W[5\��,#U>��5=���BY%��؉s�X����r��Nú��b9�tL�+-o5,p��ÍQv�hV�=��"g��Nq#�o�7#�-]Tice=c��գ/rZm�M^Ō���Yu���5RN�@Ā,����Y(H��4*y��s��t��゚�x	Q���q���Bj,��	��4��P����m�S�����4$F� %��+;k�k?G�",]�YWp��M���UZD�E�z�R���Y�7��[�V��H�hS��|���<Ѱ���YH�>l~��P������ �(�/σa�0���u�ф+���<g�����=��S���G��ݢ�k8;;b<���px?��uꆃ|2��7��BLz�X�e����0�.���[����9�<>�r��|�k�+���U�zY$52^�u�yܐ��%�ƈ��F=�5L�Oi'x^xD#Ou�Z,%Efw���C:7h:����Zݨ��t����J��Q>3O�Y8�(�u�H'�B���dR�uk�q�c�i�?QЖ�BL�d���xǲX��i}�^��6@����9J62kYoE��Vj�
ߪAl�$�6�I��A��B,;�1 �C�
�2\�h�f�$��0پ^D/P������V�n������M�|��E)I.��՝���.�h�$x��ސ�y�%�[�$Ռi��Eg���I����M� Y�7f�\�;�U<ə�j_1܆�EO����#���١�`�g!ʅu�ڹ��!zͶ�P��v�k������ƈ���/'���`Q��׷�(2E}��::<b����m�F����h��s?��X�����v��C��Z���h-�:����&����f-دU���ŀ�X�:��x1��=�"A��LB��iIȝ�K�F��w�#ΆV��Q��t�"����*��V";�y��t���pm���;�6(��ܿ���g�֓O].n���ԍ-x��F6(NQMA/XL �%K���&|�w8U�r��ױ��Pu�x����ђ� �=#�k��*;ᱠB�	�U����ެw����\S^|�g�H4A#�ex�
Q�g�����F�K�p���4�mr���I!�*��C��a��Tl�����fa6�V�V�ד>20�hA�.kv�L�K�F`8N��8'ooN<F��� c��8کCC%5%�P2 k�����
g1�ر�x
oV��{_��mY��j�&�Β���b�	���U�(��5&$F��)�w��?lM6�=tk숱j�@+�m� �WZ�.lomq��:�!�]��B�w�ݣ��㎸�k�/ѥ����}o\���FQJ����!�=���X��v2���^O�zG��v�����ǞE��v��*@:?Wwe��NE�A��Dl������";�6�b�
���w+m����G����d�"�V��W��4(Nc��b 9���z�jZq�&ϭ��t��f�X3�uJ�/1n����5[�	>{&�e.�\s��U�5]����gAwF:�Rp��p��}m�.@8������7-ãV���#{�Ʒ�g��",�W�rWv/�MޕjNl���z����iQc�������eW9�[mm���d�wP���§>N�[�\��5���y��]z���4���y0�%L�(���iCd�r�+��lv����,c�Z짦!O���Kz��>�c.�4�[�L�c�Ț՛72>�o�`<���f@�jx6������w�3��º \Хݝ]	��G�ةt떼���G'p��	�p8��ϸf	*|���t�]0=(�a��R!�5Z=�N#��v>^�%�O������}�Wu"����d�J��%���e��	40�e��b �5��\a�l��2:�9�:��٥^�Z(I���a����k�D�ӭ ���>�O}��Ͻțfm�����{���z���b��Kȷ��j��(19���߂c�'�����>��[�8Ƥ�'��{�e�woO�4��U1��$��n̈́&(^�5]�X���_���k���k�)phF�޺�>���9��ޗ~��� ��{ �_kK	&(� �ʋf&H�/|�c����.]�r���#���T���ŷ��K�LB��a�ͬ؈��H�+�"Î9����Ԉ�D�U�:�t��+'Ƥ�l�����)Aۏ^^���J{�9Jjg�p�0tV��cM���:���gYΖ�5Ɂ��m)ռa��� ���xI���L�$l�G�@z8�8���#$�-�L�X�� 7�0pD�!��H}������<;&y�����tD}ǒf�W���\9�Ԁh�5�-�
Ǭ$�,�y%rxf��w<zIt-�D��K/���h9�h6�E4Um��|\]��n1H�h��B���售<6���>}��O����/=�ċs�;��ɔ ��0�@�q��lD/�#���ǀ:��������/|������Xn)[L����>ݼs@w���(�ā�U0V�Z�fm�`|3����hcs3�ǝ�%|�����G�p2��p�{���ݡ�n@�޻t�������k-Op�(�Τ��Z����~I_��o�Ͽ$!b���!��k��/����?�{go3>���D��*���a�q}HVL@s�7!���2f����G\�<���ӥ��a^ȯ��g��j�/c0�B�u
�����Ax0
��41�x8X��U����\u�M͆��1qu��O�Ym@V6��H#�p��$vk�Ttü�gՑb@�0t�sh`�ǲ�'�
��z�(���pâ���X�]ڠ�G�����F-�x)yf�a�`q����ד�k)Ʋ�C�i|�3��S<A|��{��Y�-Y|rB�kn/���r,�/�4�_H�O�S����g���^���<��n-����KW�ُ}��x�f8u��'��3��r�i �zhְ���7�_����ݥ��!g&p"]��7��U���oҽ��`�p�=�{�֤:�kG p���'POt����3�}�
�w�6{!�&6.��'>��?i��1Z@�89,��_2�.�5b@�H�k��]6�U0�<��`4Ft*��uL��O�0n�'�y�~~s�N'5��D�D�*R�#�'H�[7y���wH�����^|^F��k���6}����>q5�I�b��+2cB�x�i���������1����3G�R��JI�����³�K�N\��I���a���u��s���������]��ǯ&����3���O��LψG�%2WlĐf�ZA��~u�tO�Gg��8����ġP�x"����N(n��
�aRJ�Y	��C�N���G�a?�a�W�6C����]��������s+N׭fj`P)`�.|-톍v㙧Y�rb��+*�`4���s�͝�����K��{\VWـ�u�ai^�c�p�;ۛ��O}�n�x���O����}9�B�jB��K��{5\K����RZ'�z*�H1y��)IxO��W���'������ZL�c�� f��)Bس>�(��p���	#�H�x�bBcAM������?IO����)ZR0BU��j`9������j��[;4�O�o�x"��j]`��(5d-R�b���7_ܾi�z= V9G�#Id�D�2㑆Iן7z��g>�-�+ˑ]A���h�RΌ�	�z�`#^���OYX,ز��^BA�� ���� �����l�|x��;!�Y!�J�k��X�8���]�>�Z:�K=���:?;c��z���-Seur�}���EUO|Wq�IbL`
x���N���ZlaJ��ӫ�v��ha�9�.�(5Y��̵�۪��#��uz3�4�?F�ak�#l��t���aPr��%:>9��a��l<����8��ai��<.��Ҳ ��$dm��섗�����;��?<9jr8)N��b��<x�*t��8�|B, �Y�kW.ӵ�W��pʅU�'�tVMx�'�s.�;<8�۷���<Ľ!Li�P�i4�V��g-�r�x�}�_���	��ݻwdFJ� �������F��4GS�	Wv�\�VJ��CmYA�&'�F;y��婍���f6��y�7|~@��b�G5<�-���t�˒������(�{1z&��Mʰ^���"#���I��x2��.��Y���޹����K��SO�lOxh�H��:�8l���5�!M�5ݖ3]�z��2�h�ɭ{���Ʀ�VJ�o��������I�<�Uh��zݞt
�9>9�~��� �̧y�q� �ax��K�+��nU�~�R;S�D"�4N!�D���h�ӡ��%*Y��hn�\��[QO���������jZH�����"���w���)����v |P�2�#�%��O�N��~�}|�-�
��5���W`�ᯋ���f[�/��������pY�|~&�J~.���Ox���� ��lrNǇ\�'l���i��H���F@K��X�����`\j�Qg��=��"�B(�ςS�p��.͎Ap3�yY����2��͝�fC�3\goƴ�Y&T`��B+���q�^GB0"��z��}��ޡ���्ym ��b��S�8���n�����t��>{"��[(��i�Mv��S{��Nҭq��i8J|���z��ͮ�H)�ZH�%�9�~D���k��TY�F��UXSH�b,v�{4	�_��~2�K�!y��t<n�'P�������B�'��Y��+����٦�=�|8|.�YX3���:-xU<��<�{����:g�C�+�AG�F�����c�uZ[�5��,�;T�^�|9�հ�¡@�Q�	aƚ`�P/U
�ǐ���F/bࣽJHƭ����9�����+�C���Cx��s�GB����T��<��̌�C.v�g�%4J
�*V�Z��61F��b��K�(?z�Ċ�Pad���Il�^%'��۷Y�a{s�]��|Ɔ��p�G�!�=
�@pC|y���0������p,m�%K#ԢC�����������O}�]�(��I ��0�g���Y���3Q�F+���o�H�2'����o��^������p�A���΋48+��R�֋R��\��wYJwn@o����O� �n(Nd��0M�p��m�E���00��f�i�(���|�r�ë�<�RG��������@��l��@��[s�+%�9]}6b
H���5�qR�M�^�4^T\W�Hp�$�,C8<�)0�VtZ�� @��$����.���P�)dQg��X�z��MS}z�����n��)���r�O�Ť��WW�,p��^A����ާ�)ntoU�N<3���
O�wx͚: �5�Ue�G#b�_�(,�N%e���v��j���w&���������Z�N
8�9�'k!)��گ�H���'`��G�hHp�"��9���ۜ��N
ǥ$�7�u
!ܰ���w�_��_��Z��^�����9A��7Z_#�֦Sʜ��>fC3�34h��%����g��v�\ڢ��-��0�È;<�B���ɐ=Bc�I����}n�����D"�8���	m*��yçh��0�hC��$<��=:��^aN��@��gx�E�O�忉Q�X_��41θo`S5���-l�(�w��VY����>>�$<���6Z&�9>�>�"�#��w�y��J(?'�!T0Шj��'�Y�c+�aN��N��/��y���,�r�{�QZl��<Ud0su�C꜅9�"�:�i�h`kc���!���Bgd���&�t��ƕl�A��]�h�fൎC�	!I��	���Y��~�%�#�q,�GM�o�XI�Z�{��p�_O>�����	���j�#/m�t�Q�\�IE�M���(��K&�'�zrRC&S���'����vu�>?��~6ǂ	;�q8�������v0
ga������usk�&����&@uG`29����u��{��?����Բp�	��;���f��U�^����a،��@1�`��ސ�@=?�ܰ�aH�޽�c�`l�l��Ù:�X'!�D����DO�p���ޥjH�|�>��0�I�4�y�滌�Ԫʛ͓R6���T6�ڬ���Tw��F��ѣ�QQ�r��h$\^Bqq!�"�K�y\�#����O>z++/�O+���{I��O2��k,גU��e���_٢��o�[o���\zՐKEm��nl�[����C���Y0@�q���yl$�Z�ʕz��g��ڤw�A��gg�Nng@�'u�jN��ru/�ң�*��=�ӥ��%SpADd��_6H��E����~��\�D6�����W�O�VZҘ�x�F��Z�eY(.�h�X�Y�)��B�I���I��Q���#�>| Mp�
@&��
ܡ+�V�B����o�g�7N��l��c<9e�0	�=��;���72Fh�4`l Ђ�V�����y�^�˗vY�ʝ�I�Q-a̽;���`3�S[�(mm�p����@��C�G�a/����]q�\;N����Y��	��	�����Cv|t��u��뜪���<xX�w3
S�c�p��a�Hq�~�6���ۼ`��`��� ]�(�/R�8�J������渿l&�!B���R��51�C����h��ўۇZ@w+�aw�i8�.|��k�|KU�~��8���*a��F#6�U+���NK�=���������0F��qI�~G�I�ؠ+��bT�XO�8���aL�����%���$�?J�zJgcVͲ�瞼�Ͱ ��Y�qXS��G�m�úA����AX{��1�n�1��џFE�:�Jm!m"@�i��Z�
4R��
<V���Q�S��X&C�૗P���J�}d�#)��sʛ�,�dY�Q��%�P��(?d��!9�iZ+U/��f>;;`�&^����� �Y��r��z��l�cׯ�M~�C!&����i=l�ɬ�m?'�y�;�aC�T�6���DȰ��&M����)����' �_ �}4/ڸDG�P���	���+t��j:�z�]^O<�K;;۱D�䤠�;�<�0
�>�TX�O�f�>����R�	�)���&���e�cZ�]���MV2GM�����nT[c���]��F��d@��5�a��E0)�i�#o�AC��*qy�-�/".�ߡMp�3���e<%�
�"Vn��-��q����NC�z��Q0�_��/�Gǽ����y�"]8z��"�����`0�L��F�|�Z�ٱ���0,0Ͽ�,��x=���,8���&;OZ?��	z�̚9�\XU�b�\僫��cb;���Ջ���q0葙�3bI�9�X�2�ԋ�f�:����hHr�Vؓ77�9-(��t�²����D�B2v*E㖓����'�M�lɎ�8�y�[��  ��(���,�L��/-��/����˟$yٴ$��H�E���F7��~�T��;ߛy{G�̬ׯ�����U]������9qvD������O�xOX�ei�D���.E[��O������x�.�}�����$�u�Ԫ#%{i�@�kj����t.����{�  ��IDAT
����&�+�Rx�ɼp�����@�$�}�� @�������ʺ��-^�]�ׄ����`�2ML2Z���|a8d׻_}�t��@��t��5YN����#��X�L����c��Q�x$]�LHè"&��o�um1�r�]�&��=���&|&�@�BI��
v�C�n��m<cHDB�0����A��5�m_�9Hx��$��s�J�W�AkV� &J���څj�X>�$1V���s�z'��&�P�
Y���'}�(3� �~¦pB��@$٪�d1�Ө  ���<�]Arf��Xԥ�|RT��(Mw��u�Q�x���資1wEN���-�E�h��	U������q�u��}z*3��M~�18��,�g�ڴb|��uro��s�y�VnoA7��L���2V�R���p�c��@�i��G��N���n����A	[���H����t]?I�%� 34�}cJ��YE�r���1�3.8f���B�_�.�n�b�SR��8pGn�~Cn<�)~��� �,���o�S�P;��-8%@(X��LOMF"<_���d��w��0�D���޸ Ǉ'r���F�������A{b��"59@��t���c��q':I�(_}�]y�cv|r�;TO�䘋\=u�ཏd5�x>,(�Z 5ٮ'���9&����K�/q,N����]�][[��?��~��e+�ӏA��˲�u1��^ɨ|m�|</�A��+Y���D�'�8�@��!�y�׏,I�\�Ʋ�i!v��q�(���]E�a�bf�wH�B�������;�+��M���)7�%�X�qO:��(�+�ؘ��B6a�{y=:���&7Ӑ�[[R+���G3p�����t2.f$��+Ĺ�H��;�y�n�RǮn\�ء��d�Z�\��q\>��������㩢�dMu^\�[ϯn���X��^6�d��*)�k-��:���2UN�|���jظ�,�$�h𞇯�������1��cUO��>��1m��\T��,�XАp�*Rc�4E0t,�Vd(+k�����k��+�|E��}N�D�D@������PZ͏��6:(䤽���r��O�{t|H�k��`�՟�/[�m5d7dW��3[�C����;��Q�f��x/��磌q��UF��G��/�ru��u9|x��ED��R��j3���w�Ɍ�`�ˋp��qD);�=4-0���`<��������=�CAw�Aƪ�@k����"�vyS�K�]�a�h���}����We�f�����_�����Ƒ�Ǩ�n��c�@*}h)T�u�-6;p4c�w
�Q�]?{xx*����/�P]�o~��뱚BGŐCIV�3f��:a��B�VEs}6]5H����%�CʰB0��ۀ���y�U�X.�m��.�����rs��d����s�ȣO�Kr�R������M/����K���"���':�{a2b]��tx��<T�B0Kd7�uL�~�[a�Ĵ3�>yJ�BD�t5M���eX7~k��ɱ|ūQsvl�<��Ie�+7xJ^Ji�1J*��?���`��c��̚��R�w�CP�(\bE*�^�;"����hDD��;���Ů����ɄM�����1�
�E��M�[�j�n޼�ڇ��ǡP�����5����,�R����br��������[�Q#�,
v�^� ó!Q)��b"�(g�h��K�^z�`t{ ���枀�$���:�!g�Κ��!4�Ƙ����y�
59�i�D��":�I�"/~�Y��7F��͍M���V�c�@�b�@�O�� �/'����Lo*%��揕�D.����������/հi4@$�4g��"Ml�iLal0�����XY���.�2{��aѢ�D/tû8ږ�4ѧz�R;f����#����Y�麅;��.�" ��M"#����{6��6�N
�Sq�jy���2eA`DHըU�Z-#j�5|0\d�R��h��{�Y	�/.�豕���!�Ey��93���b�xOU��'�&I��c�2@�nr|���ӭ��HDSX:��t�9��㉌G;��3b<�֚7g����ʐ	bv&>DD���f�lp_������J��ڜNҪ\l��C���d��(ȓ�	��ҩNBCL*�t6l���Y�y�k��1�E�߁ሞ;&�;���s���1&2�\Y����[�P�/��d���d:׉��40Ί�;{04s��O����+���U�>�(e��cHc�H�u[s��({f��.Ȣ�1�o2G���aD����Èx�P�q���Cy��>ӝ@���f�L~S��Mn](�*�1�:��8������[*��0g6�ϲS�npC�=-V2��S��{GK�F9�H��(R��+ɷ��S��ydn
������Gc��'�enD`����گڈ$��j�ZCJ]#b�`	ɂ`�3W�ܭ�_+Ew��G�,��U7�����t�|��w��l}��@h���
e����3�����(J��v��}h_>�O;�.��K���Ng3<�H����m�Pb�P�M��C/9'��a6Z���x��HmN�eĭ�g�u7
��0b#�,Ҭ�
��;V�؆�.2]d�P����A@5f�H� ����8tE"TA�$vQ0PQٌ��:����9y,�3]u	��Ј�HC"���C�4�dK��^���n��R/9/*��H�5�I|*P��璲X3	��PNRI�"ba��!x�F<�2eaihb7��)�[-!ͭ���[ ���V��2ǁ�o�"�.$�͢Ϗ���p�	���6�x��
=6â0��\��j��u�z�k�ش�s�  �b㽑�� 7Y�����z5�4�N/�t�[�<D#�aͳ�74���k��(Qz�?h�f�5�7o�K�jWO[���1&�Dj
i�|��nnu�%0#�I�q��GS���� ���08���8U?nV�^oi2c�^�x�Tv�R^4T�}�I�����:ֿ�ĳ��.���S�a�y�n@�������� ���d2k<��r�n�z�0�1�D)�H4
���E+�C6`-<t��١+�ӟ��w�}��<=|J>	P��������i^g����ﱣ.��r��A��n��kj;%�F� F���˲�]��jl�==��֑-���U�&���7����r)|q'#�6:��5,M�1"sj=�l7e��=X*
5E�I���D(����-].&�YT��p�0�`"�H��}��M�`f.:!�P�.�ը@�
�C�)����>"j���YFMX���fF�3��l^�
J�c!v�Z�����bkh&KH��~2C�4pV5l�*�9T Vb|�vB0�6�������s�jc��_q��M����-nV�Z�?������F")���j9<IY��X�;LI[U+O���]��Ԟ�u7m�����ӕ���x 7�_�d9QT�֙���
��C��@�N��Hݛ;w�Ł�
k�,i�aDP��EW��;���@}���!ks��M]dV��pz���l�Y� D�����{|,���ӹm�W�2^#�����y �>D�VԵ����ӧj(,���}����l%�E&��<>�GOO���T,u�";����/t��
��(�h0��W/_�5(���͈)���}5�=<��z��i��wJ�:�[Q[��Q�?ߘ�Q%m6���.p�����Ew��@>=�#y[Hl�!+�x�S4�/7�z�Qwa&�V��������x�q΅�1��a���1Z�u��C4W�T#]d&lM��o�H��B��N:�@m@>�iV�PU�x�Y6���"#31��q:��l��������Z�<�qG�����Z�T�����UM�E[��0Z���:ee���F���f�(�g�U��Qa��f<�ں�f��]��~`	�����\���Y݀ʅ���	I��M9��k� �`c��ѽ�.�:�Y����zm=9��������ﾡ0v&���S3;ׅt"S��oݐw�����'��3{:���<���]ϕ{wu�ZA���W����D�^�aW��X������Iԣ��[�m�ۺ/}�����{r�H݆� "UY ����������Rd��ݕ+��}S'���ۏ�PQ�[o��_o��辜�K��GS��G+2������.�Mi�:� F���@�l�Aؖw��\�q��D�3�N4,4�ٖ�+��G?�7r��m);cNtT 봵��#�"�M��&�&��Jj��8�i#i�$�,�+-�)Je,�+���`s�Fec�Z2GA�BU������f@؛��Z�<>e�x�tj!Č�b�)�`
�cI�%dif��l���7��B�~Y����-��ơ)��:�Jyt�q(T��fz�9,Z��
1?}vV��9��P�4{d��a3t̕VD�\?b�n�V�*^m��ryʬ%~O�0b���˵=ki�x[��V%o���%ݑ�6�E���r�^mznd]R�Sl@�������'g�Δ�:?���A1�M鱒��.(*M���������޿-���eY���3�4R���h]��{w�ѣ;�'�Wx�]jl����j\�]��s㒼�����d���$�ܽ-�aW~��U�y�5�S����19$p�6PT��f.��!(�\�OE�׌��ڵ���͛r��E��|O>���2��'5�֭�j`����/�������~0"45=)��\�*JlPs:{��7��wޒ7޼�������@�a��o|�;l�4ީ��_~HR���&��҄�S�D�������ب�sm�� /���ߡ�����YFL�٥.�J��t����	l�3�6p�vd�o�[L&���ř.��͌�Lƙ9������r�����}a��"�A/^E�8?٨�HtMͷ�ͻ�*�����#��MŘ���F��1]h�� ���)y�u��i͵1p���Ԁ�7��l��5H$6���P�*Č���{����vӮbͫ�y��3��Hc���nԞP��q�
�n�d�܃��c�����)]0�)�Q���ʾN�.!���@^�yE>���٣��
;��p5.]�_6������ݼ~M�%u+f��?�X���9<��б�鐩�U��x'�jx����(Z���$���W���=�կ�ݾ\�~A��ծtF{򉢆����nwK��3JPO�+V$��7,B P�o�!��η�ʕr��O�����������vGN�����%�wuq�!�oث�,��\��+�<S����҂�+[&$4�=�b�T�\Ij�`4r����Y��Q�b���A��dE��.�x۴]I�z�Y�P��e)iiO�<n�~�O�����1�@�]��ݼ^�\ܕ�S�:��L��it0ǡ����CY��+��J�'��ڸ
7��X[�����v�����Ǎ�s���3. ��C�a�r���bڠ/{5rrM\,ԍ�Bm�ڥ�fL^�k��AI�D���[k�F��H�!����O:��5�>@'e�.�Y�p'�j.�_����U�~�3�����}����W��$ 8;SX����-TY�&���=y,7՘l����G#D�ՠ �pL*��\&41�h�V\ۅ�����7IX�w���w�m@
e��jn�>�f�O�N�������l�7�%�Xf����������;k~�𮢞+���7���n�w1a�^z��Z��}P�)E�F6ZZ0�g&k"�g�NH���k69�i��s����1�S�M�"�Y�:�����q��7fH�we�O�`3�)���I��D]^5K�C����d����v��{l���@���My]M�Bn�b^[ ٴ^�ñL܈����=r������Hɔ���Ϭ@�(�m&��^̈8Q[��H7�� AZ{ L#Bm��ʅ�3u��+2<�Dj��B%���ٛ���ƥi�g�5�,�m�CG�uT�B����C]���+k�z�l&.]ܕk�o���t'�\�}���Y�ҽkf#X��;:vӎ���=����t�]�.]�(Y��:��������{3�Z@��Bixen�לJ�tY�#��H��2Q���&��hTwg>[ɨ;���(����c��K㪲i�������5��ӓG�9��=���L&�:6��^�`���C��B+h�X��ө�A�x6��uBo����u��lM��rI�i��۲��o�+�0w���r+/}>��[WR��A��E�(���o,m�1Xn���r�x��\�.�T_�C����UUg�H�(���$������2���C}s�7��M��b�Вa� ���|>e,�d�$�jW��0�H�g�Rk܂ua"Xk�����Xo�N�m���	��'dqȅ�AY���8��e�ZkE?J:/]���6��v��X��O���òs��T�aD�P.\8��
^��Q5	�G!\]x���Rw���w\?���R� x!P;[��U!��x�w�F�;���
v42���/�X ���ߝ>�F4�����sp�����r�Q����2�F����������@ݜ}[��T��l�",��t�ۅ�����qbޚ�z��1�5H�I40���`�E���cg���9
r �\Y�ZT�;���sӝ-ݒ@�ӭ���s�]�ּ
�b�[�(����-o(��$t'�>�M��3#��tu�����q@:��@)B���Z����.U�(Sh��5����[�=�fO��ٗ��L�Kv#�`���B!����!����JQeTW3��*Z���?���P��D1n(���RHimZ�+3tD&���$��O�y^�X��2��OC��}�pdQ�9��s�E�N|����t�	��X�`�����v������rx�Ԣ�`���W�j��Dv�v���	�NA��/
�8�ør�
�ȝ{�����.�),��/�7P�:PW�	zp7�m>Ioh��k4l���"�Jޒ,�n>`�&d�L|�qʺ�2 �{��H.]����1��cp��d��)� |���d����!���D�̝{H���=�ۂt��x"�߹/Ý�,�[,�DY��M��������3K�:c���l�����X�� 5����6M3w��Y�4����W���Uʢ1��8)
;�u�x ��G�E�BL3d�(&��ѸD;Y�����єY���Ƨ�����[k	���g'��6.d�z�T�g�cƀj2D�/y^��Y@�M�ͫ��*E���CZsX�@H�l����ɱ����޸�jf���/Y�1"���r��b�������+^0k����c���.���Z0����XT�sM�9Y:�e]�U��}����*e�K����氳CbM�"��n��dr2}&?���:�s�xm������u
�ݗ�r4;щ���@YF&�?�Ĥ�
�W�	��A2CaW����O~z��i��̖�����;����dQf�qNٶ�əZ�ԁ@jP�Y�D��Od|E%G���n�;��r�����\͈>���O��K#�	��� b����3p ���7�!a�/��S���n����U8��{�ٜ�#�ӥ<x|,O��Rv�X�X6]��\$<����u(A���G.�ks����ߞ/�l�j�+��[�O�����t��3a�P�V���K�)��!� R��he� /̣�n(j�g��@9v|��t!^ԫs��6����?xR�\	���c��)��1bոѱ2"28S������u�2��'w�3�)L�
�/^dSr��ӓ)��R�}��b��apC��ƃѧa�bȰe�V�b�˕�@�
���\�4� X�z{��{9ܫV��O-@�2K�c{K�X�Ng�4�����.�pjo�j��G'��B�N�����.��^:).\�$�5�z�BZV�̅�e{ z�v���nb�r �^G7BX�B>%	�p^��g�D�=aL��>k�ݖ���LV��+uD�Bv����Z�F��	@ t�荟�� z�Ό�(8�Sf����Gk��X�51���ƙ�ꒈ5#�"�c���GG����ל�x�c������>��PN�kNZvqsȽ	Yc4�{��l�{��>^�*���|�֎/�y���J]dbJ�M	�Qٝ#�YYp���b�3��P�U�S��c691W�S� u㩑p�,�x��Đ��9"�4Mʱ�B�|#�y�4䆤H��%�V��ڀI}�ʉ{��/]�DT��ȍ9tlBq6�����d3��� �k����� ~���}S7�v\#����^a@��Wj����w��ͤCU�+�[Y���ˬ��rU�G��7�{O�RYC��fz��y����ɧ��������2�c"�-���������9qZ~���+��;���	���sy���t�z㡺ۺx{���c�l!�<k�Ak�����H�ͣ�����OeZ�r<Y�A9�T��yi��k�N�{�.�R�d�ᚗ�O�CXY��J�X�z��Xw�3�ﾧ��X�(�O1B�D��O��v��^@��(�j��fN��|V�ˌHڱ��H�3���	.$v����v��7�<dd-S(C#j��Ȏ�t
_d�!R+��hL#�>�ԒMF+J�Ton��߳W�G'�U�1�F[��,�L�;~N̤�6�o"ZBw��(�@)(�Ok��@�}�3;O�@֛A�6k���S��A֌�4;ۻ�ǲ����+"�dDѐ��-�7����3){Q�E/��jj.2/�����v8XP���?���{|CNPF��eb*W� �tQ�Yݖ���a1�j�0�:� O�9�S���y�FU1��'���~����?NNA^�1ҝ{����B~��O��gw��T����$M��f�rlp�@9ә�џ�'�y"K=��7��Q��l�莕�?=W�c&3�ƠKg6&��5(��\��|�l�^�=�u�.�X0a%/�����Ʃ3�b^	�V����lәx����·I���Y3����X��Vk��6�(n�����~)")�S����	u/�#A-5h�y�+c���!��M��D�|��}��'�.k�ҝ����ꏋ�����*-��J ��J����3ހ���F�<���C�����Ms������9c�^�*ҥ$߬>Uh.�w{�Ces�*��.<���qf(_�΄D�?�ëz�I��V,Ŭ�����8���{��@�jE�Ka������0b�J�Ogl �]��D�K,8q$�8�N@�.ZY��#��0h�w��l��4U�~UG�ߪ�	�<`�Ed5���h��{����zmO��d����TɊ�����'S�
���5�xF4tv�i~n夢��J��Z�µdIt械�EA��H=OEn3�E��������c��2Ck��B�>�,���yߡeC8��r9��DↃ	���Jhh��4%.)ԐP��uߚh�kğVk�³6�"�U�x��؏7o����@����ȩ��Q|�B%�ڮ�V���֑b#�py�u�㋸�$��� �֍�}z]�%�7��	qu���h[ɺ �Z�ɞE
��A�T�V���cFn>v�|�q4Q��wY��%_�j�C�Z�KQ��A�b󗐻���¢8jk�϶Gˊ� ��.�˔�%�*c� ��1�400�]���`���ϛ~KF�Pz+ 5#`ɹ���2P��a������9�4!�{W'F���ؐ.��R@�5Gx,�2ECH%�,P��s�,Q;��Ԯ���҈�D�4b�gei��"L�]�S�Z�������{�d^�-�Q�J����7�����Ջ����PJ.�B]�gF�@R���kn�|U�fUD-Y�Q�h�=�	�U��Imk�PgS�̬z]Y�H���2�1� ��̯豿�I����*������7��4"��I1�/nĉ�RY�0Vi�zd���MbҚ��g��"d��Lw2c����T�AJ�� :�����Ey4��O%�N�L�.ULw"5����״3�s�[V$�զ�w_����ԃ��yˊ�:���ر�b�*Z6@�u������'���"l=� u��DP����z�T5��?Ia֨�P>���q���NQ����e�nE�����\;#R�K�7��{
M��OV:q{t_��)�P�(��ذ��"4��ԯ�TQ|��H�þ�g.�C�gCi0|�+9�r�򵩔g^�Fq�h���b�Y:���A��N����M������v��}���s�_b��A�& � '���a��*�g�J�T��A���F,le-)G[¢I̅Ui�+|���@㈝`��u����9�������W�M5z��Օ�ϭ����ܩh�'�y-��\Ն��ѓ�/uV�X�eZ'LW�{�ژ��8M��,O=�{-X{�2ڻBڋ�̹k#���P�
��[��N���A�4h-]N?�^GC�J�PE�jl̨���?����͌DC�n�r8"eu&�|f���h`�̙���3�j	�9�)Pv��;Ϥ� �s����y���G�V'�$F)M*&VŘC?�.B&V7�Ѱ��Pj�PX^��5@ E|��Z��J��-/*t��
���y2��A')h�[;C��PH�Rx����t��wR��s�XJ��a��5
�IM���f*��lt�&1E��7ei�:�Wl�k�`U���Tk�vDqw����I�!���vl�U�2��&1A��t(�4ō9����(�cOdLj[t�����%�%26>�2T�#_Bv 
u�ө�*
��<����͢���֕�����C�ڼ+�"�[�v���G��H����b��^�t���O����躁W2=)�d��E�-��T�Jg�gnȩ�=ؾQJ��s7��rJa���f��٬�&C�+~we)ੂ%��0 Q(dP)c񐉶��3ʙy���\f .��9������O�0����Kp���s���R<�� ����n�.�Tv�2&׮uN��=�XVnŌ,��B*o&!7��>���F�gD^{�uȽ[�K'���U�Ҁ������<f����
��8hf�k��0�=�d��v}�+`i���8I���G�wy�$6�`{�u}�hH��(�Ӓ��qU�s��uJ���e����+��Enh{'P	�33�y
���A�Jv�3�%�$�ږ�vL�
��j����,�Y~nl]M�4�Tq�{n}��`7�1)ۗ�,�Qtq�^ �?tʺ�?���6�^�S�A:��+����N��D�c>����+�3I]�^B��k}5bHJ�w�7��p|�L�3`xW!�u �]�ɟX�:�|�(�<S�Y��LIh�[��t��]��-�����/ ��1��E]j�b�]�(ߠ��������=fhY %7�Whns��S�e���^>����\qmo���3^k+��^�ϾL/�Q�����B�z2oJC���mK6�H����sfF���fQ��,j+�u�\J���9����_�rC*m�!�7���ɐ$T��gM`ȍ|&��ϙJy�O�h�N��
u��
A+�Ԝ�|�҈ m	y���~k���X�}S���B���x�t-u5qk��S�!w
$#����~���3&/��1!�,c�jd;GTuJ[�#���A$ԕ`}04���L?�P�sY�	"tCa$��HLH'���W���m��F{�+<^�����8&��V�;k��5&A��ׂ��F�u<���ZG��yY���'Z���j3Ʀ��؟��;���Z���.[x��עl`l׊
��!��x����x?s�?����iK$�X�v����1i.U�6�ҳ��ׁ���[(��@��Z��^�o�Ӗ8y������ UQjN�yU�XJ���Ox��ě�P���+��\�Y�{�o02R�hT����J�����妥X�	ŵ*��CL��,��i�O�nBe����d�]�tB�ڏ�ln�ƠWW �rA Ϛ���뎉LR}��h�ŲwJa��E� ��{n0������4��O����˶��0W��<�&��G�S��E�&�6o� ,�1��&��p������`�����;�-Y��Wy��\JF$�-%2$��P�4A<��Яg�$�ЌKlj���&M�4�(*�
S��W����Ǉ2��,�]Y���U��"ш�ĥO��W��W��[�Nc�TK�1�Te�ĥE����B���0��^x>1��m� PL��oi��!bt�\�>#Y�s��3�Am��� v\X��2As��D�u9�1����G.����G�ueK�;20���`S���B
^kq��}����DZ���o�݌�K���?��?j�Η}0���R�?��p���:\��N�I$M�(/���(�X�
������&��/$���K�C�@�����^�'�T�z=�r]��6Q2����IQ�q�*�O�e�;C��ɰ���Fĺ�����#����V�˾�ƭ�j�d����L�-T�V�J��\�IĨ���!@\�����/��i7����2�L�6u��g��L�����XY�+���+��E��"�8��p~d�����<EiE_�������n�`\`|�4H-I(�Q�13c�&ž��~���|���&{َ�2�8������k�C݌`��w�iͭ!�ŋ�uQm��6�J�PT
 �V�Ő�u��Kj�󳬎f	�����Fh�o�Y����{��k�^$Hf�$����t��#u�D�3���4�Mأ�#*_%K�7]wе߳�ZI ��O����ۤReIr��UR���TܕY��%��Z��P�^� ��B�]jB�W�]�v�5JfuC"��מR�S�,Ye+��/���<&��`#�f����u; ���O+�~d�li`��1%W:�P�� �Q��4a�?�eZ����B-+��0݋��O��/��2�Z0�� ������ h�xz$�Ӊ���.���&��g=VТSp����$�Fvь�G��E�ҿ����=?��O���r�mH�5��Xnl��,�+}�A	��
�&��
Ж!C*6)�Πo�gd�Pd��t�C��-:�XZ�t+C��k�$Ru{���d�65h�Y���@����ӆ�b5��$��-�$P50���\��b&HM���r��R�(�eU0�@f�l������XW.�3`���VBe-��g�)�FJ���z�T
�6�Z2���?}a��ema[����_r���R�1�]p�A\�!Ԫ󶳺�M��= Q�Һ���b|�˥�I0��Z}�X�POpTA�g�i���I���j-IS�f��'1��$1���K9�+��X�I Ʊ�
�Je�����'��걦h�ཀ��o˥+`��\!��EO�y��Hr��,��_�e<�v�48*Lm*R�ҿ{�BB�SG��$�(!��h�(��T���5\�'z��&��5Ȧ��S��gC�(��,e}��K����Y���s��y�t����T.E���Q6k��F�<�G�ra�ռ�e_^��ô�h+��,�}�W�5|v� N�ϞY0���1��CZ�uL!�ę�M�w��x-��} jry��%H�L�K��w]q�ģ�C���`ǚ��k��hvT��Cl��R�{H_-8�Tn�2a����Z�v�E�dC�S��O@U.i��������p��m�e�g�#�4Q�Ə�:��H�_�0�D<�μ;�x4������nb$��O%��>~���A#i�0���4'a�S�1k2kd�zyj�J�'���+�Ir��.u^�R8��}9{���Iu�r&��QmT�z�Ϻw"�ސ���lTY�����n��*^J$��nx>�ƀ�hk �=�ui>>��u
R��ac<^����5b���դ���?7�)�C>�ٲ�&CQ��N�m[ؐ�ΒҪ��E�%�y�b/3䑹�J*��!����F4�Rt�ύ�&\�v����0��F��Z�V�ՙ\���Ku���S�=0s��/
��Zzɭ j��g8<��2KP4�byxŀ.ݙ�lZYr͞]�g�l�OA�x�c��Llb%)���Wt[�}�5ȧ�_�}��'�\�C������7���N�/c�kN�����,Sb!}�R����8&ه�QK�y|&��l�Y�g����Z2��Z×6�3����[ߨ�IS����b1@[��8����,���������+� V�z��~^}-	Y�:-�|��5���*I�(�	�v�R�$�&a��$������������p�]�:��V��q�4�������%�M��g~���3�)��)\���*��x~�J� �2��5k�}6�v�ǅ*)�\�ƪ\��j��ER4��UI��A�������-��;�t�M���9�±����f���C�Z���{�4'cCpk�e����}}������R����w��ݙ�?cEg�{*�3d3��59I�c�qv�F+i���U4��Jd��MJ��6R6���EiCnPtB}#�Ķ��z�����]��Pr������c,&��V��!�@
v�#Ȳvp<�]���Ϡ��f���ko[�����{/��4���o�C_r�d��4� \����H�a���vXd]�э���S6a��Iٷ���A%��u5$�� �cl/�ٸ�@Aw�*SCj��T� PC�u\���-�!LD#S>�����>#����a0X�z/�@�p���̘�e� ���62���sTVЇ:R�\P�g�����<���&�h��ޭ�΄�q��b��9H�7�p����/�&Z�m�w{����&�k���hR?��Y��:C�\b���bJ�� 3!&t�����O|R���=�[A�)�OH&GT�[��)�ⶡv�DR�7��8��2���^�̊�*O�>��k) J�EY5���q!�F �	��w���}򗽢�OP�-m�H|5����xM��s�f��]P���pA/����~�ݼ��3�VU.Ē����*������o���sf;�qj��x�+2Q9(�B�҂�c��2�fæAC0X]'�����HivK��+k�'NR'�E�1+���Tȅ,v��kB���ŇA\���������ژSh	�(���B��5n觍�hl��-	5Js�@L��n���	��Ƨ���+#2��tN��qj�7PӔ�/���-mFQ� /��sJG*�B)F���s-;�FȂ�oP5Ǣ7���!��r�ئ�آ�] �·lG=������j��ژT�68�PՇ8���_4�����2���/2"6,kQ9ܣ����5�P��1�i��w]��n"٨�IA��7�	�i #�'�����d�iM��tS����.i�Z�D
yp�GOyR~����l��j#��B{d' �3=��d*�%�N�R��U'��˗d~�6i�;��LRK����Wh���@�p�B��ͻz/�\]h6����Hkk*��]������?�8��>;F�Y�j�y�e�q�Ya��YymO�>��G ��.R��SY�C��$��tiH'�����&�@�'Kt��V��vw$�vd��D�*���:���*(���D�偘�,��ײ�n]��ґ���o��_�:�N���`qLce2]�L���N\��HA"�Y�.ǡ���h$������p"r����M�V����.�z����S��n���R�*f+�be��-(ޝ��Hsc�l�eYQfw�J]�AdA�FC�4b.�`���T���oED�]t',�K�,\����}���f��Ȭ�p�L�U�;[�Y�\X���Kk��
������%�bsEZ�������I�7���h�D����+�����;GH�B���μ�ϡV��5!�o\yj5�cvÑ����t�6D��7iG�7FETĴ�I;�X�z!��#Y�>��ڬ,�߽~��%d�m�	���I3�҅uUo��:��G�X�hT���P�3���Ieh�0:=�3��r���h`��ذKت9{�
zX�t;:� m�3;����T0�g;�f��8�uFC=a
j���U����b��}��N:*�pg][�zf<
�X�,v���o6[R�u�5���@�����B�]�:���t��R�n��;:��U��vn��!�9���/��>/t���)�P�d�I}�]u�����v^��Ρ錨�R#�__�o��8��3a�Hin���k����7V��9�>�%����رY;��n=#C8�6b�X�q�����O��X�5��`U����xPn����Z���,=��.cQ��|��x�J]���6Q�~��M�6d�tá�jb~�eclH��-7j���&�J�PbG��Ȁf��p��	�u�n 	@��0�Yll�St�L-|��h�v��|VO����q�Y��D�۸�q�m��&��Y�^���"@��uE�l�}@�~J��eSg�츥7�fz���{�+�=��|������PվY�lW�]�p$/����Q�Lb�ZD>g���\kJGR>�� 6z�B��}w��:��֖�{����+�rN�]YN��xeͧтdop �B�XD7��A6}�:]�Èb���D%>_��/0R��ֆ��\���-�XF�OԆ��H#��#f�˰WXLL?�5P�C's���ڞD���j��WQ�dA0u@N54#���>ǲ�s��{
��G���yl�k|B�r�i�>fɅ�jg
݁r��ƿ�:�$Ϻ1��JS�ԭJ}��s/��Ŧ ����C�犬�:q�,!��M~���q�l*�꘷{�"��#
N�<�{Ƅ)�A�P���)oW�k��aL�Dw%,�l�H�OQ�����2�� ot���N>R7a1c�B�Z��@�%��b�@�n�*d��Ɔ�뎜\쌊tV�� �"C4(�N�7]դ��}�ٜ`uT�H�X�y�� ��.(����, �jҟ��.��:C�#�	�u��sB��x*��}��{TU����J�$<��={Ν<et^��|�Y�����jt,~#~1,f�0�z�nFݑ�z�
�O
��ߺ�]��qJZv�����U�.#���n�����:��
�xj��X[S�����b��ӗ�Ih��EB�Q���ZO$��=~|"��ǵ�M���֧���b���El��{$�K҅���ԑ���C��ni���Ep�]�ME���]�x���:��d����껮Lk>x\G� ��ա4NL2 �H�kp0@kG�����T.NNt!U��R%�=�f�u��"���
��F��ס�n ��W�!q���؄9K�`�w��z�j!���-b���3��f2�5�fX�oCdU���,w���h]���� q�o�=� �9��	T�z��9��Ǟ��2���૧�hD�<cE����R�}-}�p��T�P�(Y�^�3�Z>�
�KI;����]��T���:�<����*_L�A�h�kf(�Z3n�8�8�@ǅ�U��+�r�`(�H$��M�Ag .)�m �V/+�9$"� �Ycj�|N<�g|%O��3n���J#�C��b#�?7U��OQ4�n�f���N�c	m��yM��-H�����/����d�p�ETS.l��D���R�L��l��&�h��ů����l��D�bjUt�t����ef��R���C�T@�⇾��pC�	��XI�v��~G:;�h�\�����q�P9Bq�a��W���XA�K<H�2ydz��F�]sL���9�7u ��O���"ܮ�?�C�}[��8��ў�SyO�ܩ�%?nf2PWr4��=���R��`nmSm��hg�{@;|�y�`p�;�aI��|%�Z�zN��v�u�z3�Ɔ��cP��\*V(f�0)�a,�;%n6�[*(�@2��H���B�u�E���Ɂ�n�k�2
8��x�=�I��S�1=�WfJ_9N�Ϛ�x��4"dY"CSSr=�P��jNPw�kPȹ/�wLH�y_��YCB}��`�&�$Uٳ_([C�4(k5ʹu�]�W�t�{:Y��E�R'G�g{����R�{�{��e�l$��+L�_y�EĈ�j`��du��i�l���'�!ޱ�֡l,�����e��Z��,X�/�C���lR�j�e�G� 0�E=�y�������3]s6��1-�M�Yk-�(��݋��}u�^d��,��"���ƥ,7s���P�C�^�HO�8j��l�3&�v�)`2�AZZOo����Sx���*so�ܫ�lg��M�g@V�d{� �V��wu��T7f�����`腩��+Y1��u���Z1�JI΍�i5�&�@��M�,���*+�t,y�ZJ?<���GE�8/X�韵�\R��e�	�ɏ?��шM�H:���5�\�z�pk�v���������R1\M4�M�"�)a�QuYQ�r�gf�� `�l��ߗ��D����#�pJ��vF�L\�t�6�Q���@��ua�.;���Th[Z}M��C�UD����� `��.H�+7f\�D�s�d��h�ׁ���e>P�eT\p�=P?�ߓ���#l���!���Ib�gG�� ��X���m;�]8HB�:�A�r:/�
#���@���߀��{<9��.��<�-W���p���ի�9�<��#��sUy,��^!�mj�xns�:�i8�zlt���Ϩ�n''�<��A�E�@���n�2�WA��cf\��\�,	N6���F[rrt���'��=��a��i��%�r��2�62�ų�����1TD�M���{oC���N't#��(�Z� �x5����;d
NwP�o�o1\FfjvLa�sB8	tH6$%x�e���vNB�B�;zl����th�bN�d=Roar�b����=:z_�	����ig� �tb��dB%(��z�֝��D�&4n��L�8m�.iwo\���Bh\�р���LV3���X��z��"������UaB4k�֬,t"L`�=��C�1S#�B�q#C4vFX����<��
םΆ�4R�{d�FtU6$�&e�r����bT�_��k]wk�7[L9i�u�s�Θ�����(�@ չ5���Z.-�&�l�`�2�������R�Y�'1�h���N��&0���R��'�2c��q�Z��6�Q�|5���UD�u~Mu�.�/�6W��Wtg��*Bn`�P���͊n	��@\��fLE~0j�(:��qq��V�XN������S��a����z���
6?�r�T����#��������П�rr���(ڳ��m
�bnq
������	E����DQ�&5fjD*��w����*�`�����e9�m���HQ�70sXS�&�� �vZ�P�qiR-R�O��-�~�_��QG�x)��z��(	/���c�FP��n�k�q>;��z���`�9͊� G�_��kg/���+H�����tw�̧l���(�+� �M��j��܈�PlV2k�����Dm��!]@�M�a*=k��%R��EȆz=�I��w���h�Dz0�J@���<���.M@�}?F=��1zX�������x���Tp�0s]�e'��@a4��V��I�"�� @��q��<�je�޶^sGwbд��3#�����{}<_S�7��Pt`���;��A��?�2ޝ���� �Rd3[�pԁ҅���1�C���V��%mtg�>��8`�H�[��p<P�:t5vhut����z���5"c��m�"�%��x[��E/<&�2�Xr�����L�r�|����θ/;��|3R��	nW�6�=���s��/�J.^8�X�!A��B���	�@���s����?��Z7�������sDh���q����Gڌ��9>����U|Y�&���8]N�Z�B"��5"�����ߗkW�k�����<�:�oD.�$Rgk졇�������`j����nzz�.WO:ܬ�r�:������@F�X��V�k�kL��Joi�YɢZ��:ؕ+��<ZҤ�� m�*2S��ɴ*Q�
�=$�H.[[�/�w��_ZSq�����H6+5b��w��&]L���\�rY�]��"��K4�Bv1���}���8@Cj���b��L�
&9X�b�)���&�i��,x|�;`�7�)��+5|�T�N�f^tMu��@�����yTC6W7 ʥ���^�ݭ-�+�.^���Hn߻#�oߖ��X�a[��]r���P]���\���}��)�:��۲5ئ�t颞f!O�=��>�>�X~��'�h:��[�,����O�k�����Ywc*�o~K���[���+z?]�6Ē�:ߎNNXyЖ4��7�v��1��jdi���q�~�X�+��њD�������������.�g���Qt�����Ʌ4J�H�" ����Y��b$���5"��Є	R5s;�ZF�
���W��>vU�����X3	��]BS�>�C�ڠ�<��ߕAj�(�tl�
��_���kW��!gV���Ԯ�*W.�X����Syz|_:Cp1r��V$ב��C��뷮�b��n�W�.uҪߩ��Tw����������>+(��94ܖ:8�.�ی�1a,�}o��s�n����M��oC.]��`%Џ���Q�QE���5==���=������{��t��Hw�9�轃,bT@Oy�1�W�2��?�@�����*��'N������!�[)��t�d4�@ll/��`s��颾uyO~�7ޕ_���v��o��z� zx����V)�2��dF���]��Sui�v��03�	wn�4����u�PC|]��P����_��ߕ��_���Nݜ���L��Y������>���7�����|��7d~�L�t��~>`|
�9ۖ��D�>̠���K'��� i<�r�(���#}é���M����?Vw��?�����{��Jm���de/�P�ܞ1(^�<��
/�)1-�3߿�+����M��@�їi�~x������P���-/�RK:�9���Dmҍ���Q!p�.a���|���W�%�]����ϟ��S�$�v/�H�œǇ2߼�^F�0�S���
M�uG�R�=���#}�FT���4H�/t����#��?��iȭCZ]��rژ1���� n!��D��H?_����M����ȷ��ק�lw�K���gW�X��|&��C�����}b]"��rCw��-��W`Pr��ϯ�j����O~"�>��~�Z�VwP�|�X��X�U��&jH@�[���ڨQ}��e�G���w�r���g6��FOc���L.t��.�8���~����)ٺڱxN�e� ��L\2Y�� e��Ż�g���_�����_�����c�X�/��y^+�zR�A��A)��C���ߔ��I��y�s,��|Q(��d��t��ŋ��o@8�L]8�G��!�e�cMp7n^ڑ�F��}�;�(���o����I�Uϵ�m���ڡ��6oR��r��\V4���J�U��2��=���s)^��̼��'�����7nȵ�2� ����l~v���f��H����4�N^]p'v���#y�k��έ����E�W�&�cF��𭁺����{�>�L�=�]Y��P�P�8��A�F��몿|邼v��� u;�����M��2�軼)�NY:��X�n�����m��Eݤ��'�P�|�b�q��e�}bGr�Tц̘��R� ��т�mh*�D�Ȩƥ����
�jЯ���{I]�~``:����v�0jWz����w�B2�
C��{��
�$���o��/�ޖ.��3�,a4�2m�������G�@�#��VRO�ص"$���[ç��,ut��9"�"��tt �@V�-5:���:'�YJߞ�9�7Mc�b�ݺuK�P�q��H�����|��#���#9<�ʍ���>:|J��L��d�Hr8b����{jx����}��!ҿϞ>����}�M����-���v\D����XQ�@砹�+�	2aZ�%I�c=��]�9�ъϭ��"{��r>�F(���F�>�d��t��q]`�;��r]��x ��Ӫ>=F�Z!O�i�A����������	Uf���)�h�+�4� �����>b��[Y�Z�1ĘnP���'�>���P�>=�m���X<W1a�d0� Ȣb�GϞɠcy����k�ur�O�PDy��5���o�.�!=~���8��Kz�
W+k�=t�V�^G/rc;Ka�&�hT����[=��2;��b� �}��Ňȃ������>�I�mX8���	+���(��sM@h�����8A2B:����|�k��/�-�A�M�h_��12	m��������NYHz�t�FE_��@�͍7���Ş�N轨{������u����e=�P颻��>�+ҽ$��K�=bDcE��;|�H�?;6�&��j��_����ߑ��}C�	�^+���Fb.w�y �름BlAB�t)I��K��A�ɱl��t�?||,��������x�mJ��A����7B_����u�uz���La���opG&:����>�g�?���Hv���C�h��_D�ʰﳻYV虑)�C$�4�{���
�L/�7�E��&:%#3�r*�e��`k/+���,��lP���%L�gGO���ɒq�$ҶI�.N���(Z� 
o�6j7T�;]��/����&�Q�	,���-(h�%���O�뒏3_�f���W�q�h�<���|������C��_~,�<|&�р��x+�=1
A��#N�n����O��G����Ç,�/e����n������g��F#�êV+N���$�?�0J��,+�F��d�D�����Eu�~�@�տ��rgcɽM���*rt@ƲN�s���:�����d��(X6N��������x2��n^�k�^��X�ѩ�U�>"Y���i�� �p<��z�|���~�'�"��}E��������{��=]�c9Q� ȿf�ɆnQ_��޾.Xuúk]|y��X݀J3�Yv�u����/r�ꮼu��p���X�I�~16��:�yi�i��-�?���m�u��r���~����W��|v8�����Wu�)����18��`4�aƾ���)$\�S�M�"8�
k�����o?��I!�v:�����-9E��hLd�c�*�.f#5G])vj���~r�c"�1��4�V����[����ޔ��hDR�2g(d��XZ��j�3����Y`�T&��]2�zI+���j���$�s�.t��x$o&�;{��$���I�kF��%�K�s�s��O�+1%/,�ao ��X��؛ʸ#Ȳ���$Ef�љ"���C9=:�A��϶Z���S��T������?YB+ē�)P\�f�<�"-<V+�)iF����so�l��y)�QO�zꪝ���]�D00Xt�]:����2��X`5�dP5�=HXAw�~_}���Ǜ �������Y%r΢����ג���8��r�����d;ߑI6�b�Up�ϦCm� ��^�v��W0nGęДY*�OH��(.��H5A�D�c��6��tܖ�
&_E38��l#)Ζ�Z���8��BO��`�i�78�>�a��ZP�ډVܘ�`*����xGv�7��>���o�
0/��e",B�E��~�ZJ���C��a^ur#�6�ʤSQ/ĲjD��&��3������Nh^��x`�DAp�K�� Q;'��4�5���5�����ԑZ+'7���	Kt�0���>�%Ӑ@"�$��k�45z�LD�{����g���t��s�3�AG����;����k��G���5ʊ�y
M������r�J-��r��������iǭLn\?P���ә��ݑ���BJ�Z2�X��k���c.�s�4]G�_�F���U���d1=���lײ�mV���ka�?)xg-+�+~U�f!غ:=����o1�����؀��a���.wǙ�w�Ŕ�n�{K��R�$6�kz,9��r�߉.�<�>�����z5��r�
a����Ʉp�@�<U��X,e����Ξ��v�P7V��:�[����O ��b^nm��+O�Z�|;%���C+���E��S4b��mE@��Ȅ�2k2�^�!�+/{5򐍻����u|�xh\������_mD�[!^��L?�J�ė�ry����m����8? k`�&�hB �@�[�/�3�vE�t�E��.�!`p !˲��u3c��N�
�L����4_��F�����\��AcC"�͂59F��4�J]�%��7�P�8�<��],��KXT$t��N�F�ky��"��Q���DI@n:��-"PN��� t�`=��>�B�.�+'gYi�)cY�+U��C��Z������-@$��F{��'a.K� �eIM�H��@(��{�}��w������=�+Y���/�O0�.υ�)�	k՗�=���*h�FM� -grz�L]<uQ�[���]��_�5dKyvr_���sq�.�@�1����}Y�LY
0Tw.����yKpGy%�I&r���;j��CZ&gY��:[S�Z5lH��P>H��"Z\���?��/��ۗ�&#"�NI~��J�@�J��SB&��.I#A�xI����t� w՟EK��9�3�+��,X��[j_�2��b����?����\�:&ө��;�@t�C50���1��x ҴJ�
�����h��om"+D=t�c����T�.\j��|�P]��\�F*t��p���ymW��>{P���z�����˿�ţϸ�2��zlt
9�����3��@�'��I�:ژ��f[�?F6*x]�H'Og2_��?�d��A�w�z]vw{�T����@�}kg�,a]�\<� =5�W�_��)Қ��?����zO�=��C�����t��V�A���r��C�Nc���3B+�F�/�6�$B��/}��[�7���rt|������\�r��X�>�z������l ������=��쩶�s���5�}a�$�	����YΉB
ts)�����o������;��F:0�y��Z��R����J�9�]�Փ���J������_d�:�� $�W}n�^��_��*=#�ݨd,���U��(���������ԏ��~��X������c�Sd�T�����Ǯ�l
�bƪ����9^���#C�wI�^0"HK�Ҹ����w����-Y��::�ɥ��k�䭷���ܹ�;�3���#����M�{��ʃ�6rЃT���hJ�ծ%\�>ɒH�&.� �˨�
�Sy|��2s�VD]5^@��+"�����v
�UzNEs��~I~������}���]���U�.��p�h��uy�w䙎��GGr�����-y�Ҏ<��r��Lu�-ԎM�>���]������3��e�bFu]����X�F��!
Z?��NrC���w��\��-'�����ܒK��Q�}z�����>9|"�*{�L�|�:}���{r|�@d�ʀu?�(�2TWvoo��h1�ӝ	u|��\�=�$Vݜ06����.bE��1�����W������\Ip��PX�4��M&qy��9-&u�ft���Yyu�K��Z*Q���8A�`7� 2���d�8� ,�cDdq";[}y��u���?�/�x�^㕃��7ޑ��H����G?�X���|�ޑ˗oȃ�s��O��9I���r���L��!�n����/X�F���N���74S�,��V�P��=��O#�@5�'�����~�����{2?}*�}����{�y�s����*(b�����s�ۿ�K��ٜu&}�����'���V�PMC�ke�e��)���?�Y�wҳ6��V Ja%���j��XM<�/X!����A��l%o�ؓ�{{�ke����c������t,Nt|/˶�;����c����}y��w�׿�+���fS�����?��ߗO��uF$xa�=R�"Xc��^u����o�er����h@�=cY����9u^��U:n��(4��?�?��+���3�|���2ݭ��z/WnHkG���ٿ�F��o��������2P�Qy ��D�K#P�漕z��P.B�F�;&"��9���y�,`B�[����3kNB=�����^�ϳfh�2";?$#Ӕ�҈PKoP���UAPs�n�30O�\�E��l!��|9�� 5��+<���i񬫃A-�[�T�M�M��2���t�����?��������|��{z�s��������_�}�P�.�J�����D��W�z]~��ߐ�>��;��*:����(�|(�Vh���}�j~&�C�!ذ��(����+�6C�ڪd��c,Ԉ`���/��٫׮����} 35��������d<��s����+�u\�t�c9��W�u������� '��J�a0�Nۇ3.+���L�=����d���&�l������������ޫɒ4��Z�%��ZM�LOϴؑ���� �x `�4�G�Ƈ��F��H��$ �5r��;�#Zk�ե�2+���ވ���_ĽY���m�Y��yoD|��~���qU�Rȗ���ɍ����<.�RQv.\������o��{=\k��g��n�#��o���T��ݡ��W�a3oJ5��Wޒ�MD�L_t*�6������d���j_�ANrAH������[rxr"��k䪜�c�z�̥;���o�&w?�T~�ۗe[ﭱu��a�� ���ΚGj$����晢��&��L�#̐	K�s�ߣ1�,�����Ҟ������I��ߡv�s�3���܇�IB+s�D/)X���������6>-������G�A�c�d�b-�I>y��M?�9D�Y���j�,VQ-�fNy����+�G?���W/x��=9<=��������/�+�����$���?�S�/��%�}�'��Ι�E�\I��������z��Ha����K��=���@"@F8<HJBd(&�*�sVQP�e�S7�2���3���wE�l�nK�qC��=ill�K?�������t�9��j}�iE1c��:rxt_��@�7�YQ�����B�e���̉Lh<`<����&��v�q
����;w���{��sߑF)/��~�@N�}����t�}�rQZz(�������˻�ܹy[.*J|��jL��W�_d��g���^�g��`fT�<�=C(�i��È2�R�~�x�
y�;J7!��S�3����OԐܐ�<��n�ID������z��-�uѲ_�ߨC�Rý�� ��ۛ��V���#Mը���?�p���8��'��W���B�|�^"g�6R���92��;;鿻3��%u�s��X�,]֦=G����8!"qq3����7�D�JP��?#v���¯��?�#�\l�TM��y��7�"È��T9k�m5y �ф��H�7ߐ]`�l��E><k���-iu�r�����ɩ9>=��?�T.=�ܽ{"c�Ցz�)���7�6&��D�Z���-tKx0�a��Bt�p 
A�F�w3Db�)i?���z�VO�x�Iy�[ߖ�o���?%a��&�)����[����;�n_���m5�9=;������EhIo����e� ��Gdm)�1�𵖘L�sɪ|!�c���0��W@c�n����y��OdU����
5H�[gy��{o�i����R�����k�ʛo���כ��GI��+C���Ӗ$,���z��ÀL�zcRj@��|�Bpn_�ϛy�pJ�!]؏xV8�Pr/�!F�O�٢t㕫��Rk�5t��Ƞ�ˠy_V�U*b��æ��S�Gs5���-G'=i��)RO1�8X���~���D��K�����g�@���p���$NYU����G���%C���+"c���Lr��1��dc[~�+x^b!�ra	����??L)��b���8�P
kȑ˳	�Mx���"��Z��z��>x���ΧGG�{�<���wޕ�G��n��,CJ9�}=���8���}��,h;��V�ga�� �!�� � ��$�@G%�_T=��>�����hپxYv.^���C�?��'�2dyR��KWc��
\������-�|,뛛r6�����S
X=a���]<�t6_�I��ɍ��7��-B�/�z�	�EQT�Tn��]�v"O<q�r����?깜�����5l��s�]��rN��ēz({��ǟ������Äޚ�B�ӡ>�HrlFX�(RAN��;4��8D��F����PI�xy�����l鳂tc�~��z�����}�?riM��[wE)���CTi�Z���E}F%�<V\V*5������2�TI��(��r8�p��\y$�T|x0?d�L�&��.��JKcW���r����
}����d�N�G�f����c=T�L��wɀ��DinuV��S�-�U��TP�6��e��C�u��s��հ�o� �#�󤔍��u��}9:�îׂ��W._�v�Tڝ���9k�АFC_76.���9O>������akx.�c<KNMt��0�띳�^����Ϲ|�0��{z���qs�֏�����z�j_<�^pE�	��p@�7��9���Bxwrv��{�_��0�Jw�T��!����q�rI�����s���8�P�phČgD(�A�����dk%�sK���Idy�7_C�/7o|,�bF����<��s��������/��lsuM.n�H�K1�Y25"j�b5�=JdQ�sR+U�����-�Ʊ%��WM��K(7�����.q���{+�����|g�nh<"5����F*�����l�D�:�F���I��vw����:�,N�C���+�vs��	��|!k󘁪+4=��,x"4��2�IϚ��Ck��X�8J���-��<7��]�!6�aK������!Ùd��U�.
���q����Շȉ8D���Pa88~�"�=8H��WF��P.z�6�I�Ts�Y/ȳO^�o�'�N'3�gS5�r��U���t�&a�J�:#�h�X���'�CE#6���]E�5���f�	�>J��[�L.WU$Y0�;$gHP���l���Ǥ�7OO�ݷ�$��zs�����Y���1:'���� K_C���9�ҹ?a8��ȋ�YA��0�7H��!"14 _
��L~�-����@��;���� l:�S�����#�Z^6V���&��}meM
Q�JME�Վ�8��P�=$GҨ6�[Kg�!I@�u>��q�H�qIr"ҟ,}�\b�h`nz�0�z����T��]ݐ�"���+X�!�ύ|�� ܄-PV���-��A����C�Иy�ae�H�Xg�*"00@A�+抬lR�?^������$u�KNy)�8w���gȜ6�f����s����� ^�Bu�_�'p]��!��K�PhHR9ɍ�@|�/Gx�E\\��\��dȑM����9Vr��닓y�SB��ޟ#Փ�PN�[k=�i�X!藍1DG�҉��ƅZ��ɩ��֤^��%���{�	�V����UC2-��RN�z�[j|VVw%�R���:S����������� ����7Ɲ��4#W�d�'�'@�.�9�Xx�P�M=�����^Iz�#=�]��st�$��@����,QY���T�D6�E����B=T��Q6��k�V�R*d��q3c�}�6��
���_�i�h�`ݤ9���_h	���0��il#%����D1�x�'W'�2olЉ��=e�H�V�jc���r�!�('1�E�Ԩ��ᘌ��(R,���[��l��Ӄ7�Aؖq�s97*�=J�����n�4=���?D����}e�}JS��M��FCo�5��7{��� w�\B��>ʲ�h�S����'�g99�(2��F;B_�dQÚ����"����5�
d��5ĉ	m�]g2c�Ȧz���o�em,OlڻiXg"G8Ж{�ZC��ca�I�1��`w�dÉ'��K)���!H��_�DҊ�jƦ���2��H�ڿ�w拚�K	��;����PF��d¯���K8X�(J�ђ���CRj,�5�Tr��C��������+ץZi0���#{|r��-'͖z�6Y���+����J�^&���XJ�QH#&�9;�!��<���!EbןѠp�v�jp \a�8{h�W�y�̰�~i������R��W�UI�O�Y��53�t8�Lr�6�*h}���1��`�Q���P�l�"/ 6�ȣ���B�$S�Pd�.�4��~����*✤��nHq�C�=5p.*@o3$q[|�|iMç��gH����&���"�����a����m�:�C`�!u�2�r��t0��^�1�Ƈ��S�dD������!sb�!a�8W,���`l}��@�35T\wE�Q�ˉ�!����R;$�jq��lU+j佩�>�ҩ>{��b>�T�%L(���zU���i(������qP��k�`�`�Z�n��g�,s�P"�\#�U������֘�<��[�b�Z�ȞO(څ�4�j|��U͂�I�F6�s":�D�E[�Yy�L<�������.�RT��pa���'��س1��	��c��;�H�s����P@�FW������g����"}�G{�r|�Hz���N�2<�)ʙK0����}.��_�l}E7����4�0@�T���6N�`K2)MΡ1��K8��i�2+s�iY_��j����!0)�0n�]�kԫ��+z��&N��'���C�����
ɛj0Τ�jIg�!A��J��~���?�[y��0��wd��p&M\���y���ĩ ��3���>���2-YiT٨7V�Ű�^GJ��䢑�Ի߽ѧ7o�Ak(�Y)2�����Mi �� D���D*�C�c�S�)���eV��s"X��4��C�SC[�C"-5c(�k8�D7d/�՚�l�ȥ]��f��?�!x�s�Q��Ѱ��?���N�_�����Jj4�2����t!]���5��4AR����T]��p���C1�1������{n���M�H#���c��'���Fg~��ǲu��� t�N9-^8�����2x����l"�A$Lf��!��>��P��]
�l��������u��Ey��k�N g�Wo���D�AN�Ū��Eh�s�c��͜�GCWse�����؆���K]r��2!�[�NW�����o<?Ӑ^q�?`_Ϙ��V��Z��ǣ'����H��AGeTv�s>#h���}9=:T#�)�JQl6N����fKQ��Y���H���\h�P��	 ����S��BAj	ȇ�*b{������N� �]-Q���%U��#5�G~�<����}���@j���EEd�|V�
E����˧	�!s�:]7�5U��¬0���� oxQ��W/˥KWdcuS��F�t�}���aM"��V�rQ6_����@�hh9
��ys�l�H��jU��$˙8���%K��XX����3��� b�������I��FRK��GA��yC��������5"���]`<�&�9	2����x�E��w�t���gycj[�n� ��b�͆cYpE��g�}F�z�q�����mv����!9`y�]����˜����p�)��k���Yxx���D
v����E�,R�/�&i��������ʢ�2�7!�����^�X`Lb�p�y��������z�>+"TG��z:��΍��z��!O�3���M�uw_�����-}����6n9�1R�˥e���&%>�3��n���g�b��'!�
�����'?�)�/h�F$�����Z�2��1!s%S���5=��Z�˧7�2g��R�b�9�H�fU�XI��9�����M9#9�$����T<5V��n4��Xֈ$��R.�$S@�1K2&%�w:gl8/��a�^��fkҟx2:<c�
V0~A�3�S=E�!�]��~{��/�K�v��ԲaY�cJ�p�E$⒵���E�I<p��7S�-���!�xus����(�R�	h�ǂx����;Q���E�Gn|���C�J�	�61��ި�:��c�ޫG�X(�4��Q�K�40�QQ(�gˠ|X�Rp���-Ҡ�p-V����?����
��}�>��1�s���Z}K�F֡.ŖL�o�L��ə��V�Lt�M��G{��oQ"%D���*�������5ʱ���jՆ466��k"�r	j��~�����kd�Z�ܳ<B�H���6`z���ă�Oe�탙O��6-����A�0�-���:�M�c3c8�J�����D=��u8���Q�*��u�=9��e0����Xh�:��dc��øO�3�����:E�p]z�\�&�y���b�*;�r1�8ǜׄܤ8�ƴ��o0]���^�i��,�5q���x����(��9+Ҩ�S��i,;��{��Ӄ��2!-A��"���&I4G$➙�}DD�ah��  ����p��Ym4VfoĄ��eo���zCB�� @�-��a嫈/v�GN÷��w�TS��f?�6��(��qM���� oQ)W9m�5���������8e��� 4�_�
ٸku�c�SO7����X����*WozC��I���y�ːz?��)�(�AM�1q��F�L�VOêj�ArHc1��ȟd��qŬ�YY��ǔ�óm}8����ID��ýXZ��i[�Ȍ��3�O1bX�d���Z܏�Õ��ƶ�L${�E �^�I��Y�-g힔*uE
5�]�̑�9I�8��r~���z����@�?���	ƹ���0�$_]�['��;���ƪ����!�����s�*I����@_&�3,+"x���ȸ�{����ux�QH�!:T�n���g�ܠ!�ss�}�T�գ�>g�����rr��g�fXP��@�罃Cy����G���1�d��wa����/����$Qg_�HL�?Y�T;+	��Ő�$?	'����yqL��/ %&pވ��5!��j�Y�l�}� P�u�5qriV���a���і���*V$���}	�7�%c�q�F`�8�6#�GM�s��%��&x"��3S؄<ݧ�ސFm���>�1'fz���Hxy4�B�ڹo����ce�����D��>�r�ɶ|t�����Wz�Ջ�׏瑤#���ڸ+hT��N�ME�%�ю��E���D��|���q�s�����d.gݩ�v��Y���C/�8���p����Y�C�2P�yt���nƱ����Wޔ��E����U���H�A�D*�[�u��eV�Mi������`�7ޒ������M��$������e�g'�'���j��Ji�|���2�i��<O>��y�Ct�t�J�w�@��?��Ri������h�/��(H��:g�@[	�v;o���ƅB��7ߕ�7>�u	���^���t��cWZ|ݜ:(�4���
aЌH*�9A��y�����Weg犢���cݓ�h��[8"+��t��K�2'Y��g�w]���]n��^��ȹ�e�_�0��S��MK%M8��9�S'�(���E��ˌ��g|�=ml���bY�DN�o�8��Onb�ʥ'�%}�e�r9˔ �N�J�����59e��T>�����o��n�@>���S���t�+���dw)�s���dX���"Q[�C:���jUv/\d�j�JUZ�my��7��-�'��;�'-P�'N7j�2$P=���+|��Q��s�i�q
]�����>���}�sE�ҟVCБ����3ET��.QS6b�	a��nN�IA��R�h8����&gДt3�t=R��z������ޑ��"�ֳ�g24!{�u��M"�J�z��
�G��d(�@!�$Oq]��P^}�e��x��<�!��G	ñ�u[j<���'���!���M�E%B��Z��nݕ|��v0�_�;ɞ����_�J�2y=z��y�\�"��z�s}`PG�Y<P�M�`�f� �ը� �,�9��a�GjL�����}R�]{���o�	Ԇ���A�!6�AU��N]W�3y�����D�'Y�N�����9'�%=F��J��-�]�3�>_�oI��F���g1:A�P9

�9;w�_�h�_�5�9=�d}/)�.� -�Ѓ"�n>[�^�D~��kT�Bн��M���uc���G����C�|@X����jඉr�a�ÙڭC��ھ@x�(HV����;�������N��v;��� ����c��	�B~����wd��}Y[��c�^����ەi�T�n7Ոې���x*Ș-���P|�P)r@t�XW�TҿWǏ���g7�27�S�9����èT$QI@����lL��y�؅�nt�|������֠����ʩD3� �5��z����s�F���A^�R*3t��X c��aĪQ���q��,i�#z�ȥ� �d��6s.Ug�F����̑{�מs�]��ռ����-B������"%jq�(�~F�p�V��!����j�t ��Y_��@�ܳϜ�τk"���M�ңi`��e##qz^ù|�i�PZ�q�O��e2�g�@p���7�7"K�L��"�@[I�iz�$v��i_F�_�a��_6<�%������(��J�Jk�r��� �`��V��)�0)~ln��*\g
��	ٛL���6�Q	��z��|x�ɠ#�B�l���a`��L�%���;cO.�`���˅?�p(�"g�q^�D$K�ar�x���d��E�*9=�C�G�F#&bC�Ǉ&��F�o2�Ѕ��j�<uz2n/\��3PO�-F��(�Z���X���w4Z"yB��Xo�Ԍ|3��Dθ|`�%��¦�l�4�w��21ٔ舭UD.x��a�ٖ���;D��i9����&f�1�Qhd,�IE���YFQ����M�|�k6Ŗ�X�M�Ll�#U��>#� h�����?��`L��Ķ�����޻rC�B�\�{��s��f�61�l�+n��r[���peVw�A��(>g$�%�Gr��t�%e�:$���ۯ�\���cE��,�,z�L2�)T���GK������o�H[��n�^�OXr=�7�@&���xfR��ĴP�D*Kfԃ��ع�F�^����*�:Fv%��>髡88:T�QX]�<X��
�UxVb���I������$���E��q�]�����5��8du"r4fxA.�z7>�r֓��<�fׯ\�'�xL�67��FgD�
���ɑ�Zc��@�pc81�͆EH�uh ϑ�Ny4v2s�q��b�=�z2���C
2��hk�x �G�v.x֐��!����&�<�eP� K���2�����k�7��[��l��M�+BA�-�ù�"Vբ�U^�?�@���I�u�GD�k��yo>��$쓧S���ql���_����ͽ�����%��&���ȸsaG�vM������$i�i :�fH�G�X��h����v��$��׈Iu�iy����r:ܗK���8�_�o� �?��:/,�}�x��D��<�� �	I��C�H��L�$	�8�)���$[Q�D�)XӉ�V=g��۬�n�.L���"�v������SH�q�������v���_����U�&����+�^ߕ�z��|Kh|0r"�������ǒq4���H`��Q���j��{gQJ��m�x_llЉ���M~z��z�~�����5�f-���E���<(#���'���_K�u��� �NOO��X���q���A� U1��1�w������IAfӒ: �)�o����/�YMBS�ln�zR��I�?��OY��𣏤��.[��������y�����?�Sy��w�֝})�V(6yi�Y�r
4�<[��&x��y��Rb^���9���.�^�A��3���9 ��|a8U�< H�g��˯�[o�%�{�{�:9y�����������ܽ,��u��J�ސL�*Gͮ�i���p�<��ASh�	O� ���ӛ�2I�7 <N��<|���(�~B�O�t��|�\NL<�Ƴ��F$v����"���!\0�u�ҤM,k�H��(i�;צC�%}=0�Ը3�2ԧ�@k�� �dE|
������-�#y��u��w_���yW�����o=-e��w�~Ht��_�B��H�z�s5DhD���dE/4�^wD�/�xDe�_%s/���Z� !!� ���C�� �[t��L�	�l�
��1觾�H�-�K��&ovS�x�y���}Q>�?�W_{]�x�)��͛���ɩŪkH*2�s��\�f���D��I�H8j\��1���� ��V���9�78C�9�!Dw�h4W�7���O�X��<&��o������)T�w?��_���?x�&��A�<�gRx��JPZ�8NP<���=|E�\���}w>g`3�=k�w��l���,� d�7�D�A�h���o�����;����z]U�B�������*��au����>��k2�cw�̊UJ�A#�1�vz�+$��"4mZW�'��8��Xށ�O��"%��+`�.����������aNqf��A�#LE�@�}b�th��@�I����k�|�8������r����A��1�,��-�7'�ѳ*"w�! �O�M)^��X<�ٜHH$�M�4����o��o���=�����O>��P}eK��ɱ���f���=75�dĒ�I�ݒ�M�f�;��T�X�(Wu�H�pq�Q6���e`ǵo�8+V���5S<'E�NW��w/�rݾs����3=����\U�>Ǽ���!$M���"��Ɩ�ȏ�7���,���\��� 6Tu�ȍs�iC	<�3���V�ch�S��Fނ��~�g��$d_��?���t��ɾ���QWÁ�2�g�����9��&0�͢�����H��?��(��d>���BJ2M�:7�(D���yK7;�'�$ ǅ>�S>Pm<�{d�5�@$�Q�ý�q;C�읏��k���!��H��JU�텭mik8����*B,�c�+�ɥ��*Ev�c�� ۠�;[(�	`�ya%���h�����P�%_�&��I�2�I`r�/�����}��]��o�^M�By61�b��Q+X�?��F�A������A�iI��4˙���X��$Ќ	�D�ų��.CgMC��^��v�B�f�$Y����sÊ�֜��D��%:�l�
�c��0�C���Ts�޽'��.�=���nG���}��236������ck��=_�3�B}�1��z�d�ZL�őCn����px����ea
�����	����d3.���,W��t�\#���>��^qK�r��������h��)C=�j]y�8CH$ϧ
����ʚz��0Q�Nh��9̇�:�<V7�4��ꉤ|:1X�.Q�u��XI5 p8cB��Q��Ǡʃj�j�&�{�:��jjK�;��D�����Ciu��xC�c�k<�|_?�s��01�?���r(�B'����W1��^3ۻa �n���S��E�D�
�/���-��z���OȓO<%�ٌ	%���X�0P�L�B����Ќ��l�G�WJ�i���91��	PZǵ����g��*�5Ϭ�
z��A��6��3-d�!a_Ŗ"��$o���|�;IJ{�3Td-��E�)�
(�z�+�C�� ND^�5fݟ��)����Dj��#I�$9h���{�@�<+g�Mh�6S�l��FnC����b�9u�C������t��ぜ��t�K�~�B40H#]�ѠO�sT�~�m)��T�;1lZ��pڕYm�1�3P�!\��
��n<��K���4ľ[�e#��t��2(�f�0s�qM�u̍ŉ�8�ȁ\{D�CX�{��D5fkxYC�9�s��H6{}��'��:�I���y*x�x���a�f&�xV�q"���-C'#��B����a��G����7\�^]�o}�yy��y�ꡡ/��)�¹�P玴�������_��?�%U7���Е^��=��5�~-���Z���͗�w��G�d �!�&�B�	��[���?��z^����(v��]5|m�uM�jscM}��R^)��˼SA�UQ�]V��̑3I����m$����p2IZ��%q��<'?(��gq�g���B�×���;�#�W�z�Xf8@��<���>zAN��
$�0F��J�kw�7�H�ZLG�dQ���M]:т�&$�`E0����xOgN�R��A���5m��B�c��wm�&�����r���l�C��}���I�ف=���.���q�٢-�>��BҘef�ɨ?�H�p��� ���eD��cS�2%�c��Iq��
s�����5$�V,tE~�ӟ�����ܺ{�m����K�X\�pI��g���=$��AJE��
s���<��
h�����M/T� &:���/=Sh�^Y[#  �N�3�=r(�YF����JcU����e�ѐ7_{U�ܺM�U�duuU��"�/]�7_y]�dssKCƈ��b&'/#eX$5|Ӟ:��:�ܘ��z�F	�p#��/�@b3bGā��Ki�=��@��V�ǉx�e�� ��"�3����'�g��!t�~�<��㲹�I�.�0c�[��+��(�E���k��(y�z�!Q�g]q
�p�D$5Vޕ41���P�+T������I$�g(pl�:����S"{���b�r�^E+����(�!f��� �Z��"��1T�P��s����L��]<��zd\�MՒ�ļs����=�}μ�|�پvY>?ړW_����J]�y�)���U��?�3y坷(#�}�U��`�W����=�C����<e��IZlQ�[^̥�e&�fDA P�\z(Wk|�������~�ԐiHV,�gEz���^������l�����l���zcM���}P� �l}sG�	� q��[re[��JSܢ��"�'a�4iǺ��g�3%'4(;���7|$�[=5�J^SC����z����t/�!`T)("�B�Rq�t�j�Pa��"9�����W{��4*5����?�KT$�JzD
���7��Ӵ�m/���K�%$�����9ϊ�P}�L�=rqk[~��u)��L�w�`�ʙ�{:���eG�@�g��਄]�|A�O>�^��>��PdL������B�$I���ĩ��&+� y,���#i��Y �!��к�1�A���{1��=���c4A���l�t��ɐ�d�o�X.'0�Z��!X���
���$Nz�L�Kqy!S�Dӱ�jE2=��\!����ꬥu�r��s�>\]��>@K���l��{��ѰA|�@E�z0G�Ӊ���I!�"��X\t�ґ'f$-+��;/�0a�g��8i�3�H���R/H!�0M�3ʻ+A�������%/\�c�P��d��t[m�ՋRѽ�HD��Kz��O˕���ן��+j��᭦�U��ĮD� �����W/4H"�<�ɪ"��^|V.�����y��؞�bB���~C2�yV��6�0��|��g����ޗ�3����#��.�]��c殞~�	���dg}]����������b1�-؆���B�$��4P-˧�;�=���ş�DN��䕗ߐ���I��:����3�،#��ׇJaO7�'B�b�a-@�{P/��}V�����e$����+y��w%W��`.'ø̚H�c�L�m�{��H�=�8^|?Aqqz���A^*����Ђ�p�x�|<4A�C��n���x 9�a|�K,��%���� ��,#G�q���B��po�ռ97u��3�2�V��4�G���~���~��e��}����X}獷9;���z�al%f��������;��@�V5�e�ROW����)��Z���~�3B�����	D
K�..-�C���p��є�_�;l���_R8|I>����ݑ��q�%:��|���j�ʱ�jq2Z��3�:�%w>�����6FhB��1����@y���(�����w�s�u�,���@I�3b#�m'�,rIq`D;�����v���~K6K�|0�I���L�m�ACd���g�2����K���W�����Q�Lm�ٹ���>D� ����3O�3�>�h�*?��/�߽��4�3gl�%�.}��J��>	�!yG/������$���~��;rz֕J�n�FviN�VE�e�k�;�Q������@�ˇ�5p�~����߳��"ۊܪWv��O>&/���r�:ǮK�)m�}iR�r��~���H���ܷ��HR������<����>_�c����\��r�iD� 4����ș�YW>[$�]PR��=���C��L*)%1��Q�0L��R����q��l ��w.�rP�������7����n�!�]+f�%��Ï>�d�I��� �K��)����z�t�ru�"U���Y��b��[�_����k��膚�M=5:�� w��s۝8��=9����ll��/~�s���E�M&���;ҝ��.���k��$ �z�0&�W#&��FDEO�ܐ�}"<䮆��z_�H��Y����!e�'d�	�+\.o#I#�C����=�u�SЧ55]�r�Lm�R~F���ɩ��M?���#+���Xy :h���c8�y�A-7ɉ��5N��׫To�8���*e/��0|Z���%��,r
In�Z��M�C^K�*��uZ1��G̎t�N�Z"�X�0�<��^G�>Ƴ)�ʷ	d��r�9�b��e>�E� �/�_tU��Y�U�����$�B;��qh�A�C��(?v]�qڤ�RD�u#���Ҳ����1�����d_\��pFD�!���3d'��~�|���n����b����s��<��d��	yA"c��n��(�gB��(���>k
��6W�wv,�b��?��|V?l�`��>z].]�*����W���������|��Mf�q�
�4@�|e4�l��&��P��޷�%+��n�W$t��E���r,'�
I[z̦�\>�q��L�q����l�J�=ѐ!(d��Z��[�!O��c$R ߈I�8��:���
��Y�,��ϙ�����T���CIbp��)��H��Μ8����� �9 �Uku=`c�LO�>wV��ք:��x�P�������=6B��n _$2B���OJfzhHeR1u2q�B��q�����b�`�k1��_ �ZY����"؊"��5���J�u�\RQ^����ى�S�t���r�&�э���<PX�0�1�'�!����2 o�ITbl�'��G��L�(��dD&99cqR�\�{bG��4�o�3�)��P�K�2�$���!��$�26�-��"�³��4�h��y�4�t�f]�`�x��\�p�f�`���
��s�7�Q��V�Nt�f<�* �W����ɀQ��r���D������[�Oh���c݄{��IGGKٔ�b��%�W+rt�/�aO�|��vS��pТ����F�N�9���Ej��o
-�����`?L��$1 N'_��= �ӓf�����8z����?�;r��-&u�!�\��.R뤉�{����]R��Y��_�oǜ]3yV5�]��|�A�bW�K�'x�c�������x��٨���ʊ��C�� ����?k��{�nɡ�i�����F��\���E40�`���ڷ�6EY�n:@�,��y��!FO��4+�\�8���_-Oy[C���o�s�=��n/"'�2�3齜� ��P�K�쾌��9�d:��p>�L@�i�ޞ5~�Vפ���f
v>V��c�&��e ��We����U�HX?ML�~�)�����6&�qv;�YĵNv��6�r�&kv��!��X␜��M����{X#ⱖ��1i���$6`�� ��5lx��M򲋱C��emӂN��S�\N֊��BK�d&U�������3�~��64;�.�Jw/��W]�m89��y�M'{��׈4z�!�������BtY_��!
*�����5�3�])��Q�G�&�A�=3�0���zI�'�1�}�$P�ńn�� /��R�5}O��=�Z���PN?�('���>�Ս5pv,F5�	�QM �Ǵ��jT���Z�yV���� 
q�az�
s>=2E��0�,Bn��g�6�rj�*����p�����no��`�1J�1���(`4еUd89�ċ����3V�N@!�bXM"h�Qo®j��Q��Mm�`
����҄�,�_�/r~C'��4kb�05e�+�5dG؁���*����>Tar,C(�'EyV�����У��u�vT5}���N(+�gB��	#`��(]����r2$'ƺ�^�KQC�
�{!�
Z��y/��8H���\HB�?��O���Ġ�採,����=O�;hD��KXgohD�XR�ǋqH�s��Ă�@�5LX�-�eIQ��;�7�h��M]��z��.b§0sl;Ȥ�����u��$+�}�̐BS��\&���I����9/�,SQc��C_�jVV�zw1fR=�{Y5$�z�O��|x]d�
�H_��!�eB[,t�.�#^�T,gĄ0�Ʈ��*/_��7>��#�о���"%D��A����Ϝ�!i(�.W��O[�ǂr�h"!�ԋ_�z�9	o$TxZ'��`2�YP%�b4�o�5	��0g��6�^���9�w�$8�g�VH-�(�VH��)��X��|4����=�I�ٔ���Q�X����wdJB��\U0{��^��{�H�B|�OOx�jǩ�����,=�zx��?r�Ƹ�+����p����u��P���Յ��a�|^#�6�kNf#�#��i�/�:<:�K����v�+���Cq�n�4�c5*ǜ&�e9�BE{|�i�ǡ+߆t�)Aa�m�ˉQ.ͩ����]Z�Ir)q�0�����ր�$x����).9��y &AW�.&vrm�u�f�=����p����o�����Z�	/`(`Z���t���ɔ��s"��,���G�B��cNj�onnHo8e](c��:^��x���<4�36����\,�gMֶ.��7�1��c\�*�A`�}h�|�vd��Ӌ�HD%�ю�LI���W�s���ac��$5@}�}BZ���'�v�l��h_3�1�2.��
�����H�j�6�x�����+y/�^!�2��X����c��X�]Bx3�Nq6��g���r��H	{�H�ҁ��U�v�1��١��Zqn�Xn�	�v�ԑ@W5X����{�M�����!�4�����+"�������-��6��~"������m �g�Z�5ǌ_|�R����sk{K._��Ф!�ש'�}�=� ���h��"���o���t�s�?n
Z�
z͘^���dU�S��S�5�����sm �_%J���s�"A	���J�3��e�5�L�N,<N'Zb�"���/�������Aa$�3E���g"'����D��*��7l���Tlg�96c��*چFDV_�TΒ�N��K��%���2����
[�sֽ�ɕR�X���"�	�q�Q�A�iش��+��>*�H��'��a��|�IMľE4���V�9z����qK����D�����l{��H=*��g�:�	r�QƳb	?R�<O��c��|<5�Ny��#v�������`eֶ9�swkK�z�Q�|���Sa�q���m�Rl4�y&�^[J����@)=�Y�S��j�0��A�V��C���Ŷ�$��;�R���T@t��>#TtC�Ԑ���� �*YE���z$Sӡ�������Y�(k���Y�HnR�`�UO�(��j-��Eﵥ�)T��K<�e�?�jU�$�Rb5r�Y�����gbP�0�O(�1��C�N��ܑ0���6@Ϫ��z/�黙��}t�� ��)�q���ͭ����e�џ��n6P��Lc^ӵڼ�+GZ�T_��QR�s�/^h�zt�3Q��J�9�{W�i�`r������wc����X�z���5Ò�ɛa�a��F$E/Iu��s�cY>�`�x���x݇�p�=���M;óɘ���2"�J��&�0�&�V�M��S��[[����L�F%�WX5P���{̤��t�juԂ���h8aȱ��-E5,u݌+�u�a��:�EL�j�B����F���wN���m��^�3�p��<��6�d�R+_Q��F$LPY�fDh@%r��ݐNL��/��0�X���a@^�c���F��(c���+2�C>�mb��z�B���r�; )�赇�A*�jm[�ب��۳�,7QKtf"�%�q��i���dݧkL��+���g�*Ɣ��sRŘ��֚�)1%~�G g�_�p΄'TϘ�5����"�x�j+l�#��YN�O�)����5���)����Ęl3���f�R���"L.��4�b�1�u`߹$���m��_�3�;�5��dԗ��&�b �^eVN;c9���u�<�R@ ��e2�ׄ�}>4���f;S�H��gadZ"�o�p`cT�ԑa��"�ڥj�碂ت��m�6�2Q_�
k�ժ>��0RC�A�Q�����ܿtx���g�dYΉ�+W���*dևY�B�(�)��F��4o��[r3B�bh��zH��)�AF�b�Oa܃ؒٜ���x��eL/�~.��2�]��	T�f�X������7?���2y�eu�`�<���H�b��v ��ĪB[� s��S��Q6��zƌ���F�"���j�9�s�8�;��c��#�0��)
�����=Pl�c����{���;�󃒷���J�����~O��}al��
�<6;��A����1�O'��/*0��!S�DVc�E�`��(	�`6�˥T���$~����!Q4 >�������P��D�d�ڡo{�٢3*�B˛ �'P��!��3P�K�i�=t�V��D��5�˼?1�S�u�8"��X���2�H;��rn�j�I
�pz�&�{a��!LeE�\%G�ʲ���e�dE["V˩aQ�х����]��Ϥ
�5�9j���QO���k��;	�J�
�:�.�X&��N���� h�d�<�$x���M{(��ƥbId!t��%�<thrя&��le~c?;9��Hg�8��V`1��C��-F�V��R#q�1X&�v8�l^G�g�<(��U�"� � c�
��H�&0@c�Q����0'��l��'�K�z��p����g�#Li�鞔�p��@M6�ES?r�h�����}�b���<�v��O���f��W��Űi_���rHtfm���ӆEU#��1�O�������1o��@�=zW0�:�p��9�?�M�Aq&wu�6ju��X��:��g�&DHt�u����-Vl0��HC�0[r��g>���Vb<&5�ZN�p��ܳ���49�`� ������9h�f�U�=��tΤx��oll��y�^���o���X
h4�u���(g�<5��񙆒�&@41Nb�ķșh��x�!�"JN���D��j)���S���jC&�.���c��o��e� T�A]��a�"���}i��mg{{�!��޾|���G3پ���գh�P���e�8�b62t9���p&��3�0  ��A�s�����g�ݍ�g�s�D?�O��|e�YRb��s	�:����)2�ň���^TbRt6/���\LQ��F��\1{a���s!���2bM�,}��)+���A'�lb�����4��|b�T��۴��<g����Ǯ�\nR=��	�3��M���r��x��l�\��I�T���5j�a���r�Q8�������݉"$}�Pg�Q���&�렅��.d�LӁ؝�A�8"��nx� KOȿ��!%d�[g�t[�I�M�җ���p�l赢����-����=y��	g�`�%���2Է�4�~��{���IhFƒw"�4��BK�Ch��L�"� y9�9	i��`t�6�x����Υ�
�SC���`z��{UP���W�@i�1���G�/����4�L�vp ��;>��}?#��� �<x�2L(����H����\���h���ڦ~n�K�ݫ��@�V�e��{c{��'R�W��K,�C���ޱ�@Z"�}���Xk�5#��0 =b:���ԟ����Ix8 ���1��d��F�.pM�諊<�q ��~!�t���_�q�xxi���;�<��<�I���ċ���3�f]�шK�rd��L]�od�3�<�EP��̝�?(xT��%�	�Xp!��pa@�!�+�l��G�M�rS Ήz$ք�9����j-�ZL4A���!��S�M�+z_y�"�e1P�'yg&�����D��FC�gaU>;:�����Cfv8�.ce�D�22���Cw3��?$��
�[ �2/P��7��w;=Ee"@���m:��RaPv�P`�����V�x���p�	�����������N!3���A���I�e�RlR&�]R��T�8��<�&�y=tC�v���[+�t@�vGN���h��'A�����G�J���\��������w�w)+�#ҽNN�_�_�F)��5��N�9�|�P���挗<U�K�Q*S�����!ǆ9�j�P!Ґ���f#i���"z�̓���ZQ��g��⣗��gf��u:]5�u',{�`�2$	d�;��M��Eh��H���BV#1d~���H��^aRs�T$>�Ѐ��&�����xP�Č���	&��|���7;:9�B�aMqn1��B ���\�k2æ(���qa�r]���Ib�x�$�X��ML�Kf�
_�î����	�ћs��\(m���Z��zM676�6���8ph"Օ52q�"1>�PÀv��]�W/_�b[�_�����?j� C�0��j��G�0��3r�Q����s�ma�o$Tr1ї�3<>5LCW�)��q��T�ixլ���$�e3V���2BA7?�ߚ��n�vW����ݺ%g��\ܢ�Ci�	o/N߆F��D�孕��8U�،a�9��ؐ���H��$X�z���>v��>NON�'�4[WJvp��8AN��1��$����v��H�E��A!��{�4�� ?ª�,���"\����RS�sd�p��yh&#��Y�ы�Y���V
� �A�f�uLb\��Q8��1L�w{gSj�?��/{'���3�J��$��YF/�k2JY��`"?�z2!�f�Q9������P�kbOBu�D�u��d��"̗~�kp�F����, �QLZ��ւ���F���T����ILa:~ۏ���C�c˦��F��%[�`������x�Bu�d��"�9&YN�cU�����!���a"���P*ژOx�z�AI=�I �^he\Xt����c^t�QP!��ee�*�g����Ƿe�~�H'�b�ShD-�����1:10��Us��.!�[�I"'��.{.)l�m�e5x�����A�X����^V��ﰞ!��q��h�`���>�o���TV����r�~[�޻�.=n�\�J��bjjdc��W!�b�Ej�L=c\�%�b����P��3o�S
$���f�>;S�ےK�/������*����z����JC��z�lN&�����c���+�%:�b1�27�Na��&D��<�>a�r΀��A& �,b5�B���=�LĞA�q�m�qQQ�:����惂HulAL�V��!)�5�^���e�� �N_�j�}5���l�+�k���W���5�ԡ��B�m8}�u�)JA5*�F�b��*���P�	1�gn٢o
g���u����DK�Xo��fTĕ�=:��o4"Y��ޖ��6;yI4qcz������j?Ip��,�ʘHB�;1	����H�9�!��3Mqˇ��	Db��H��1�\����q��1�}(�I�q�Tu�keݔ�&�д0��;��T�N#��Y��A�8ʪ�t������,(���6�J�+Ő

I�(���P�D�d�8L��`��w����A=��2X���H���ϝ��Ԡ��ˮ����:{Q [G�� �a�0�	9���P-�q�p�Q$g4IU7�J����$>V�]!LDq�$$M}�����ɧ0�p�dN�yU�.�m�z�%YO��˱" �D`/]�D^Ɍ1���^Cԙ T�3y=�٢�x�ss� �W�V�����Ր��B��obM�nfO,�I�r:�O��8MĂ�NQju.��ryw[�*�]j�	�?��U��إm
Y��f�%��|S:4pH�UgJu��1O9��**Đ���$k���xo���p�#�ya�r�e;@"�zSv�c�%�C�	ʘ����u���ԜJ����Q��T���oc�&BZq��g���� gܘ"Y�>LND7����8�YnF�E��Y�$A[U"d�<�1L�D��9ċ(�a��<[ĒC97�����Ǉ`>�G
h6��2$�M�]��z�I�X�R�r���֭;�/�˲s�2� ���F���5%W$��m_�&��Z� @򿒢��p"ͳ6QSM�(�@�Я�A�cBg�S���8
 ��iئf%F,ε��>�4������t��/���|�s����z��M�\eϺ�&�}E"�������^���M���?��� ���z�x�N�\B��i3���$k4��L�dSV�""�@۰۔bC�(D(���U�����H7�ܪ��yu�*��9�6x����Ԩ��V\eb��xǣA_�P638�q?�)d�;�"'2Иxθ'�/)gg���C�Q%�骬TK�);��ʥ�"��0�#N�jtG�1�{C��9�M�������TY�G{J��Y�{�Cn)��h5Pt�x�hcC�z��jdh�D�m/e��}��	��3_��b�d;Ki..u�3	+�?�ʒ|��B�a4�A8���CTg�:���0&�I`68Cd Tu
���1��&��Nd�ơZ^�N0q��X���>r'��Q���@&Ƶ �lU@b5����^��XbC�a���z�X6�w�a�a��ݎ��>�&9�����>�	^_7��fM�6� ��J>奁�"��8T�Uf��jh���x���F���g:�\�`}Fl6�'q��0Nj�2�Nc�O�`)��=a�$�h�U���2���[ �5)(L .���g��A���@Uk`����-\Ewt�m$�W�,�Mށ$�J�!"d*��q����n�%~S���I��]��L�ՐQ5�]�	�F��,����q`��u(y�+�ϒ��߯��-��yBE;��:g���NZ3N$ݡI�	�l,�3"@�0��Ʉ�b���S����Z���۽���'�E�B�*4"����{l�ueu��fsO��H�о+mw��Hr��GC!�n�<�h����jH,g(t�V���,��	R�3�I���s�"iW���$��xQ��D��b��3���'b�����aB;�@�B=0���Ɍ��s
!�@V��RL��Lꡲ�.��y!�;R�(f�L�_.U���U����T���Z���7�kª�r('�1)��F�aT�����{{-��D7$A�ڮaO�� 	IA���\]C���Zgz�}D����t�"��!d&x&V�2�É���cyf=߱A-A8��6���B�^�3��U<��)���hXsr(���Ո��l$�
��OI21�lw���k�����G.D��`7V=�0���[��hd�S����M�sW�����Gej�Ty �7�� ��أQ�qyAz�w����]]�c9�{�߫�AA%��!�l$�{=�{���I�?�����	�}v��AQ�N���'0�T��Hr�=H�J�6�J�:G9�9���4Шt�q�M�5ۻ;�R$�k�u�q�ly��B��H$�ԙ ?�$+_�|����ݶ�c��cY�ޒg�s]j5T#�Uٕ��(_���2e�0%��sF�?�&��y�Y���駤�sN	0�nv��}ߥ���k��+�x5�d��у]��P�f�(���P���XDru��5����!QT�<uI�FG$IRsf��L��~Q�Q���$�k���˯�������n�Q�y ���ʅ�F4(!Ûp�u`	^lZ�H�xgG��[o���>X&6M,Pϩ�ő�����WP���ޓnw(�n~(>+G00e= كO0��D�Mm*rt�|H��C��y -����9&���:�Q284���m�@ڭ.=�g�#Gw?����#WU��4�*��#H{�TP�W�kT/fC�vq]��G?�<��"?3�,c����4�^�ysϩ�'9a~}��QHޡJq�l2�W�
1����\���(�9�����S��<(J�@bh�G�S�\�Ze���Ed���O�C��H��|�o��f]�P|��@_����OG��*yn2_��cw��`�G��21�٠��C���Rm�^�����|W�b�l����&sB\�V�@&���l e-�pP�c��?a.��k�r2�p4���c]��D�u�%3ck�Ll�?'Wd��!؜�_!��~����^S��mK�D���%�b�J�2o$��G��ĸ��2"n�y�/\�@���� ���o��2�bdc��d^
��"ˌ���J�{��$OcrysC���ɿ�ӗ���]����U+���@~��ȿ�w�^>����� �����,9�J�n�����)��>Ō�]�(�~�	�����mi5�u#X�g�� .�O8�O&��;{>��+����!O�i=�n*d�)��Pf����&S���x���tT21�� �AAM!1�"��@"/��H`�~�+�e�N�%�r/ls�PC�F���e�́�*��\��#;kk��~�9�W.)̮�����J�[ �`����V&�\X�g`d�01���aԌ�(yV�o�g���O~*/|�y+�ц���l�6�
�)$#c�\��Z�����8؅B��(���?�Wt��+�?h�5 �O�ޛ�gcH�f e��i/G����s��D����Ǳ�`#� .��jU�?�4�	�~qA��y݋@�0>��)AٌS"vt��/@�
��<^Wߦ���'�qA�T�C^D�S�s�HM_'N�,�������Q��h�NAϡ^�WY󒲭90N���kΉ�/��RDc��Pґo:<���9�K�6�H<����l'�������Y�����u�������{�&;�4[le��|�{��#� 軛�6$�gn��E��Eҋ��'�~��J��ޘ�w����}ӓ 	 $��@���m������ȹ�	e7X0U��ٹ�g׷9�`������ߵYO�6���sWXߐEz@½������k��_~�&���9���3yu�A�R��\Ds��H�	�?}�<�̳��ͶB���
�C[�+�*��2�3�h�<�Z<��R��(�!��:������I̋Ǣ�q�%lQ�!X]�3��c�W��r�:��lr���Cf��b���ŋ/��{��k�s�QId\ҎE[g�j:�e0s����^��qV����Ǣ�>�\^�]SgS�D&;6J���zO#3?���͙H��,6���Qt'kcԓ#y[�L�˛W��`��SS�,�>��s?)!@#��xr����0�P���P��&3�t��b3ON�Q�}5���B|7��bA\*ck!n�0
Al�p�^:���&�z�d��W�Wm�V�Z������K�m-�C͵�Rh\�t�����p=xn:Q�FU��d��8�@C�
>?6��gQ\�^��9B�+����<S�HTh ��F�4p�� ���u��3�p������+��πD�&x�B�3uM_�Ü|�52�j"�ۣ��%���R�F�
�X(^�`�
Lt�������Ŗ-��0/h���~۶lƦ5k�ꫯ�k=��nl߶U���a�O���B�������?ѩ�_����9I9s%�x�|���K�=�e]�>��K�_��9�T�Գ&�0^�Q#3�i=���-���D���	F�4�DF��+��>��k�$�o�m+6O����5����ַB��kW4���u���<��C�Zg����a��������kZa�����Dz�	R`���X��/��Yk�E�P�V�$�8;��)�[i_��ۜ�!����s�$��ex�i�:l�3��F`������U+%�[+�� D�#�b�J(�{��D@��ʄ&
S:0I���-��.�8�;B�_���r_,X�NQ��p��y���!�w�{�&�t��<�:ׂ���Q��)�u�5�d-1��kx���Q��^�f9FG�竊sa����gŪ�J���v�\��O)�ӻ�֜�bt���@��.�,{��n7U�d����0>?z
��r�����sP�x����~f�����!�u���K���2��'�+�,�����������\�V�]"�|C��u9�ɛsb���ҁ)���!��EkT��G�7�]!9o Q�x`	!�~h'��K?�M=�CVmr��&gB��b��F�����q�0$�gS�.Q���%蚊��lr��e�>��|~� .��ʍ�%D ^������{%�|�_ņ�ˍ4!��ʥ*oeWR�W@���&��$��i�u`��8&8H�����'���*^~���������"�4���J0yB�������dF`_�<��� �������x)����Y9�Y2��'G�Y�LtX���8%;^l{j*��v���ʙ*�-�ϧ�aUֻ�657�)���+�f��w�ǕF�x^<��Ԡ���#*������TY�``�4�����:��HS���*F�����7"��(����K�`IJ�c��?�ں����� RN�Ej�uy6u���$BBE����WQ"��yF��<H���0�MQ���GAC�$ԏI��~x�,_���pA�����J�Z��,ׅO��4��ت�k���j�����Rlׄ EF�$�&�2�u�\|�[ĕ ��֧k��VC������w�	u̩q�'n|pf�0ag]z��6_��%��g���;i����NE��6?;UA�Њy���M�^���,SE��,���$���;��O��ز1�C��Tk�>
s��ؐ�JC���$��̗��//`��+*F�W˒7�^>��}����cɚ����~�S�5e&:�2�"�|Zgp�^��?��M�\2�>�2�`Je���R�֎Y��`�7Ӽ�fC��߰���������[6xU�ًWq��9�1 �3�4���4��@:��m�q��ԂZrh.\�����p�ˣ
�fk[93��#4߳,U|�GZ7i�xtr���4�+�̖*7%?7��v����ƭT��aJ֝Q�9�� �� �@#��;����i(1�R���ck����FA�(�r�J�\*jj��M'S*|��.J2��Á�uz]֢���%� L���"qH�$n�3��ɴ.&������ +{
eO+{�՚'x�>������5��b8چ,��w:�Z����#�7t�@#��|�L��ȩ�G`�v� [)�LN`RZ�ް�փ�5��� }���C�aqAs��vWO0�����I�ƌ�>�ֳxN|�c��h�9�_I���+�n���.���x�a��.�s�?�ek�bzvZ�0�]��{`jrJ��ux`�l\�TG��aK�w�a��r�x�c���y�T�xچ,��W'.�o��El[�LrE`��'�չ	̞��Pޓ�����L�!34"�h�:���ZAD��T� )C�O
�e(a�`E��(�����Z�m8�Lh9���D���F�D�(<�3�;EN�L��Z�R#N�5��lRE\�6#��m�r��z��)����|���١Q�g('�F�������kGL��+8�TϛLhњS�J
N��T�����<�r���	���X�� ��i�P�\Ȧ+KJ@���	Ȉ�Q	�NS���:�9vҨ��s��V�)��/�S6�65��9�����w������yv�t�*��-W5&��Ii��f��I���`��|1*��3-���4"ӾO;�N�΁8�����*IS´d=3�ukik6��4�3�蕆���[�F�	GG���G�3��N�g�W��0�:4]u�4"�n�ʈ�;V��!&�^Lh�=���}�z�.��?��M|v�Z�Cg&�����!9�O�,6�Z�`��<�w_� ���G����M�<oE�.LM�+�n4�{��OQ�C�|�2�� �k1�FI��#�vҚO��OR7Jh4\�����tz��V�+aG�kZ�1�g:�]7Z��� ��\�u�@;
$���#�d
N���ww��<j��=(�F(��BNc�S5�h͂�<�-�#^�1�*LY�oI���� 1�0tͪΓ]�HۓQ�cBi=���|��Wd�A��;��xS�b�"�U�Io���B#)�4c��y�]�I���9��e���֜¤&~Q(�'�u!�\Ef&��Z����k����V`f�#�#��)L��)G�|�n�H�kE0#kIZ�e�ݬ���H������jd����,P&��������	I��)�H�|1mP�]�fF#�w4}��6�˳����#�_5��oz)$>�X�(�е~wf�'x�ϋ������w:F��D��#0C$�?׈�?�q�\}X�����'%�M��O���E�X9���n �&/����_�PÓ�+@���L��$jI�8}��ʌ������L�˶/)I:��6�9��Myf�2�07I2`N���l^/�ө��Ї��7`�l�*�^=#���xA�ޒ
H��[&R���Ԕ�'-ٵ0�&���k;rJ���?�J��4Jt��e-���3iD��SɢV�	�S�'�w�V�}�d�i5�c"�C�
��� �.�<;P�*��b�I�3�f�z�(7�e���+�d��O��69�F��b��Z'�0%!�O3-;L�m���TF�䌑��+�Z�����(���鎙��=���ꍳ=q�"�y���ά�<Y^p�9ž�D�#�4�k��FA�����gc䮯��Kܒt�,?�H��<ˡp�H�
��0.}{�_^��G��pd���ڟ�ZZ#�+�O~�;Q=Q2�|Zּ�4�Q���1�8-,�T�
ŢD"E����gxF����9�{�j8s�ҿ��&�q[:7�@� ��
d$U�U��Z	����PP��z�Y���ާg�����a���*~m4C�qY�l8ϋ-8�1��bN7��Ye���@��P<�
��C���s(	���X�^+�7^Q�2q��V���}�t���lG��9��=��pzN����<\굘a�WB�\I;��P�1�Ab;8Uu��GG`��K���Ij�$B���K�܆3o�HF�����mFǨm�%�N)��Uo�-�E��c���\R�oi*��)�����m&�%����ֶ�kk�ϣƻ7�ա�u�{���_��➩*k}�ԛTH�7�gH�I�C�|C�9HT5Py�6���W���Ĭ�v$��h��V�FA�sċ4��<��k����x����
"�N��?�3.�gZfD��s���2*�fg"5���c(�"��� k������'J���Jn_`�0xɡ��	L��b�BV����%<W�S9�������ݚ��z��F"�X��|	A6��{I�b��d7���d-g���¹5dԾ��8��c�Aʀ��^��";�଄��0�5!mK�'M�]���BL��xrM�Qv�f0�7�ET?#N�����'���Jj�IZSH���1�4t2rXOk�mSW���x�^2ab���m
~oб�MJR��h�p��Q��ik��z��^���O�RcJ&�1��?����	d<#jm6_G��Y�Q����`���gMDD:���y|q�(N\8�Cz*+�������	N�������^1��c\�m�3
�����4R��16s��ٲ���T�����t���(�����.��ޣx�������o�ĉ�*Ud�=�LToqBP����`�j	��"�-�~��7�4۲��n�?��?�E�����|n���*��:һ4"��N�K�V~��zOE2��%��ޕxda#Jն.1��
⍞yz��Ck`p4������<*��J"f(1��g�)I��᱇����������$ZJ�K�E��Df���.��n���(��{�he۠�:I3���f�LU�
��3��B�?������ѹ��10�~-���'Ƒ�u�0�'��ʹsox�իm8�|�hYM���x�|���ˊlX9�lj�%`[v�T�UI�ϔ��y�����4�#;���;kV-CQ,υױP���T� #�U��t��h�D_+[t���ѐ�2���q�������n^�kF�����9\�>�R�!�"�7��+�����?�y����PFeA;��$�� ;�3fp}vN6���M��kd�s�N7�C�{zsf}���0����(4u Xj�Ku�;��l����Io}S���U�n(���4�_�?��w�a�=7k|��`jj��*f�Ζ�*�$��H�<R����մEF+���E���e/r��3�A �΋k��������jD���E{��_��"�(��c̨ڹ�߲u#���i�;2�C���_�p�ެ!W��ѧ����%�h�lI����C`�-�.
�9Ȇ�%9ՙ&�S����S/r=q(x�k٩)0��Α),��ڔ��a�mW�rÅ����y��F6~"�Q[�z��c�j�b=�X-[O7�9��A�@�á8��=fm��F����gհfy?~�<��V�~�YI��JS�P���s���G�p��#��͢!����O�x&<߱s��g/ /?��k������L���I�Z<������Eoڥ��+Th?׋c�66޻
��/��uÊ���^Ƨ��g���\��-���y>�yIu˭:j�e%\bY�b��-xa�<��#ػ� ��/^�\sAe.�Yj](nyO�F�+������e����}@C�������� Q���8�lZ�5��8��-Pv�T������:ܲiJ��s�=�˿�31��j�Pi���},�p@� S���@C�#�y���G�Έ���=�|h�i��z]�8"��u�2J��I )����)u�� ���a3_���r.v�4��8�G��� ���h5�qj&]y�[�˥��0��tb9X���>vv���bp&��^��6��p�#7�f�:&H�bX��#Л���S�aت��<0��7bX͂�{؅"c#���4�b�2�n���\�U~���;�w�`=gdzxfm����.؇�8I?�N	��Z��}H<���W1!��q6n����F
X�t O?��.\�>��K3(�G��W��~�(vmY������)|�����G�$vD�|�-�)���)y8���o�����cd8����F>������M+�bt���Tj�X�|H~�Q�[~q�?����t���I`��<���زa�7�Ոヽc�̔�f(5U�gs���?rc:����8*�,L[^���@����I�6�Ɵ��Gx���di�2Kj2H�	N�����2�'_��M�����d-������s8v�8Ju5���1J�t���5��!�����z�MӍ踿�#�߅�q�\{?`yGz�qwQX5�=Λ�45p)�G��������CT���l�4�:��J�j�@J�u���ݛ]��i�J��7x�(f��Sw��,�H���^`	m�C�q��#jF�)rDQ�$�(y���w0�	#���[�9Gʀ���P6QWY.����	i��6S�ۧj܈��F7F���aH/$�GvV}��QT��Pm�-�z�6/�����ޞG�z|	���x���ś{��G���
�õa��Dp���C���c	lܸ?���q��)Y��bY������<��R0��Ͷb#]Cb�Q���~&#�7��)�Fd;:!���V3;?$=jԵvP��EV�ǖ]��eQ��P��˓���yN�GI�J6�Z	d��bg�����G����Z�Ṋ�y��5v�a�&W\���w֨F�(�ޕmڲ� J�Qj�|fP������4���+�d�T�Rא���pER��� <[k����|C�Զ���Ӛc�nS���w����Ge���K� 1&���x}E�ѽ�<:Z��'����j /B["zfS��aVB�-�P-�Ց�8{��T�pD�(F�R��ŭ`dhX�Gj� �G0ݒ�oT�g����rI#��<�}3vl���4��$.7���"��If�5�3���i�r�s�:�4�QQ�B&bq����e�s|�q�*dC&��)���ؽ�~<��A5J�����贄�9��*րCw�����l<�Q+���ƽ�1Nì537���,ڶb.��?�8��ڡ�|%��o_ǡ3Ө'gqb�޻X;^���k�;[6����S>�T�[|��Q��Y��P
UB�LB;�
X�k *�	����u�W���>fx���ĥ�TA��T ���~r�+�WBl{�1,_5�-ߦ��=�C�.�FJ@9�͐�ۼ�8t
#6�Ɗ��$.��oS��7� w��ܿ���-�lnF*N��Q@zλ��YP(�������?��º��������ch�(iWCS2Ý<v�$���~��'04>���GN��~�'�䳷T��\2a��t|�O����V]�ލ[LQ_��.��DJ���͝�#���7zш��^���H~��m��P�ѨMMM��E'�N�=��%�;y�d̍ATk&�o94784��S��''��u�N���=��q��)��>��>���V�ĩ��pzv%��$�L�j`�/�M8KJO�u��5f�z�(�Y�ٰ��|��f���̐1/�/�q�݄l֮]'g��ӫ�O�=�CGI�ER�R��\�5��~5���]:��⊐Z�3vOmLؗ��y���Oqp@�vd
*��������Wcx�V�>s��k3S�>ç���G/��=��<� V�����p���رI_��%몙C�^�S*"ő�pR�-�\ק��n�����Pa;��7� �J0=yo��1N_���S%l���� ��x�Տ�Cu���{��Y*03��.�<��KG堕d���.�J�M�e�\n~����z�dچ�P���05��ь�2U������<��6��3ظj���X"�a~�

b���Rc� �O�ć�(3�r[J��@z�r�4�dG}���۵����nJ<���b��X�½4�1�� ��<��^lD��M�VM�_��O
���,\��o�%�ILN/`v���;��H ҈�^���o�BWK�heo��(v(�hq�6����QG6���,^}�}�H��"���4nZ��j�����Q:��6f�##��K/��<��,��m��Ol٠�l^>KV��+�5-�H�)q4͒JtT����O`p �󻑑uTЎ-����,ݰ�O;2^M�{V
#�o/?�FG��rG�^��u+14:�m;���%�{I�X%��$�.'����c�1U�*�~��{�g������Д���V�I�R(�!oc-����lm-)F��}p;yr��!�",ZY�2��,�1/���/��!����٨�k����)��ġx����bX2B`b�������RE����i��ׯ>	��/��}��1
�*^��q[�][y~#*�2�|m�~�:~��xP���<��۴��6`l��)OyG8W��~Q����#*��'�Έ��8E"KjNu �R&��bz4q͂����M/�q�ߥ+��]�������j�_��	E�>��<sjD�]��غ7���"�2��+��Nʒj��q��Fs
�o�T:���mٸ���n1�:�d[�]2��atdH=��B�\��BS�Ɔ�JW�Mt��J�� �i^<eđ�з�#�h �a����Q\:��v>��hFR��x�
	���F�:�m��,���ו�&�?74U�s��d��@���QV]��v������Bs/fw�hĊ)��ƦQ?��m:70��jc+��(�G~s�q�^�nY�=�<����9;����Ǯ�%�����{��4�����K��'��uc�^�*�[&7$�i�UM�!�)�5�������㢚����#���*I�<J���l��RW֍͐�!�i*�A`�hIchT	7�(�ob��Q<��:l߾�V��ĥ���5Y��eTY�­#�[��q�r�������'UG'-���jꙈ�m+:Z�/�� �پ�pa�wm��Ƕc�%
��/J��cf���'�}���%��v[Z���(KZ��{#S0ST=I��Ȳ���]}�5}0�����B��2�� _��5dMFA_$��ɺ)P��Ӛ,�%���vfF�rX52 ��+�u��9cb��(X��AN��J
�ھq-֌���[q�ֵ:�I#P��q��u?s_�8��g� l��<���}�5Iw8��G詌�f�L��ܝb|��+xo�粑7c�� +�S��̊q:}��l��D U�rU1�:A:46���Mٰ��׮^���K�+�v��@;)�_֡*p>����]��ZZ��P�M�	V���;!�_�<�_���x�gqϊ���|L�~_��� +�a�+w��y6�gf��;�x�g��7I$�/� idMN�1�3�Y~]>CF�g�h��,N<�i�Rv��b�ⱊ�����?�۶��G���|M�U*�Le]�&�T�,S�Aɐ.E��2
K�x�����}@#@"W?=p�&��M'�L0#yW����<�P=����P��<�5ӚY2PQzVC�Z��\���.�L�۰f|����bz�����N5���d�����ۚG�.g)�ڲ��K�pյ�]Z���hT8�?D�EVۥ�<���u��W=����hՄ�!���{��vazz�{g�~y-�����;�*l�]�`�� ���w����0RH!?$iL!T4=�ܿ�lݺ	{��;��ko}���y+�F�y$��00I ��C��{�=J�ł(E�*b~��;����عc5���3�+����>: )���u�n��<��S�H"�����!<�k�����Ө��اl�k�5<,]���Vu� e��z�[=��4������6���<,)J?~zvm����lϲ�L�rMt�V� Q����B~���9��G��[��#���U�ٙ��m���R塞�_^���H�F�2^�����[]�I"�!�=�IbZ�������`�.]g��H������HJQ�^��d���S-X�Q�hpF�ܕY|�O����Q��	�J����B�N˥*���,sz�}9Z�Ib���i��ڒ�m:uL#�k$��w���e�#H��k��S*nN�F��d�3�L-M֚��ဟ�5�@�ܗ�	�O�Y�p)5�r����Q��%O2E�p�ª��v8$�IG�����{�o�'/^�gǎȦo�<����a\�t���̞�a��qtҒ.H��'�Kw]]� �aIf)^���İd�����x֌��䄉�0���n��CRq"��#G�l�ɒ���s�<u3ծ
3���s	C�(�K�;��hi���p��S�*�@F~�z���<}ICι����s�HR�����3�Ab(�ͬKؽ�76��y1"�=C(�a�|q׮U�ɖ����[�a�,���]�n���R�����	���py�/N���Y��8&ϩ�M(EG�n]k%��<�VX��S,B8	x�&M�r�����LE�<'���r�2l'�
ƙ쀦B-���E�TZx��q���&�q���,���XT-��'��۶>�!u�)Ϡ�I����*�<u$��ߐ}��H*,�2 5$���5TJ%�б~�v@�F��S�<�49�=����{��g�s$��$�\���0������I��ֈ��e���d�E��H�w����)	�Ed3,��UP��lղ1�KV�}�=��X���-v��J��)��`��7�nrH�;�K��#9hG���8?]�ΣC����D���
��p�(�$��P	*�Q��I�qP\�BYdݢ��"{�31ͪ!I���4ay;	�#��B�h�P�J%�ɓJP�&&v�Rjjî�q��r 3�y�w���������L�u$M��lT'�(AQ]�S���U����|�Y��|�NU�|~z9�u~V����}ҁL�r����#]>}����r ;~WE��jG��i��|�\&'��,���~�dg��*yybĨ��<�����I�<uNɗ|y�	14,�W*UI�SZ�$�Q�N��^���ǿ׉'r��<Ӣ��=��F��mU�m��e8/�t�b���̛���Ē;�tɄ��Z��d�'����gO%=��C��=�G:����������C�|�r�tu�ܮJTt'�*V�*�D~��_��y I��j]@�j�eޗ���]6�=m��)�$����U8ue��~����(�]W���`C�E<)��%���>���/_G��a&7���>#]	�AH��>��C��̥���+3-����lL"[��Bm�r��Ij���U�he��b�y�$�I����*a���Q`I_���u����Z�����b�\�a�*5}�A�T�JzC��'M�=��IT"���Q���`3�tmi(�MET2kʑh�`�!��-h�3Bf�����D�2l��H�L���"9<�ʌN'SZ+��&N!����-�K�kֵV��7'
/ɩ�
���1%�nSC9L+\@)���if ��Z�p�Vc��q"�2�5���R-l^?�m۶����2^V��\aebA�/C�P�NV�g V2 �,Y*)zW��!�V��+{;�O��h�]��������lOB5�˥��#'��%,�$6"nZ�����D	1�m!%(��&����J:82;�2��q���p:1��<�U+F0PK�á�g�������J�-�v�#�ˋE6u�SW&�7��9�.�0�Ů�����µӒ��t1t�k@KT�jB
4Q�T�A��je$%dX�|PS�T[���c�8�.�ϊ�x72��u*��Z�� �q������<9�����h�v[ۧr����j���߭�Bn4�]�ߡfT����ע�X1��P$k��Bʾs��+��%ge&�B$�x����]hV�l����!I	0]�^����T��hxO�v'\��{�����>Cz�T&�+�-Q^�\��]�Ke��D�*�K�(M�03;��1lC����jsA"B1&�F�$Nab�*i�lf1J��Yq**�~���eٿ�0�1����c��_�kr��>N�!/`�ƍعm5�}�-]�����s�h�!=}�(e�|䵚59t�y�Z�Ͼ��߄��ރg���B�9��2�g4�Ȅ3tfݺ����a�\���X�T+
��ī��f���c|��R�Ĕ���a��Y�F��#��F��w�_��ޅX�T��|����w���u��Q���|�AS5\|� �%�|o������#��d
$x4�$!�*ݨZ�ƀ�fRH^�1��E�ne�S�}�1�V��h���xw�g���5���*o��zUi����r:�����0q}��/�`F����_��a�"�#S?��U�E}����p��: �N�FF�(�qT�KU"��+�I���=x��{�c�AO�"w����[��S�d}h���q<A^c�P/���ؾy�±O�;���[8~iN�mAS���C״N�ƪq7\�I���{��Hz�lN#Tv�8�Z�Ğ���o��'شZ���F*k�F����x�w���qez)R(�A$�oO�y�>�K�v
�z�m����gפ^B>3Lo�Z�\T��q�;�M�-����e�St��g��8L(�I�����xL�j쏲D��7��j1,�v���~�:>ڻ_�9e��2�y�!|�G�~�V�1�zc����H���H+�T�(����U�/
���E\6��neV��p�"��'ƒ�_��0���*�N�<w6w�܆��䫖��q,�>mk���*W�*�u%�X�tV�Y�R��U�مy\�t��D!�h�F.��!'��H�ۑP����hJ��̔Z`�CU@Gջff%tR ��g��[`��ЮaêQ�ں��o�#��G�HI���+V���U+1��}���	,̋׬�=��{uxl�}��mQƹ�5|��W���19$�0�4�L�L�T�c`��3�q�o�D�ϖm�k�f������َ��Ƃx�
:'%����[2�߾�N\��D�Ǻkp��mx���p���jC<p|j�x���=V��f�I��<���cJz*�Dxu�<'� �� )�}�6$��7pir�C#U��~�<Ɨ���'U;yt|)FGǰ|�vܷ�cE	�KX��er�$Ne�Rc6��%	�nȺ\�����1w-��iq�t��F:OQ���5Y�&�}b�D�0(�x���I�  �5IDAT><rV�6�^��l������~�֍���˒�b���ز}�,Ӛӵ�)1���7�C�&�?'xY�RϞPU� @�V��Њt˭�����/Z0���7���&}+��s6��t���8Vuf&r�i�Vj�'����9+R:#At)ѩ$Z)�˸:1)�4�l����g�޾S���Nt$\��w]I+(�X��������M*�eQaO��2G#���z/a'w僷K(����{��Ƃ���檒ߕ0�Ϡ ���MX>8���ΦxQ{�<���كq9�AV>G����f��᫸pmB�Y��qO��0j*�H{�&��{N3�w7__��1�Q����%�{��ؽ{+X�:;��ׯ+K���$�Z%�惻6#�p��Ɩ-��#cKU��)��38~�2^���8~yJ9VՈX� 7�f �w��0�(^P�hՀ�;]Õz���&Ƙ!�\i����|u�W��·��K�9$��Ɠ;�аI�*v�rWǗ�/�-�T����FVig�$��QlM�����#n��� �9��lSs#eg��Ä��+ܟ�qj����W�][1$���S��k||1�q�uK��˟<����(�"�g�܎vw�D[�c����켜�9|q�>��w��|��N�3�=7D�u��9���ix�f�[��}���oqh~/r��m74#�&[��fg�N/�1�,ґ��AړCޕ�gR�V�N_Z���X7��x�V�X���Y�g��]W�(I9t^�(��`�dm���6�jX��E���z7�3J�C�2��M���C�S��ё"�K�L���_~v	���&�g0>�Ó��#�")�K�G�����k��%� �u��5|�ɧ8��y\�0���f�ˌ�U�\�(�Ջ���@Ԉxv%­�.�Z�'���'F�x�-�lĞG��hg������=���ĆM����>��Da�#Q��ڰZ�G�W�BS6��������<��r�&K�!r�9Rf�,�(7����M��nߋf@#�m*�-a��.�O~�����T���7>�?��.͇ȟ��T���5/(��'��T^�t�N]��}��ȱ��t}s�6J]I�d/��3#�+�!a�A����M[�B�Ȓ�k�zx�	�,	�F'n��H��R��D�$�`�z��1|�?j��*gy��U�|�o�9@"���	*$�p���'���ǟI�5�-�N�+QԀN87�YCR�t��^#Ro+"�<i��񁏣���1�7"�o̹�}ˇ���L��3�w�� �yQ�!1�#��~���P�"?���oǂx��IRڗ҆�+)�o��!��}>:rN����$�شv96�\n���k}��'T<�-�"���ٚ��n��l����`���qͶ��G$�|Õ�����?�o>�b4P��qi��\q;���ؼc+2r �-�<3��G�����̅�h��Ȩfj��!��ɟ�,�aop+�%���n�"�	�"��Ơ�o�e��(/��_��7?´��l�S�a0?�c#ȋ� �S~d�2�=�����ȉ����D� ���=�-_������$3�k6j�g�n���w�Ϭ���P6�H�[�f+�m�tdZ�%�`�AL���f��4��3W17_���"ʍ���NL��ԥ	��� ~uJ��<�}h�-,�##S�ɟ�3Sǘ��n-�z��o 2�E)mJϏ��smU�
$5Ob���BR X���+��c~��s`��"�F�s`I\:;��'������c�JyQWI�I5H ���RZ"򻊿P����9U]k 3�c����֔|-��Y��=����H8�޷��/WhѠ�#�9���P%ea��5��/�/���B(^#h{,)0����kQ�E_�j%��g/�z�W��0�{x���������%T��oJI>�99s�6>�\��YHMti�۱��Ƿ\����x�V�%��X)'/���i�᯾Ċ�2T�M�%�����W����b��gqqj���	ސ_W&JP�h�ک0�R�FU�FEE
k�Z��E��yq0��j���4f����7��ϖ�60�
2��JH?U�\)�/�$��"�"ݜ�Կ{� ^��+;?�f��BnX�9Z�wr0"�xx�,mpe��ݚz��ڈ7x�>Қ�^9�=;�d�AS�/�,���0��;'����3b�F�����o��W'.�T���p�ȸ!{�0_���¼�,�AZe:�L�����E���[��!�b'��p��F������C�Ƈ-��K�Bq@�9��B�+EؑhchI�W'��ۿ}.���� �$]��!�@�����i#?�сl	R@�p6.��?S���1�:���|��ۙ�h�a��<vn�F���P�A�#����n�o�:�I���b=�9���������'��RsY�t�:�;"D����#�BF�?ɿ1$�j��V�[�O�}��|�Zl�+�Co�+��DF��q��Χ�/�zMrK���H贬������³G�:�[���U4$z]�H�SCs႒�h�'�"���-��/^�������{�uԿ����'��$O��K�564$�uUs��@^%M��R/:���?�L��tu<�����КS^~[��"8����ha�zX�|3�����_���ʞr�K4��^-aP��FW�Pԁ+,ZV|��������sK9����%#�$P����!�)Y�NI��o�^�<��z��c:��|��{����K3�%4��ƆPC��0���Q���ߧ)��8k]z��T�v\"&:�8�J[B��"���8r�dD����1j9Iɗi
��(�!N�U1Zءå�3Ts�}[���dO��fp���8K_� 	0ʔ��ZCl����uF���]"/>�3����-|�@�V��;_�����T4��Ϳ%�R��a�e�H`s�xO�w�+Rd�Z��o�f�Q�˿�Lr�.�Q��բ��=�%d��=�*�D�hN�ʫ��<�/$���f,��r8ONLcÚQE�������s��_�+�B�BA'wU�)4l�ʪNlC<f������솧$GL::Imr�z�><tZ��	�ڸq5�._�t��,�ԅk�r�F����~E1�7�����N�fE����H�ͣDh��˨1�mҨ#��RRe�(ő�Yi�S�_����L�� �m��ǰ�iYD���`x0�X����y�]�D=ۖ�o���Ϋ	#�͹����r��5��	Հ	���`�,2��`�V4�>M��<+j�,l�?�	ګ�׫It�J���?��G{���X����S�[�&��e�J���)�����FF�PC^�qq��޼� '�8���AN�#�~-4�7_{�B�I���tԶ|U1N�@� 枫4��e0U�`������g�rqW�\Ú����g�H&g8`
#��?�)��ߤS̅�:�RiA��'&;x���"�:��ZH�Ϡ^�ۂz�W��R/&��=��2����-�o^���"� {5���H�����bf3R�����(bݦ�y{�����f�dF�#��ݏK��eyoXg�������KU��l)6�5L�7�Ϗ�Z����Kx��w��w���<y�|r��^�D��dvLk-��b�
!�u	t\E;�s'��?��K��/࡝W�C,C��e#h�J�|ؼa��g?��b߷��Z���;�ĥ��!�Q�� ��_|���
��^�݅��Z����+WqF6����X'i��w+�;4��<�+�)a��rt	������G�k�MMyC�d�E�ʼvh~��^�]�0�8x�%��Tc%��Dsq�O�M��3)G����|W�(О@*;����#<��3�[7�~3ق���Y��X�mVm�Oi�_��f���r�YI-��O�~���Byni�qkt�=�[xa�Q3�����pmv^�ƭ�%��5K�� �F�s�t8�Z���S�Ia&�u�����Ζ,����Q����&�o�����W�W�p��T�=��"�
�������{�7��؀�=l&�����L��Dts�G�E(�0��kʨ��N���,����D;ˮŦl�F�0N�f�7i$� �+m| )DyvZ��>���MH����UB�Psфx[�x���-F��w��.B��6�A%b��>��q��*m�+�D-�JEJZ�5�>�S�ѼB�]�\�Hs�99�/_�91")��3��U0���.^T�V��!��>������WpM��(�Y6��GuJW�PH�DYɶ�=E�%�͏`t����ӝnS���r��2�Q�K��]�E,	I˘���6����h7�8M��n��gj8|�����c��!�)�h�%�$�ZY�� UO�15�V
�H��𚘺V�5N�$�+v3smL�("f��	�������Q3���#S\6�=Q����1r�|���ݻi-�F���]U���"�9�j4I4Fâ�!�g�/���"{grjRɽ��w)�ʕ&�m�tg�`�;VoDs��7J��x1�Bk"�A�r#ҳ||o�hDh t�Q�H�E�Ad_��瀰��D�ۅJ� 3A5�"%���14�S��"_����G�l���<�Ӄƒ@�UJW��PC�bXw\��K�|���2�u����h��`V���ǈDC�zR��*-� ��]�m��*�_����D>'az$��Rj%ص�\�r����n�uq9��q���p��U�]{K%��J�!kҪ*��
H'}e�g*���c ^1lJ$����JUrvY�C_ũ�b�sf &�҂�c�or�ָťD�mr٦uib���_{�ސ�2�T�:�T��~�k�(���(� ��U��ɛ�����ԌD���<�����Y��ou�N�-�خT�Û��r�߫3e\~�C�?�U��K%4�m�}�z1m6�����YҨ)r�P��F��ƕ^#i�ؕV4���>Cr�x��>ʭ,����M.�������f5�DGk$Qz��%����Q\h�*K�1=5�ED��q)l��U�g�ޭE���.���K�Oubr3�%�� E�39�u"3M�'��+��G>�U���LUҤ\�,cZҠPٰȼ�Q^�Ћk��.��4�> �ԗ�N�~�
��8�]�:ZV�ʭ<Z�ؿ�Q�s�?#W:�bn��_�Ԗ#�G;�p-lԫ��\�0ns��m��(6-�Gg�f��#��h[�Ǟ,qsq�dU�Kᐞ�	-�|��W�K�l�y����YhN%���F��E����~yv*�wswڄ�f�]�V�S�s�����5o�k�h)�ͪ~O;O�b��9T��N������*���D�_q*8i��� Ĺ�e�-L�geQ�3�l�hF���%�jMz�&�mc$�z��9�'̆���f�?E�f�	#v���X�/�Q�"����9�ۯ�w��ãs�c"����P��MzԈ �A����ٙ��}��F>��l��׮�^�(y�4"	�[�Fr���l���wl��-��g�8v�$�=�c'.`���^�!6��B�<y�U�V�'��'xl�R�oT�%�^��W���}k��5"	c�L�0��)2!9'!�K�.�DB_?�#��%�x=/X$�P}Ԅz�L���k�	=�%Щ�Ʈ��#�EGŦ�r���g��U���s���G{:�2���u�9{'Zu�7qB�ґM��MX|����*u�ԑܠpx#��h�4��U\�ʚٴ���0�dc���w�(]���U9Y,)L���:�V�#]��AOj�P"Y�M�H����Lѓ�Pb&Z0�����vM	m5[�1�?W�pR���f��=��f�Hρ?��)��ϕ��T�Gd)�8c˴�uM�R�T��cGIf/�A�����q��6�n�������{ME���o7�Q��7z�Mg̻�8KB�\�����2o��&Q(��{�<���g�
d�c����w�����P}��_��U������4��'�|�5j�0�j5�I�
���s��`��?}�)������Y�h�\�v �uC\y�i�f,�1ܤ���D�M̟봺�_ᰞ�:����7�hM�_���Hg�G���^JŤYDN��e�^�}:V��1�������_̑[�~��.U����A�H�-ҎJ>W��U']z�3^]u]3��|�-��e��ջ�ԁ^�~��z�<?e���m?�S����J��B1��M�6��L�ȶꪈ�����%	j:F/��}E�r�X(�K�c�_����-�+d�5�V_0�|�P�t�B{H|G�m�o�G��_�g��=@u���/��Rd�5��K0�'SH��� 
����Tԛ��dV�I+z��b��M�o�i�hDn�������_�.%�1�ә���۬g
c�.�|��S���-�w��X6<�zeAd�$�ն���$<����쏰v�2���^��|��d��t�������������eX5`��#�h»����E�E�kC�H2x�F���i�Y��}����0�dD�0|�m"�I���!P����%�׋taL�}O�����ЀqL$Å�=SP�=�z44r�i����(��epw��·���)��e��L�x��4�rd�:G���kZ�����^YH����n��q�� �N�o�p����s �Вv��SA�D_6[5s�9*�h�Է�R��V�7hCgC�;�zS?_72m����dV����Q0�\��֗KG����t���679Ӣc��7�|�X��jv�/�db|�5���vC+�Z�q�஢�m� ����~Z�A�6�$�SЛ\���M��gϨ��Db��_I�X!�H.�ІY�h���w��虔�fr��Ԉ$���+J���S�b�h��Wd
(�h&ӊp[ gQ���\�=�]�޽{?ދ_JTrv����MM����=g�����;��u�T�H1��W"�N	�X_��(r��a7�K"�ݚ	On6>+���v��h���%{�{1�M�x����ƸV��^�&���[��s��yB��M�L�x�/]Xn?��^��^����Y���������o|����8҆��Āt�V��|F�gx=,9���{�3r��y���R���b:D.W�ֿVQ�o���8��eQ��WI���{�t������q�P�����8��7ܥ.�OD]�C�ں�83�q�=�{�O�g�/�.��N�ĥk3yo��m�J�_�CVN���Q���4_~�ͽ8~u�L�(��骎⟽2�U����TQ���1�%�n�lT��iŢ,X��!�N�i��l]'��>#�^A�����a��m�w5�y:��t�.�w�A]�)�k��>6�'��x�. 6[l�k���7k b@�ۦ�n�g�^�Cux���v�!�z5[Wq����hn�N��mD��yF�.���~�R&	m��5���{��̋�)~ޑ�S�ׯ���������a3��[���[�� �[�|��\�0�ͪ
I�X�$���!�q��=�Bۙ�lV��KƖ�/� ��W
��2���s���!\�����8d��w疍x���f���y����'�Pޑ_���j�f#X�D�4��˗�zh���܂D��(Ƀ�B��҄�p�U����5�e�i��O�m�B��o��!�ۍ�h8�WcCb7��_�g7�}8-�[�n���?��$�kd�\�D�:;1�������-�4�.�xq��m����Z�~�1��D��ܡ��<�U�+���z{�3�`�;C�9� ��^�����r��Ư�=�~���Z��g�@��X��nз9ޞ�',�����M�����x#�����^���W��p2�0'O��b|l�ּr���l~��ۘ���h�N�F�n4j+����#زn	^|�I%qI���Cۑ�%�y�u8qU�\��󓘗���ꈸ:�@uB��ML�!q&bqb�x�q���EtԀ8�Z��s�î&,�a��N��FΌ���۟�U�o,n&1�o.5�{v�צ-mZ˶�m��SO�\~�\o���_|��9z�u�$�tsX�^���s�QtӲ�CjjZ����!��5���W������"Cx}2�f��-/ƉD&]v�<������I�����[�5�����m��g;JF�����N��~E�y�*�I&Q�51�Mc�R��/���)d�V�E,��45D8��N�
����q�Rf��^�~��.%}���0�B�zG�_�X!����'� 5>�VP@�y���z~^�a��Ȍ���&b�o�w�ҹ.H�y�Y��=3r��e��^@��&�7�]�Ⱦn���C���	;-Fs]���
�+NG�A��Y=��h)�=�*o�ݟ�bRh�o{��Σ�үk�oۥ�R��{]�e�;��ȴo�S�����C�_�oG&̉!�^\����e�:�����=�5�K��̢{C[��V�o����m^�]MxC�	�[d��#�8��3?Z!�8�ʕ�uq�;L��N�K'��(%����nE:��j�Cl�O_��/^~O���[����w�yǎ���`c錌�"��'k�^�ZE�k�r�:�.�����zoJL�g6�V�����f��zu�^�bPhi�b����Rg;zc�_}���~��z݆ȹ��t��,���!m����d��a�/ډ��ޣ�."��+�~���p!í=߭O�Ϥ��v�"5.Y">D�?ꙩ^:f�Υo�+���@�Y��g" 
�š�z6E��K}-S�[�7��=O`ɂlty�Q���ת�	Fn��!����݋n�苯��!���L�3٬Nd�.�[Ȅ�N�\���p��[�%��dP�D���V�񃍶2Z�KJ�S���-ƥ� ���+11?�D*-?�B����9����5�� ��ɇ0.7�{�NI|���܌��1<M��R�cD+�gW����NE
3�$$ub�^�˃�X��T�#�Y�(S�D��|jJ�i�׷!���l��������k
�	�����4I�\,��RH��z�F�?n�����e���V��
v�Z�̗��Z[�M�(@g7�*+�¶(�<:a`('����t"3a����l���ꎝJ�!)�gH�Zo7qL���T�"N��᳡Qh�KÎyoJ�r\���� U�E��~�&Փ�$�#�Y�RGϑ���g�Kڊ/r�V˱*c��ѝ�eZ��n<!�^;T��Z�k����F���Z_��&������t�)��i4K�f	]�(B7 �6���V��{K�=�l�tۊ5��)�4T�����M�6�Yl�\'1��ִ�}�5��\1�݁�x��cdmLrd�E�7H�!g���>�bڌ��t�7�����.���r^꜀:�._�V���~�W��SO=�5�ى9�id
è�	>}	�)QJUY̔�f����*����&^ܳ͠���+��g����X�5$�s���륊&�ںg���8��,#�^����Au��.�7���rLW�b`�`��p���ƙ�{"�ϻu�{�ޢ�RÞ�tj�X�R��i�bs��-}`<L�xJ�D��@��;���}�%9�����0�c�Eߵ�$?N�,�ƥE�n�ͮh1F��R�rS�Uއr���)���P�@!��u��f���(w�t}�a��5��1h�v]E��!Y�M���(t�R��.��Q/r��\����wd�ut�y�V�k��l�c��-��3hg�p%Ɋ�F]��/���eR�"��z8y����T:�Ÿ~��:�m؛Q�`���!����;"V����Q�������f 5�[o�u�׊Eƽ�=�m��G{���:��C-���G��:�j5�Y���He�MQ�)�7�}�J?x�Q��Б���ߦx��dY���gQ�_�˩��5HXx��,;W�p�]{0������/g�/%���{��e!֒/���nQh�}�O=�����_r|Q��E/n2�}��M[71A>�l�����	���!�x�yO��Dh�"��0sS=�Aĺ�=q!�J~�h��"��۠k���E�D����V�k9���:{�gD!�A\����5D��H%��ד%#�ߨ�k5U��o�)�$���l'S��߇j�A���zӯ���â�S���b����N�~�� u���T�6�ȍ��G�A:H��H�5�t�}�F�9�������	`�����������o���q��R׮]W	CO��	L��O��;Y��`�C�`|`D"n�4��l�.��ޒ0H�fNR���l��HJ���?��6&������C�$������{hQn��)����?"�m
�Mp5OW�qHPg�M�a��"S�Ո�I^����^�vIL��	?r��D���yC�����cmH	����h>9J���hPy
#9`>Ѵr�C��&Ֆ�̩hzxn�h4�𓦱�o�C��N��#�H)L���sTޑw��]$@~Õd���E�S
>IڢL��,�L��؁�w����C�$��qQ���C�@Y�H��%=�@���ѸeQ���*��������=�.g@��Xۥ��CϤ�D^vr�!褴�=SN�mŞ�ޜg���I_�J����b��C��:�I��sa�@�q�\�Z���-�����F�An�Z#���<�/q��$�u�	�E�ʬ,�P(]��E͞&�g�{���^�l��yȾ����̎m�3l6�&�$� � 
��J�teV�����{��^��,� �g�:�beeFz��{���N��Ә�
����ܔ�8���Ӱ�ޓ��UYY[��:.�	R(RR͎�	.ߔ�@�r�"�΅�.�����p��Oz�N��������3rt߬�U�4�E��q��C�T��)Dl9.�p��e�X��X���pā	M9/IK�	��HǖL�ɕ���6�<�:�<��qyc�+3�Kz�������v�4��7�j��J����iXBFv�^|fxa�mh�GXaHU��A�H&�M�&��\���aF�uͨϱ�&��Df���rtd�tIN�|H�P|~N�~�7�6k��H�,74佶���!�>���{��%2?�ս��3���޹��WeX�-�f�!�{���v��`����х�yN���ɨ�`~0v�)��rݨ�um����ŽZDIM��w�����*c��N�_��wH��ϫby_��w��!����Z�E�v�*����F��kj_cJ$�$c̷ 䄺�Q��0�K)FN..ݕ���|�޻�0W�cǎ�����������eQ����S)U�٨�1�x9�^d�f����ߓ;�/��û�
�3O=�ƥ�_]��VLZF�ɘ���0L�6�	)S�M�!�kߗ>��`�x|o:o��l��`�Yx\7v���YX��q�P&�����
�,\}|�l�=R!:��KH��
#�ɪW��rt��/�C�x7�-J�Wckv�:�������vU�U�܊��	|B���c�\�2`��	�I�N�-��WQ����ɟ}���8B�TȪ�J_��?�Z�?\�H���Ln��$[̓\�א��������Yyh�NUĨL$�#OÛ��||gI:�]U�y&:�`~�7�-�8�D�{�X��1Eb�6��KC�{�M	�5ٹsJ>�K4r��o�S�5`^�U�	;R�o�#���#gO��#��x���7����^�7>�A_�3���w���s^�����y=��z"����C��I"$ɒ�æ�x�26=�hc]�_q�ڍu��/������Q*j,�rд��]�<"���@�`��C"Q7��֔7V1o�\���֪̞������X�"���6g���2C����"�c�p���+��O��u��਴|kʽ^b�.P��дMJ�T!��޶��٦HҎOh(�ݮ������>,{��Է6%����V�q�xiz��������%:L�br=�=�́l��MB��%��k\*d�\dSX�Y�Ò�ֶ�}$�gd�>�b&���|t리O�x�0�b6�}s�2�^F�R�ǳɫ�'��>�����G�<����/?kik ��-J[�}߁��;4-�?~Z�x�=�q��cA�����PjG�8
i�]k��4�5�D�=�����svR��O�*�z�Iy�ݫ����I[=Mw��oC�=�[��_K��:Io����n��<�����އ�Zs��z�d�2���Ҥ��O��?�k����2���ͬNAW)KYHa��. �E���=�X�Y4詵�߻% ���.�vKi77�n�'������ӐH�ʨ�
�M��W�e9��T��(����h,�Mz�0�02�?(W��NJ���p��AO*��lA�c��kYu��jjQ�i���K���>�S�,�z&O�k�$��èV���_��/�q$�?���������7Ԏht<��y�7yZ&c� ��8I밧�z�.ݔ�������mJ)����*��7_��^��|��?Hو���:K���η^�}�~O6UX~��
�һ^��ݽ��@ٺO��.�¿��G2�k��I�U���+��O�w���s3	1t
�gj�%����[�=�apF:���ȏ�K=��|�+'�_ϿDoxv��J�e7���U�������H�}��0J;2�"��N�zX���Srd����n1O��g��{77�G������ٽ{ABUd��ɦ��<sVS���?���HAC� �")K�"����ߥ���LZ,I���|�v��kqI�dmJ����OW�4m���S !�!1:�Se��KC�G��Lf��u1^5�.@���z�J�*��
e�X���ş�|�"�
8�آ��ߺ(?}�u=dj)�Re����p9�����bE���<y���ݚ�]�%�~�UY�j��#�?�X�b���]'�uيF~p�2��P|��^V?�I�n��	/$�rd��R�P��@^I6����v�S�0����!e�/e���R�y��︃��Q��8�E�cP��.���Ɠ�ɶ�HA����Oz�,7�7������z�����ݻv�D�<��s�4����r��u��l��9zt�\�����৿}K�i�?�F=9s�<��)*�����l|xG-'0&�]fZ��T���b���<C��z(��o�� �j@�|�|��d���z(�#���ܳsN�g���9����k��N��^]��J��D�x�;rH�f����hZ}�j������Q^��P��9�Cf�0:PϤcI���㏞��7ߖ�H_���_yK~���d�ޖ};'�_>/O?v��(��RN�L�r.�h�ӥMG�&��+��h��_��z}rǇ�x,�8��l�7wfT^�1�U������	��@?�
ݿ���/���	Rڶ�| � �;m���o3����~$���T%�U˭ڱ���]9��99��Q�����9�O~�ӗ�w>RM��)'��y���Iy�')���
6���`�D��ea�*���:#�������{�^��k�H�\y�u�p;}h�L�rm������Ԏ*��*����fF����8Q2WY��0�<x���9�LW0�<i�X���v�ܾs]
%Gv.�Ç�=sU9�o^Ψ�HB���Ɇ��-�?Tb6UI6�����!O?}V޺������Nv�j�+2Yɐ��T��^v�<�����`52��;�'���dK���ޣO̼3+~T��_V�=�)SKv��3��V%qR*%W��[���᢬7�˝ݣ�����W�eݿ��]����C??��W��t��׀�:=u��2����7)q-��������Ok՗7>�*��ǿ�7?�!��nޒɹy9��0�������@z�r��(D1k8�t��ב�����ބk����Q����K�V��!�EgN�~/d�߶DX�P J�Z�����/�v����545��U���5���^��Z �
���/6LQ��݄hLhZ����"��_I�����r&�'�?!Up�:��;�՛�%�l7kbx2~�i��%�"�{���"�q�א�:+��dv�,���Ǥ�r��>9����g�ȏ~����k��N3�ē���|��������ֵe*T5���7�M=������y�ꊸ(Cca-7'�P�-�|zlЂ]u�,����s�X�ޗK�7��+���������*g��ZCC�2yS��Z��o�U�~X�> Ǐ�W߸I�C>\hH W;hK7 ��@����@��r|�����Qu�@��!��	������m���.�8�@�����rｼ�<ȭ�k���2q
�zOC�������ڙC���)kي��je�9�9��S��z����)m}�W߽(޺+I�$�|U��%5�m�G]s��|shn<,�ߏ��m���*��������!���e��|g�X��m8��W�c�Z (�5�U�S� 3�"��$�-I]c����M���^�닛�T�2�mĀ�H�%D_:�5P�{���������ȱ}rbߌ�8sT���H���oK�1�XCC��@f8��~�C�� ��l؛*y��?+_~�
q���wk5�95%j�����%�L��7���!U0g9$AY�,ޕ+�eK��J�,O=rR���q	;����{���;F�=��Yh�?��C�>��G�5��=r}#�0O����e�'��Ic�)�>R��R���z5fU}��=y��r��nٳk�|C]�;�u��X��椾����tY.祠ᚪW[H�s*�a�bf�H�×��_�0Tc�C�&�6�����鞵���k�#��:�V5�����p�Gȵ�y��oJ���_�8��})�+�lV�l%����]z2�{˰`��4�tujF�[E��Ä6�tN>�J����+��;�Js��{woNC�Y��Y�kB�k��!��;�X*����'Vz���c3��z&�����:2Ri#��}ߍ��D>��/yñ���`fA����rp�A	��'��zC���_��
-��pNK܈�&O�z2���#�&�S�`+��7��^_�W^}S�����|dB�;.�|1�[7�V6�{R�W$�u8G���#������D� Oz��Qy��^�m�V��_�.K�k��SO�W;%;�z��^���w�]qT`�y�#�p|��?� �>.߹"�+�(�U2���#ЖR���4վ�d>�f́pPV:��!�]���:���p�rHz	_=p�jVj[m�2���Pu����5yJ=��S�G��{ݑ啗�#���灑�� �R�hY�v#�QO A0�G���6�H�/�$���9�k��ρPG�7��JVNܡ!NLro�V�s���Bg��{���ʛ�Wo�D�5���Ր�J����rE�7+^�V���?�����&.Ua����8���	�v+e���"���7ޑ+�nH6����0g am���G���4��@,�c_�����:�+��o��*C�m2eFk��5��gH���4ٛ����$�ʤk'F�8��	�r)sC}&�8��Ɔ333����K%_f��믿!?��d��VB A�A�esɍTh�@���^�L�\3P�<��DҼ�%���y��i��ܷkA��2�^��9P��R|�YaF	6��$�:]��cf�;�u����^�)�w���|Q�H��$�L��g�q"�¬�2�Dܛ�y��o��|I��:%O=~S��7c�Y�d�q�9�Ӗ�K�c�hc�ݱ�M=����af�+H10�����'�z!o�9 �!��b�^+�a�����4Kr����OL�C��GPg��������װ�\�`U(�f��W����|��q��aRj��;zh����f�/��};wȾ�	���0��Ϫ���j��klnե��HifV���z�12���H����։Ԕ��yz$M�߯* �
wϡ� ����d�klP˘��.[�6�P"�����v@/��Ⱦ��&F�y�*3����6|��l�7kxl�Y�4�ps�� ���#�éG2RT�{0E�Q5�3�D�ji��Ğ�Q��	�X������jM"i�6������UI�|�iJ���X<c'ɡi.4��W�X���(풔���G�W���=��S�����w՚y1��Òn�&�pا�G7k:{77�丆1O=rN2z?חy��iu#�l\�vY~��<r��eaaA��ҋ���Y^�m��[���Ȟ�r���Oʛ�\��7oJyR�4��ȋWā�Q�rx��Ї�}!���K"��s���jsG8HY�RQ�o<rD�U���b<�Z��%q��Pj����;8/�C�����?�˯ɇ�?sl��`U�+�)���L�!�n���`�H>>�7��;���)�3_��|�߾@���Z��*A$�g*=|�l� @�_�ʴ��N�wZ��D<��|W���5-H{3��lMz���S&����řZ�$j�%���!�%��}7K���*�c}8�<�1&�Nt}<t��Fh�͸��t_Lgd"}.x��{&�͇��k�9P�,t#����ś�UXֵ+	� h��\��%��h�l�����ø6)��E!�w4�`ƕC�PϵW�FM�a��0x&�c��7T"����C���@�3�Y��f���/�nKJB0����r��NӸQ-f��IW0��G�� ��}oD�NAÑ�����$O��#�FC��C���%�P+�Pa
�d�i��bCP�o|f^�K�Id�֔ i�A�AA'��{����&'���<!��xE޾tS�3��3��{Mi�OK��˙��4�oJ���I���N`7�HU���ظ{����P���˴�3�g0���z9g�����ȉ#z�]*��*��g��1�u�	�mY���>���ge��]�����4���N�0d�j����Q��x0?'�dM��3t�g�x�H���;5
�~$���"3�vJG׸�/1'��g��7�����+�z�MU���p�L�@n��;�x�"09���u�2"�L���O
�1���3ƣ��[F>�M7S��B��}�����ދ��W=�?UʡZT$6CՀ\~M���C�'`��5L��nlia���gp���@eegZ{��8�P�����k�u؎'cyv]�GL�r(m��7��i%h�+�1�'��<��/6�u�x*p� H��!��VՂ�+��k�d��HC��E]�ښ��"�jݰYƀ!��&���:L�,��?HsĢ�����	5���(��+=� ���*�'+J�x�*?�.<f��s�e�u��r<g���
�Z��γg�ɇ��.I9?��j].��ut���;�d����Q9|`��:��*=��Z$��}ŞG������R�����~J��?E�g�p�����c�{�.C�cG�ˋO���{vI�Jb�ա��"�umP��Рݔ0����`��^��p]���t�/�)�s����z8_���l�Ⱦ�	9�sFN�/{��5T��ǎ��\zﲜ߷S��w��?,��^��Wâ�˩IN��k�W��Ұ.g�$����V'E�&� 0��u��2����LUab^�>G.fa	dJY��r�,�B���Z*�1�)Ğ��m`
d�xŔ�91��8I�|>)i�L��.u��]��ңM�EEÛ��<�P�Zc�x��)�y�30ii�����A�3,�y++������r����;~@�}�)Y��&kM���*�����sLk=�iT�@6������r���OL�������c��'D=��@��
y6��z�p�Ŷ���j�5 ��.x�� �8�Y��4��P/�!I����m�d��eM�a��e8��fd~�>ٱW_�iG�_(KVB�k�[��:f9>e����$x6�n�|wE.�^����<���KAØBΧ c�G�?��s�NJ�R��N(wַ4�D5&'UU�U��(;f�T����E
߬S�9B�M8��xٱ*fn3�w�ݹ'w�W���~�tE��_�������uM_݇N�K#G���O<.�V~�
�F�(���.�90��ƻP�\4�}ff��kF,e�c�ʨ�;��Bo�� ��&C�3��8���� ��I������O����]Y''�꜊S��p�@�8�!g2M�D�v̍M���"�9˫��X�t�=��3=�s��xb4�cR%-S߷�_H���v餾M�g�xￎ�� N�"k|G]�+���^y��G��Bt�����W��ʦ~h�4녾x�i��Z������~D�CQ:2�P�ǟ8#���*��Y^��aHW?���Ы��&|l�/%rlY��p��˚>��R#c>'�eԫ 0�Ӭ����r��y���d�]�g1q6*?����P�f�K}g�-1�Ʃ�+�q�p�{��z�Up��%Y]�����9wb7��<<,�K�U����G�㧏������5��;���K�4>9[��ϝ�gNQ��U����
i��r('����g���A�O��	�#=}��;@"D(h^��ܐK7��ĩӒ���\-��F	[]Bbl�'
�С�R�Mgw��K�� Y�q}�TyWZ����+h��"�ӻ�m��~��4���s���U.�ђ{�����nI|l�<���߿/[�*yț�Y腞t�"u绽���.F.��Ոz�%�J=����1�� �Q�h������X.6�DRNд�� �<�W1�Y���Vƌgf.�ỳ��hF#Z��)�n�
ߌ�A>oZb;�t ��.���g��Ǟ~V�>(��~L����� �MX����ڬ��2P,䥬�@1�Z~0�8�G�}�i����V�%�+��+o��ZGU��.oh7F:~�&6���2��n�����Of�2QTjQ3�dß�hxR������=�g�9}l��ەK��e�����9�gN]�@�6[�/�0)7gJ�B�
�n�3�g��?D���pm7Z�*�e�|�ɰ�ȑ=2;;!��&�	�>��W&*�n����(?������
~-DH+�ӻ���w}u��qP�>�����j3����,(��aȪ�E(�~+{Z�0f�#�5�q��d�J�2�S%�Dn�Y��FG��e��*�t��}_�W���I5�/e��r�J��KA�QF�S��\�c�l'��Ġq��tlb�c��4FN3�1e��d���/�WrdM�P��/�:"�~�tZ���Y��Z�hT���dĀ�=�g3Fi�z�*�l����ck������I�g�vY�՛��H�<�/�M�fLOM<����U"�P$�؜eo:��Z`>�|�
�+�U��чvKY��S��r��~N�k!�1pi�;���,K'hK����HVN�N�Q�<=�Hf���Ƒ�~�wo��~Q�f\̼E)u��Sg���hQxP�@�D�$\u5K����j�%ZΗ�z]*W�矓GϞPA��{-����\�uM:zH��O�*U����oJbd�|-z�%���?�X��mޝ!�E�vrU�k���T�k̀B�q�����@]{|���;r��k�X�R�2A��z{K�-���&8�̵$� �[c��̯�[L�l�Z�Q���X$�"!l�W���L��88S�ɬ*�`KzA�-����E�݅��:���ٿK�{�U�]��=	��<�0'��9z���Z*�T��IKOFJdx�Vo�p2�^Ɩ޸�Lj��U�H�k�,m�<-u��.��l.ݸ-�n�cSy��sr���Ċ*#�D�2YBo�zL҃���:�s>-lz"����|���.ŏ��o�,���F=��kÖ�YDփ�/T*��xmK��Zҟ���J�|��U7P�o�U���SO%�Wԭ�&�-9ux��A�2YN���G� $���v�9�j3yĝ��꫊�$���7tӀ���[��ю$փ�c�<�$��e�Ҿ�����N�CW&f�&jA6kM�3}��ӳ;����5�Ц���=Uf����?��\_\��Ĭ�9xHrzPV�z����E�@�܈��xL&> 9��
5C' �┓��*�[�3�:<�ú��G��lo�;�JH��d��,��z���rg�*i�:�P訞!!��\���ݻg�ҕ���1�
ђ���T�9Y�=/�RA�͞e�w���_>���,��^�$^�2 +	� U��pzr��ay��&��:ַ�%���z��4�B´��G�ՔLiFVU1��#�Ϟ�������sd}eC@�q�r<�����B��nl������~g(쩘�
f` Si�AlҲ�`���w� !��!�!�& $A���5@���o��DF����<qB�I"���ɵ�7eb"/g5�,��^ѯ�$��*QT&���h�%.�c7o��ָ�P��<�3��=��2�?���S⌼�����	���!0�3�;�C�f+��e�G�Wj ��N@d\��)#8F�5�MR��hlI&�il=Ɍ�޻"}�̿����#��1���f�����l׉4D�*�U�5�p�+e~Ζnj���|�?V%�$�][҇/����ځZ6Ԭ-�3u�F՜�@!ځ�>�,�_�#O��+�{v˗���,��5D����˷��̩�s�n]��lav����61$�U/��K���^�`9(s���HM]b��NZE�����Q��t�"�nA�5��:�iK�:;2�Vn�
�Ҥ�������A�z����=��royEn�6T_�ʎbA�إ��.�@���p�3&<e�K��p�i(�̝P*l�#aH؇�'��o�#�߽^G���lUL�r�8"~c
@��S%���CC�7���?����w���}{u]K���A{��h��HK��wޗ��&#|9c���lg�1�!I��4�h��!=�Dp�A�HlHF6Mr�LM�f�������0^�5�7ߕ?{�	�33)O>��KE�q����3/�Ν� ֵ���Ȩ=SLɴ�����ߩB�ǀ]×A�0�ʲ)�cJ0�Es�1,�}z{�����x�E����l��]�ݾp�R
b1����`�Dkܔ\�"m]�W߽,W�V��99�n�3>|x��h�
�X���ƹ��R����<�����o�;~��{(���jasU��3� �A2��!q:�U��A-�c?R��t�0�ƍE��O~!��yh>#/|��,7W����_{IΝ;*�Ҽ|��Y]�Q�o���ڍ�*���s9�|kI���/�N���7���0��8f-:BM���#����T�q�iN���+0���]ʨ�j�����[��99q`A
@�;Y	�/�;Y�ؒ�o-���q�S�ȹ����)YYk��z�y���`�(43p/��bOrh_dXi�t9��KK�D韎�}S��[�zEUh"u5
z�U��{Yf�x��,�C驗�C�S�2���?}Ue�!�=&�J2�rv�	����˷������5��0ɍ!�L;e�4���R$]�w��W�#��p{qY޿|]��|�|Y�"	�1�����Ϊ�zeU^zz'+}��>)'yL��K$��V(��Z�U�T)U)G��?
��GUR�Oܲ����'~���7��4��8FA��C��+1��p�aȟz/i�_�0�s�F2LB��&V��B��R"����T*Db�ǡ���6`C�肭mvde����k�ӏ�=.s;�Ty�莱�(C�����B��k7o�o�%w���u���\����( �@$C>��LK���]-�E�-KG-��.��R|�Ͽ*���|��S�Z���k~N��V����~M�\%/덖���;rh�N=�s򥧞��	=���8zDrj�[�!t
R�d6Ce(�;9���v�mwF	?�LA�4�@��\�������2��H�-�{@�qI���G�<!�$/�Ҕ���t�#�^�#o^�"�3 �.ɮ��'J��@�u�2��t� l��ӏ���$�ZO�g��褚�	����]�woUo5��n4�t��p�Zz��|,7��V*C�.�h�Pe��G��;��|WC���v��y�2���UU$7�[+�9���$������R�"��@�-
�#��X
�~1gx�ޒ_�#duM��H�����	V�^"��O~-Wo�I5�ʬ�ˁ]3�Ĵz�|tcI^y��|)&.ə8���(��O���>@{�s8z��L���2�u��fr��$%c7)�4�2D��l�Q,�m�I��BJo��B�@�H3Ec�9�
|4�Z�l'���?�S>^�T�I�U�"������� HJ�{��}����%����z$�n���װ����c3Lj�53Ci�qǤ���WĬ(�I�l�ˏ�[�h�|�/�T��*�-���U���,� �˳<���GW���V����ؾy9~�Q9�Qq�q}]�*e�}kE>�{Oc��*$���&�ᾤDΟ���-�X�OLLȗ����o���#(����Z�AGU,o]����2K�Y}�[����?��Z�PN�%s�E��Z��sEi�{~��������V��$f+�B�ŷ�%?Uw�q��2��
�?�qY~��u���x��������g�Jv͌IuA�z���{K޾tLJR���
�G4f�t��`{^�x"4������]o�ϘzZ84�y�Ț�2d��?/�U&�辂%Rc�W�L��t�(?^�еY�Jݘ�Tԛ��OS��*�U��EC�Ǎ�޳���e����rT1qƘ����D�,�-�l�a��2F,�X��
�gXO�y� �#����ZD�x%�P-T��)0�RY6�M�����!�H�ju an���u�<a'0�A�X`2���4bE���Z|4����HM����XϳL�$ ����^��}[s���JWÄruJ꭮��O_��͖���� C$��.��^�;*�����%<�K=l�M9�gNv��0'㩷U�ӵ�����*ΪD~�^��QQ�;�)4�n�������ˊu~��w��U����H5[�D�v�#~1�}덋���s6?E������{������{�2�s��_`_�F�3Ӳ�׾~�\�zC:�>2\����i�g�@%2n��L&QL�i�%���fGb�U �}4]�A9��,a�0&a�'�_[��*�|�4bB�� �c(<p�f1��#��ڜ^�����!5����1��JŰB��<'�qA�}0!J� ���r��z�P�o&�ѥo0��(���fS�^ݿ g��<�r��E�\TI���G�)�}F�,�pVd,��j��4R�~Z�Iluf|j��~<B�Jڰ7vI�,x�ɍ����t��q��2�'��xN�1��P�A�������5�B��#�/@s����)y� |�Ԇ �`W|(BA� �Cx�Ia@����������f���Ȟ}��O�: 1AP�	��l���o�a#tb�@Li%ba��_@/	FE�1�w?�X�-��#���7�d�\�ջ���^��4���3��!*f���ʈ�%%t���9k� �L�F������kH����UСh0U���TܤJqs���<��ދeu��S&G�+D�K:���C	�~ )�ޚ*&P2D��� -�r��y�x�&�I�`�nb,eY���6|���L�k��t���f��`��5�GWn��<Bc�s� M�
˘O`F� E��c3f4)n�gZ(���!�8CCYF�@Qpf����pTN o1'
�}2r��U7�lh��`�g���x�	t!�u
*����	0�q���XS9�%�=�1�q���^c	�7�`Y��cO�7G�R+$c	�ȂÜ�g�+��A٢�����c*[F��C��my�d�>vY�d�K� ��S7o���B���%xPS,�%��e��@�e,�Y�M٦43��T�����M��Gc&(�ʂ�9=zaT #����hMt��E��^�ê����T@r*�@$��\	^�V�m!�j�KCdTf��U��������ix:ICC���:b�"'��=΋5eF��l��bV6���n� O�� 15dI���6.`��&���v�����&�p��70lT\��7�PJ4�J�z5e�����0�q�ci�{��P%u�9��Ra�K��F�8,�����Y�x4۷o��߻GJjl�޹%W�~��jhXڑ!�(�d]�H�H�J���r=��LO��0ֽʫ�aR;찗����B�o�C<Q�$Q�V��u��C]o4� ��E��-3j�b}ޜHF=�B�(�f�ʼ\.3G���f#z,�k�|� �@�7�]�C<~��cqi�����4"����D���aN���}��c�Q:��"���c�����&�!=U��AAt�k���U���(����lB9edy�C���\�?o[`��X�T���A�j�1~���> �:�M���A���[O�ט<r*f0�R�1�g��xj�˱���ģ��v��.�0!	�5�x�XH�{��Y�ػc�}}�g���`A�U�zQưe{�qM�#�V��P ��dNEC5�%���c�6v�8�E��
��l8������\]��ܻ6%�d�M�qP�͗��a+����6���l� �<d�"U"�DE���p\3^&���A��JE3#w`f���@j�=>g$��*�8ڔ�Ze3FĔ��v��FJ��}&T'*��ɑ,8�CV��͍M�<m�����a�.<x �x�2�<At����&����L�ã��gt'��������!�T'd]?���j�x�L6��=�ic��jr����?S;FJ���)��B����z��=���&�����`�L���0��[u3���L.�P�T�(951��z����[DU��/2��h�=��Д��@�
�x�g\Ɍ+�n��r6�y�����z��GTg\���ZG굺�Iȭ�����h���G�z�����Mc�OcߦF�����]�3[�_|I^z��OOH�X�R�(�n[?B7����Zܥ={-�����~����Ut�@�]$1n��N��Fj�����@��Zj�=Β�0a�X�!���+	a��캦��C�Uf\�Ķa'���1�A�b �0t�3�!�&�Pr��]r��싁���g�	v�SLbÒO�`Ef^)�%M��q�\���K\�,l��b���z�F�;fe��E-��i�\C���@b��|L/�者+0�C��z4K���\���T�;�B��
��� 9��g�ӫ�R .�i7�XP<PP !B�@a$v�B���cWL';�| ��L��:7m�ȍU��D�U�m̧�!��[�� s��A��Rbm�sw�ĳ�?z@.�+��.�N>R�g������������ǿX�D�a	��Ne>:���D���&�&�q1�t�y$�z2�]ev�Wr������H�$�����)��8	����;ߔ������~��D�#[(��Â���ˎ]�,pm�E�k�������@ȓ��Q0B�z)����H��1|Km(&~Dz<P�B�"����pZ�wg:�e�`��Xgb`��9��A��V��rx�!��;�"���� ��~ٍ��s7���"�A!��ω�c�>SEKƾg[Q�xkS��^�$S�pFN�obB�і��p�s���0h,�����5`�8��~���L(�yB���tr�sx#?����@��u<��x�`rG���8���d�����ƽe&Z}UB>�F?�{�h�}vUKX�t��K!?�P�4�<�� %�ci�!+Y��Q���N�F���LONJ�R�	�ݫ/�/U8C��G���Δ�.�P�%�>����[�G���~�7Ħ�ϻ�����mj�n�k� ��G���F�O�^��Ք����'�I�M4�\IKa������dj�$��*���`��!Ac�O���&�,��:}Xi�f`��yd�ʲa���a������0	mCTV�F�3�V�+҈�z"ț����D�_�1�ǡ-��t�:�t�-iʹJNQ(�0&��kÞa�������!���L���!�i=��c�����a�H6�xxSm�����.vS���r\Nb7��	����g�Xv��t��6�g H�b���a8!+>ǆ�
��g)�#�J�K�t�w"3��ņ��$Dy��pQl��6������}ۇⰚ�DQ̍�@���l���0�=K�ޖl�d|3c ��2Y�Hf�&e��i��=�Dx=���I��Ұ��:��&i�P9�߁��2o�VC�I��}{d�¼�@c���$@o�k!;)$>���^���Ǚ��i/�3�}�r��)��a����U�����DAYZo����a6x�؏�NA5۾/�w���i�t\Y�J�:���ͫ+�S78@u��n�d�P8�P;@�1s�p��گ�	pOyA���㙰��S����z&��xD��"�ѝ�Bϸ�ټG%c�}�`܃ZӾYd�*jleW��9�8I{��-r~z�X� $/6�[�_4������ӍlY�M~�Mv��BTNf,\i���ã��嗀�-bA#���jdJ{i���!��]��T�8������A��9��~�Xv8����|��~�>K�z�4̚P#[)��%�:��ā4#@�!x�����-e�^�첍��t��A��Ԋ�����J�Qg	��=�І�b	6���V`�װ����,-������azbeB�g�G;���̔�>Hī�@�
���ٍ�7eskKr�"�@�JUv�βm�V����
���Q�G�@1���7���O��������(�ł����\b@�74ɰ^���4���S_���P��a5\AÑ(�߀��qRݩ��5�y��l(�p0�0��=��(|�Y2�}�/�v�\MK[�)�^�䮿����r�lu���[� �P�:�� "�&g�����t����� .���e�]���:����� �H�e����2��4����Ɲ�A��u��g옟�;��C������>�'.�0n�>��<0
�?XC�X^e6�%��aB����_ q6%�*E��5Y�AL�F����yk��f`H�r �I
�	��um���9�0be�'�c/��e]U�(����D<��G$U�
V(������R.fYQ��,5C<�A_ת��,���ܾ}�bRm�;MU�m��Í{6��T��> )�16`�9"��?�M8�g�:��n�Ѣ�Y���n�;���,�5�F�~��@���NO�eZ���TU�P�Y�5j0A{��*�xe ����V@�Ǳ��1?>��@e�����!Z�?�SԢu�۪X�[R.dd�R�Z��P�~ r�����<��Ɉ�����ms(䮨���3iܞ���԰�,&���a:Sn[��(:Ĉ$��%S��Q�dH�2��Ps�*ϸ�(o�5���T���2�J��J���&�^�%]�X��d3y��l�Ğ��(�&=c
�=xؐ\��C�����`� �b�e ���)t��	 �T�,h�g�N� �j{���<����dr	�(�����`�}(oI�Ә�91Q��j���g¬,g�`ɠH
�<�>C]S4�m�o���7�Ĳ�1��%Ϭ���+�fHz}�������Q���6�x�^��_��π��Li�c���c$UA_ѽ�:{R�ثC[VW֌��䢮���{���r�Ï�ߗ��9v�t�M��\�� �@=�"oP8�$fy{��1+�!/�ςf�;dW��=r�"�){H�wZ[�����A A+���`�r�ekU����r�������	�Y8�&�0<����V#�!V R���+�&PՉ�T&&6���s��K���J�I�P(����_}ۥl����e����A��gi>Kك���A"ٔ�=K+0B�2�M�aY�\�6��hx6��]ߌ:J�1�
S�4D6I��`)YlbcT� H�gېGd(#Od�����TВ��d��b5vzUߗ�G��YND�8P���8��.2�17��n�$����\� �J]�{ȁW��u,D{@�*�>�Pw(b�=@eY�<'<�����9��l�/`�C NTv�҃C�v�"����Ml��!�X3�V (��ΩA):�����:"ƬH���*��=�k�@�ӂ"eR46�P�\@�B�TR!F3 <�e�:�l��!� ��������``&"����wZd��p=;�e�Ձ�Z�����jmR�����b��q0�T����[��9~�a9�I�|��~wMz;	}�B�&�\{�x8|1�{��r�E���4��Jm��!������m����n��Po�%ރp	oP4��<���*"�{4,9&�������/���g���}�h@3Òﴧ��(�\E�e�bz���vu��������8�I
*��N�?��p�;�0�v�����ji��,M����g��HL��sx�f;�$]08%���x$��*��R�	[�f���P���0�f4��K�x9����!TA�e
x]s�ƽ[fS��&f�9<d�!$*=d��S�<��~x$l	��3`z=�,rQ8�i#��F*�t2&��r����F՞^lf� I��w]��%�2w������S��-�|�X�W����#s=���{`(��ڷ�90�
�z��w���}]�@�9TB�5���D�I�R�Pk��*`P:9�-2�a��i�f�^Kޯ�kkY��4�x����r��A�I�y F[G���n��`]\kh6o�{ު񰓜{`:�#�������M)UR������mh��U
%�
�f�"F� ��*� �ݡ|���}�w�Ƨ:Sb��Nܕn�K YGe�Bl(?$M#���VE�&R�}z�}Ti �K���Z��ܣGR���>+O.�0��p���[7ysCÞ�e��ףֲ���-��Դx���[�ыAr4H�rm��[�W���$��V
]kd��;��c9J�<`4�.�m �9�\%�Zt� 4.Ab�q_��S4�cΚ=�>㘦�N��0$��lH<+C�Ʉ4)S�g�	-�a{b���-t�b�:�A�1Ywx�JE���Y���������C6ok�T�T73 It�\2]1 �=�d�a�T�TVg���1n>�eja��N���ܔ��%�zs�j���!�� ��g˻� ���(�A'�B� �zj}b�ݤR*�լK�e֗:�VTE���5]�ELR�c����p�p�6��� ��^��T�k��� AU��*��CG7�@ �џ��V����Ak����
���Wv*�	�p0��wi4��*�"��Eբq�%6�����_��|p�#�«��AY������cFhz	� � Obs8b�Ո拘O�jS�צ��Aih:�\���}��ꍓ��i0"�D;�S� e�d���'�YGĶ��+����ay��B"����TPo���z]�-�Ik�^�UM���Q%ת�o��l=�ݓ.@g0�ClUJ�d��cs���6�,��[�И��F�*`l�a.t��b�#g���<%��ب�" y^_���*��?-Y��ӆ e,?�X���|r{z����Bƀfb�I<f, �r��\��� h��u��+p�et�n#����a�Q�!F(P_�]�]���J�X��6섈��9�O�~��5V�P�]���0�
=a�GnQ}9�h�T(S@d�;��U���0y`g����o��a���`�ßA+��YW/n�G���Xt��ceѼ�J�-��"��}"��5�	<zz@o� h���q8���^���#�B.����l�z��p9 %=�����c�Ø![���@��^,=d}U�p���,�I�;ƛC7l�=(�ܺ�(7���!�ʣ��%u��!ǌ{�"�����6�h��� жVwT; f�A��dO�N��DE���8��
jX�!�g<�,����yA���SB�a,E��Hm�g�l��-�	C����J-W)�:���Iń�0��ui���R��������1�g�C���nf�����Jj���JG�����Q���C��E�5 �guS&���b9�Ɔ�:���mF�g�+��g:��a��X���*Nv�Z�0��dW�(F3a����]ǰh*=� ���Ҿ)����M�e��\��H�">gj�H��AG!��	��e�@�q�@��O���>�� ��'.ɟ�v��U���>˟��j�aN[�d4�nrL��C�ܥPQ��\��$�����d�4E�P��1�1S�U1�C^B��J7�Uo��@�UkJG�\�`G��%<87��Ν
�1/@����w]�>�v�ة^Q �z]�`(-�(��!c��A�!�`�A��AW����)�s�c<�J!'��i�W�T��X�����e��hE�#0>��j�Y!AX�v{�EД�n���C׉�8�d�l�檜#=�$�0g�G�|��J�{ʳ�����;R�����EV�"Q�ئ�Ӣ⇒Abr�^4��T~P����W��k�V$��u��T���Рt��S�0YɑN��;(�v��T}�W�kmK�&��f�â��J�[��;�X ���m)�v.�G1���~2c��B���i�;��|H�/���wS5!F��}3٣���]l��i^��,�yt?<v�ƑU��:a�{Ҙ6\�?�c%-D=vH��x�ׅ�m2����r~$AsC��*$3��qqHQ�ń3��{f2���d�윛��{�e���/�$W�!	�F�![�-YƜ�[���VS����
��}�����z��c Ċ�0	W,M�.�;	�� )�V=��吗U��&]�#�5`���8]�����v�����VO!G�fY�V$���9_:j�66�^��ܺ�*�n.J��aF��ߘ���cy1q�aP���S`Lj���J�0��R�5�ꍖ��Y�w���T/����o(Ǵ(����e�Xe���|��	��0H��f��Z)oQ�ܐ-�.��q���.�:��z�0��$<��C����~[�I��_���9~#��d\��F=���9��_�B�〹2�)Պ�{�Q�&L�����e��[���� e]S�Vo�Ҏc:`1ջ��"���#�8���/��z�
?&Nf Bxs!f%UV0h=0�k� VY�0Σ�jx���7̠s2�e���'o:{	V$�ZöB��ŭV������Fgd�<�D�{^���uQ���GH��k�bT|�j�^�V Y�A�O5+B�{x��.U�鐀��0%��a3��VbƫFaؤϰJ�?;����A�1��
\m`(С
�1�H�H9��.� ����z��.*I'��r �u�ڲcǌ��wT�{Hv�WA�JE�׀�LH�:�d�i�;�{��u�t����K�xo]�T��L��
�xz���Y�]���sU
&��H�bM�w�LN�Պ��{��	���
#�c:��D21Y�Nʉ��p��g�W�o�]@��to&�2��kigȒ���=���5��kr��41��a�U�eJf-h��2^Θ�cD�	B9Ul+�e�h����	��G�i���Pg�C�c�x���)���,�0�3���+����$��E����<�^��r�*�v��݋���&�U�5�*!(mP�@�"�i�z�=�Dd�P%��v�ϐ9���'���Y� ,��}3~���л�+@2�<5;K���kn�<i"��67�9� �j�qɠ��:Ex?X��_(��R4 �@��'LF�� �T�����R�����H�BƥqC�#�g&�W����7�Z3+|��a,��z
�*��Ec#�Y��F�E(L��R1#3�S�V�C�¿���,C��q-0e���l�(IEl r���g&��l*3���82�2��2��$��/t�"����p�
2��~�Ϲb^5���` o]i��M��n@�.�`�\N@Ʊ�gNʩ�����2==m�V��p��pFy��Opuh�P���^=��U˴%������ևd/ϫ�����#2��b�X1~�Z&�<H��.���7����m.C�N���<z_Z|�ə3gUy�J�Ze��Sd�(@i��B���8Gx�DJ(�jx�������Α��ڵk�M�V���;�t���DA-b��L�b!Kź�9�
�T��h�a��^K@8<���N���D�9OJ���8��.::Y��0�w)0��3.�ar/4��JR�2&�-p�����#�V���~O=3�Т������`��? 9��ͬ$�c�H�{�?t[v�� �F)=5�!<;�W�=����o= ct{g��+II͍�/J̈́mO��b��Zbx�bIZ��ʥX̻A�yye]=��ڽ�ecG�x};�>��{}�f�ϔ�98�����i!�����]�hf��6�m@x����O��X`���أ��|A�JB8h���K��6���0N�;��;>�*�O�o���o[Bb�|�(r��B�y�R��䔬�����!�\3�	���-����U͏�rk���ӏ˳O?'��s�]ܖ��� 	@����N���qVi�,s�ٚ��.��������~U���k�4���
�NOE�����PR���C���t��k�4d��+���:p�o0	|��9w��ٳ�k�u�~��F9<��IN�_VkQ)M���W����� =���Cp���dX漷��^�G*E'�R�P^Du�t�l7zOCp2l��U�"�D�%ޥ�
��a�|�4���^k��VMײOt0еN$�3j�g4,s�̐���|�aHΌD����]]�e����E�����q�p�٣b�$b�Ѐ��2(�]=�H^3%��<�)��\�p��t�s����v%5V�ӓ�k�$��'h+����S����9T�<��TC�0��|Ĥ5*e�'V�.�3�& ]�*ۛ���:�y�ei9�L�T�x�L+�y�Q�`!%�3��	��L�)���>��k�� )��$b�΄	eB�Fdi|}��*�Y�Q*@�Sɱ)^>/;w�`�Z��W��yH�Y6!z?�8!l�JKM����R�,��f,3�
�* ���F���n'`�~LM�{Zj��~'�%9u��|�� ��JW�&�4ph�ݟ�Ш���l���'���k�)#?&���JÛM��3tg�2�>���؄�gY��5�ƙV2��s9S�g�LY"E����g���gɻ��6V���<�K�a�~�y�s�1뙮T���Ul���}5�-�����`N���{���o�bk�{�v�h8�xt�>{9��P�(��}� �SƏ�� ރW�>����Re��ϞTohA�k	�L5�EBuϞ�R��aIU5�����8�� 2���+���bڵo7Ï�[Tή� �׌D��2�p@4T�й"�,�-���u�6|�g�ˡ�dޱcN=�I���oz~��eό��BO��V'����X��b�̼�iX`dd�������
I��)�}I�OڶT��t���!	3ރc�wy�����B`����9�	CC��0��k� ^1�Κ"��̲�B�%��/÷]� �(�o�q����	C���#?�ǉ`)�=A)6���ӊ��W2����b�7B�,�215Cm並�j�E_e��0T]<����عG����:wo5�� 3ƫ��'N��<����W���!o�)���]
<��Ԭ
ش<���z?��z�vxTy@�����$��%���=BD���T�j؄�)�*�zV��9_z�������`�d�����c�3�p�ɘ�� �j@�ct'�<B�FGmG�f����rwq�����y�F6�8B���bK��V�Ͷv�oP�����pcbFJ�"q%d�So%�-r����ٿo�옭ʎ�*	��(�#�=�e5[�4�m����JC�9�D���WJ,���l2>�$,ɾT]4dk�!�j�<׾kCuC���8l��Ȥz��RE�5&~QC-�m�nDi�\�"�jSS�23;˽�:�z��!��~!���$h;Qrmu9�����L��(!�����T'�`/�������b����B�>�8�\	����Q�XG����L�!�� ���U�����h�q:�k��Yk���/ȱj�\<=`���\|�"�%�anBh�(�82,�bY�Խ_y�I
�e�!ƭ��\[_���gzbs/���������Lt��R�:�3'�ɣ����j�+���4\!�9d=C���Y|}�p�=�[�C�஁��a
�\�h6k[z�u�97%�>(�z_�~B�7���
Zd�AdMp��6���ˤj�/�cصsZ�?�$�����vT�BS�b+~2��s��,�3�W�C�i�qb�n ��K��c���z����ڏ���׽�o5�wN�Zӄ3�	��3��0ɛ�c��/f҆��@��F5����`8��C��_o*2�8����c��gK��Y�-��~��=)U'��k��=h�``��*aClKɉVT^�.`o� ���)�e��mw3H�R����1�%<B��D��e�˱Ď��YU �9z����+���8��Ks�R�!(�	�xO[�(� �� ,9H<N	�M��G�J�ϐ�|%�(A��D*�F�:mCI��A�y:�B,�tFf#Ld�о��H�6��a'�6�`W�}Ӊ-fĈYA�b%����"�BO��l����frشm�	,IK����d�#���d�@�W�Ʊ��!F��;@�����,�䙜B��rp�ѣ�iyFwf\����]B��u~����dlω��0VE�&=��Hfa���qZ���+{�/9�,���=dj$4��������K�=�|�������r��ᴪ.�UЉT�Z�;��f4f
��h ���pw�kW|��]ai��w_�i�0s�;�����>�H!K�Z:������vǲ��p���ux�ழ-2݇j%��Ɉi���K\	ؙ�uWn�IYCx�9A�h������IC>Љ�д��F#l`J���S�"C�t[�c�nuɼ*��ͽA�ƪƖuq�Ko���VPp {m{���4*ڡtu�0��ˢ�)�-v��5z,Cgg'�'������g;��4��IE���DH�P�I��$�KߨY"�5��>���-�6�h8��z���b: 8�'S:i�!�)mX%�@�-n�X�>еQmu-+���6WG��{$�㙒%@� � '�̙�Rc��h�}�V�*^�PP� �����b���r8��I�r��[��(��Gj��೨+R�)���c�&�$ڛ��Y���dp�]�[������%f&o��UڀA�1��&DI���,n<K�..t������e ��c^�p���B�g\�.t"��&ރi�K����eC�loIj���� �ژ� ]s�=�}�axuv���+a/V�B���2�7��	��l!1��.�����/�,���
�{�0�[���i6��J�'�2����6g�N��YD(ueV6��(����\_|�y������wW�~�����6�2x�2L
�KC -6�B�M�ySƠCڑ�l[�8S���5L��y��~��G�����-���`D1
m�- ה6��%�H�%c\8
�Y㭩�l4��+��#!qv����7K��Ȍ���$���S`�_��v�Bנ�5��n��eU��nv@f�셬���G���x���F'�+��S:�:�z���	q/����&�-ux�����Bh�R�Q0���6uZ�s�
?pCTѫ�ݦ��ѧ%Mg�&c�꠱H?v���}�H��Ué�6)����-Gʥ�#{ӷS��iJ����M��G��],61|�ȸ�<�N8��@\�>�sJ����*|��O��9Fco�H�*V�RV6�C�j��IZ,26EKY��ݰ�wv�&?{��n�X5*�Р�S����KKc'K�֢!�te�B"�ĥ*r��[�̳ w��>��'Z\g�ad�ӎ��Ą�6�'T��Q���ih�b��+1����	ؽ�L�����m�\�@r�������O�� ����q��ŚOރ͂�N�L��Y�Q`%�޽s;�>�%���-=��$�Yy���W������}�n�0�Q{>sB��lLJ�9�c���c�el���28����PO+x��ɥ�M#�k,$��==6`�p� �	A��##(�������T�l�8�se�Hhٹf�:�'��}��yx��0%{{;ꁱ g��0Qu/�Ϻ\M
-o:M$+��3- 쉩��>��Z�R�_k��E���׊�9e��E���J�[s���U�3呣�U�{z7%��v���0%��	�I�OA���Fs&����Np����*h<5���0�$O�	X��{�_|����DwG=[���W����[x[�4��To�}C�vn���%#Xb2�d�'4���ޠ�q�7�kի�n��Z|��H��}^r,:|6X*�ob%�'}���V��x	IH� m�����lM��wAڂGvf�}i�6�O65�V�"�x�=��Xf�M�g�j�gރ	q����{,3����S$�����Ax��Q899� r,����N��جW��qlۦ��L�����QC��I*�L- -�H�M �R��v��M��0��Yܬ�ZY1^:&�k]��I�:!e�:u;�2���uqXp�v�`S����Q� H�-5}�<�;���u=05 �������)&u��Ђ��ݝ-���ْ�by���(qh,�Y!�ba���[ǖ �F�͍ƪ�H�J��8�񽨾f�&{��ʿ��*3��{��5�gm��^A����OE��4<pԫes򲙑�u���Z����glf/o�DD��TX��	=�Y�  �Y��qu~���vc��f� F�x&��//n��fTc�R�x�D�b�>��W߄�p��nI�ʞe
O�,���Y�:�JW�Y�O��̽��8r����RP�l��e�s��ʱ�`j�k_ �5v�im��
�?0Rm��wb	�e���MԆd	���K14m#����K��'��e�N|L�hx&��$� 똬z]�EP�}r�������VB�������V�l�q�����A���A���$<}�D��}?v{�;�Y����Č@	�W�s��F�������\�����>�Z�*w��a-��:ۚ���W���XMF�m'c�h0������3 K!��\���������{;�*q�'u�ݸ�=0�mO��̵g�d���>q���M�8i�����<jW~ЗS���u��@+����".� �Ц�CRF9�Y-�?��PR�\�򽃈Ƽ��ީɩ�h��͟�	����ko �6�'���Sˇu���[@�:�z����N����5��vv
��wnEP9�F�f�?m'L-TMC7s"�[v;[]o�j��]l.����@�-p�<���6�Tڞ(^�a2�ڋ�	x�re/]k�{� �w��7}W���ť)<��ۦ����bF(����~]�	4�~A7���G�D�&xy���e� .���l�-Nt�'j�	yp�����C�ز[ܴ�6�0I �N7��>��#࿶�0�>;����~'�Ύe]/��ľ�as�Q�6j��R�������O_)Pnww4N&�����\�ϵxS0p	PUTP/
���8`*A���ZUq�؝�]�֞�=��N�I�u�[_r�>(��� WS�Z � ��Ͱ;���Q�a��+�h	��2����X���+�	�[�����-ː���j7�-st��,���뒵D,�e����,6��Q�O����@��P"��F��N�ͪ!���Z���5�E�������=�H�g.˕�)��e����Ix��Jiҿ��KXM}yﯲ��/�8�$8KG��k��ų��wu�}�NJ����U�o��S�6�v�#�苪�r&��pp ��g�)��4Hl/��?� 窰m_7�2�Q��1��.�K*Uݶ�b�i��F��0:*��ւG���c�Ӯ=�IM`���zz�ZY������77�B�8���Ѽ\����}S�6�cMjY�DH�Nvw3�v	�x�K�x�{[v��Z�QIU�.N����սX\ΥHN�׻wOls��+� /�^�,c�{iς�XV���(cP�ꛯd��$�ރۚ, ��)װ���ڷ ��-5�gj��Ч�kح0F�(�������o�P��V��"�ý~*5U)_n�:�	�����|d�x����28J�����;S	��C;jv�k��<��ICJ�=P� �?���Yf%PO�����2�v�ܞ�T�O��P�Q�0�Z�Rw��)7:s�Dr�"�.f�Y�6W$�zc9
�C��L�넇�ɕ��,�C�6��+���y�o�D��J���D�/��_��^�5��ΫUo%5m��7�<|���N��[�D����s�g'@v`��}A�Y�,z�r��4
\ޕ��V�쫆-C%
�&�g���5�����Q�A26Ѝe7�9�8���V��:�h��1v'?-�̃.�-z�Mv���}�7⤶��ɒZvd�ǥ��.U�P�MY���j+��C�t�I-��^&ͪ������r��,PD�1 x5��NN�-[�ɢ�`MZz9R�y4�5���U�0}��|"�������ܳr����eVv�)s�A�pe�Y����D��Yp���wL�T.mS#;	����M+*��K
k�F�ci��b�.�h�j������P�\�/�B	L��3w���>�-���Ev�r�M�U�BJa��{|�HY����\�N���O�ɝc��T=<�3P���$�Z�YD �j�&��}f�ج_[C�oyG�k|�ξ�nr,U��}��W-����T¢Վ�jof1���7��� ��o�\H��5�)�D���Î����b�IJU	���R�y��]�ӈ�N�~1�l�GĶ�*Z�Ʃm���k�CW��NDШ�v����91��qa5������$L�>ׇ�r��$��tm)a߃2|yK�~D};]B�%��J���T٪L�4"F1�U���c��;�
��B
'�GX���Nǭx�B�6~���	P�)�8��qy�����Rg���%=�
�)�~v��B��n$�_CJdlܼ�9NP�0p�ZZR�o*�a'���ҙb�[���P����c+a���/�D��{e�/Ϗ�AþN���Щ�g#Q��ILx۝޶-�"Н�~%%S���manf,��2�E��$]�Q�Rc��}ur�E?�A��bն%�i��'�(fh��ܛ�Q(:����}��[0��i���?�u��ꑠ��c���^��9ݡ��l׼��'?�}�܊�hMϮ襰���>������eM	󱲻�L	��<���i���� K}G��� -C~��R8�I;���* IPnn��G� �XBB#=#�0E�w�hY�u`M�gѧ\���ۙH��o����kB쉤���;l��V�J���m��v,�\Ȁig�@���Ԁ�M5�u��(/�B����շX"i�X��M����5�U��>i�<U9�OP�����+��"�U�t9��:�~jg>�w'w��o1j��6
u�ּ
����>�k��<�`��F ����Df+y<-��6`�'4�4-ܨɪ�p�t�J�:fX�e-[��T3KaE�R`�\4Ύ��BLTd;z��p��y���ݝ���e\+lTR�v�/	�s����Q�_
�Z.�@V�)+�,�T�BP�+���4����K�L]&X1Β�f!�U�n���Hr_��e��j��A ��g��u@�o��`ϭd�O��$϶��5����=��=���u�pGv�l���C󷰲�۔"�zu������H�no��pYe*�1v��k�I[*;S9�Y�dET��d@14�M\��˿����=_�0d� S~��O:M�"���<�g9������gN)I������}�c-D��3.��d.��/�A|P;�T�4�8�*i �$��[ � �1~�kp.CsS�L.�y�NC'��ר������$��\*O�.�jx1�b"��}x˯͋omӤi�� ���uDbfA�׿���R���e �Wa�v��;���c�MRy)��L\��L��4%F���[ըØ��S��V�c��Ac*�v�TD��j}�%���j�IE��ҧ6�����B�t"�ׂ���i���U/�+Q���eA��]�N�;����A砶ֱSn�rYLq��|U�ѷB.�� ���~�࿐��5~,(�."�K�E��M�U���ct�6�����W��s���L�Y�6�y��"zU�u�����;N��L>&�ۣ�rG�����'�V��߷��T'�,��ɩ{��(nཌ�D���Xe���+��]Q���҇~ٵ�o����W�Sš	?r3�}��K�k�"T&������Cp##�j����K9\�)o��p�Yo�$�eMV���j�`ߴ�x��͠��K铐zDDk�t��S{�Lgba{��[:�\
��=�������:��F���dTp�&��E�ot�ۑȴ�ε��u�ձ�S����N�Y�������a:^�����L3����g�o��\i^f�D�oAƢT�Ѳ�kk�,������~���ޕ�)R��H,�pvq)�>B: �d�X�:��V!SO�G`W1�@���2�ϖ���a����S2��T/��x�fp6�tI��� �Y��q}R��T�<�8n�UZz�t|����  L�SWT�.�m~VU�R9Q�wPZ��4 �>1g�g�׌��J ���`ՑD � pd�ۖ�r�l[AQ��m��x;L֬l�J����1��1ڶ�����m�d#l��׭�0��_B'<+�-��ً�Md��J'������e�/:����0$B=�*WWФ��AY��N%Vz�El�����P	�YD��W5�{��x=Yy�~mh��{جJ��8��ڜ�����M~S�����.�\V�0nC���>�f�2�
$������u�G�=,��*iH�Me�8׃on0E`� k,�B?����O������o"��i�]��h�^\��Dk�h7ノ�����y@�ʡ��n��]U6���GDj��ķ��u`.�2��-����R���t���읎����c�( �\�Hz>E�z2�mS/��h%@�=dYl�Y�����3�k����a{��j�N8��e��2�Ԯ��ݫ�^Jq9hց�8>:Tf.$DQ!�&��/�L�,xc��lH0T���kJ����+��\C^i�6��}��S|"U>�i�����m�=MRZ�-�0Z��Rߊb=.�욣���d��7�ч���4���3����8����Q�g�Ά���Je��D����0�cIE�ƌ����o�[��c��eD�K�RyCe>�uϑ*$NWK��Qz���#�)���!��X�h��F��tq`J�R�O��EQ��
��ǊE���؄�����~���c�w����M��#(Ò������\ɚ;�� �x�=�2g @��������?�����/��õᶆ�%=6 S��΢+���M�ФF�L�v�Gw�Q�����%Lrd�H�~��,\��TVK��b�[��=�|�LP��Q߾�{��V
Z(�էr��t�c�m�������m"J!�82o��OǧkS#�}~}~��?hju���z!����a�4N�;'����-(�(�S���
@tz-/O��?� P��O��X^�&��� 9F���+�y��kywE���T��5eE��
Z��@	�ܯ-4�v;@� ��s]Sp>�x�� E��j�I�:�#�~m��Rk ��[��/��#D,P�m�DBP(������3������{B��gBb�Iw��:�$�麴y��h�A|a��v��)F�S��VqZ�M��)4�l���H�1o5E7~UQLv������`Zb���'R���i�1�<?���	)&m��}=
UH�R+sn@S㽃p��}�Ln>
��0XKe%3�ȿ|�$g����<��ITj�
d�v��r`���\9Df3�#�A����7K� c��۲@y0
=��
�z�K��X܅M�h��(�k�T�P����@B��v�m)��&'�y��L$0�	*O�w-X,���~
�׃�p-t��#�=N����E����C�\n�Ixm�jؿ׽{�?<����!�
��"�ax�Q�	0d%�;����'�S��y_�9a�9Y,�bTFYc'=D�j�Խw *}l'S��7�j�R�Te&u���H��]�ݺ!���Jr���+�I4H�bg��2u0.��T֐F
�%IB�Hh�ck� L��?}�4�����ͰT��19Y,����Ğ	n݇Bdy���Y��Jธ�u�u���n�)Z��\�?�ܢ�R*������L�g���	}����XqM7�B��ґ{e䰈���{) ���'.i����l�d��H6�Ye M5N��j}z��|�J�s�f\�Y��b��F�^d �2ҹࠤf�O�$���Z"�Aᯣb=�ɃX������d������ ̔���͆������\�|��0�
;l%��I8��6��iĜ]
	��.�B����iw���p�j*�����``���V�2F��(`Cg��T�I^���ޱd`�g7�a"a���=���)v�����q�Y&ջ����Y��mB��^%A�S�l�L�^P�I��B���D&��?D�����2&�@��GؗF �h�U��MΊ�ȩ>o�ܝb�U�:Xv�rei4��� E`��̉��Nn�sG��l4����,��>ݶ���E�Į �_!��6C��,|������r s���l�'�v#�ڙoe�d�u�T�"/�G�Y�~�y�1!IM�8���d�夿n�+Ux����=��m��9��W�5��qe��Tjh�q�B�T�Zui����d�v~x#��������
����g�c �'d�axqz�{z.%��p����4�}lEG��O�&{Lw�KZ"\�jƩ'�O��G���eP�V���tg��k�iJ�f�N�z�.�mΤ^NZ�Ԥf2��@��8kxZ��4��,Z{�=��Z;���&�Q�`�-���R��	\��z}�vP"�\�� D�'Ws5Pq��P�c�����b�C������K����Kꆔ�J�.��2���[`�1��5��jV*�==�{#��;�x�{Myҷ�Jv��^
#�LEsrn%$�I���n|�>��=��=�GS��2�(�L!DlVQ���\��� ���gi��-쁤7�Á��拡�1�O�i;�)��)2!�է���O�s��}�#^�"�0�L��o�
^�K��^�/��^�X��Q��BR��
s���􃽩�R�(����d��;�N�j~����Z鲊�{�4�	pK��8G@�n�a�������7�3���SP��n0� ���8G|eޝ���ֻ2ŉ:�g�,&�����Z�ק��#� a��,ܶȹ�`�H��W7�O_}�nݕ.'D��Ɩn�D�i���F^��A e�����z���X��tY߀(��r��k&/]F	����e��٩�َ���$�q	~d!h�,U>T>��\!�vs����m1��!]f
æǍnaY�����q��3��D �D.N�-�v���TX�E��E�ވ\��CY��W���P�`i���Y׺�����i��d(�3�jX���%Y��Ǐõe�,@Y���+eU1U��xt��+7�T�m��ȆP�j�m��.-�L�v3l��5��](0d�>��y�2H����B�Y]'^/5��+v��=d�m�EV�B�C^�1��J�+��؅d�M8<��^Z(��٥�WG}�j*鈴��/��><yq���=�8�i&�b��=�@蓔am�
3m �.#�=$E�\f��22�3*H;��T�y �%�i@PN\�{גm*C���UQ�_g��'���g���T�c��������F�fõ��B��s\0l���BIR�Vm�t��>#�F\T9�&���������٫����E;�D�x���]0�cJc7G��4���)�����?<y��\)�y]�5�Y�f�6v���a�ݟ���������N�t�SFr���@g�ס ����s[H�̋5h垨|�ќ<踄/^ZFq-,	�	H�*�OF���B�=�0���_m�����_?	�L�\�9���4���=�r��P�}���9�N��}{>��P�ɓ{,����F
����0N��ms�Z�/q��p��m;��*Hy�����ɉd H�و����}��2Ϟ���3Pb� ^�t2o�����x
	;D���k��F��88�b� ��ev�e�� m���I��x���O�f��W���!���2r2����"|���؁��-���o˂�R�_�=j�ol�s�g��l������DA;'���G�	My������A�%7���W�@��=����"�x9��F���?/޳'B��S0�e��ϋ8��V����m"�Ű�ݑ��X�{S�G�1������"ty2[0urbiV��aR��������'aZ=�#%R�ej����[�,�a[J&8	� G{-!%�c��j{[���B
��PZ���o~�>=�S�a7
�����i�Ѡ�71S�X�\T2W"�%s�~j�z��Sz0y�zhhA6�#ar���}���?�c��i�����!G�J����@��~������T$�~Bi1�X�������r6��S�BAg8��F �����m�_��\�Z � �7b�j	끠���D�0�����Lr ����?:
;81���joc��ǋpf��ɳ�abA�����Z�+\�	��f$��Y�
�N�H��� �\������e<L)����=�m�*��+��;J�]�0�/bc�)�ժZy3��8c`����յHv���/�o�;<d�ή�VgWe���`�,��@�����4������ס?�L�pY;��ޅ��+�r�Dx?���*	�I��s
p�$��44%�zv���ϛ�Ә}���h�&͢bR1��P�˕D ��l�&o��I�ObF)3����d'�b�(CL���.�W�C�j����솞�_ʝg�"����پ�������3�˕�5$���iA#����D(ƓW�`,�[ܿm�-��*�Qe����-�����>��?��T˱�dD����t��ZJq��d�Z�N�ِ�%�;����D���O��ܛ���(�E��ҷ��g.����L'_hx�Ѽx�4�Kbi��;mǞZM�����[�(���Q��!�|���@,-(zI��4S�F��k���2�]��/����we5����70݌S\�M�*;ozS��\���W�Ej�H66���i�×�(CY��XV��e�M��:A���c^7��&�����G�����H��[�׻�ru�0�(Z@ae)��Z2ׇq&qC��=���T����g��|�ͷ�7���p���~X��k��X��8�xǄ���Ë�W�>,ϻr����-���ק��������Wf�7��E�g晋�����^�j�dO$!���nD����)g� ��%��	�,t��z￭j�v��M~V�_��<�o ��F�R�c�:q�(x�R�ꙅ��H��x%�����p��-E)��ۖ&?�?��޲ ���ʩ��Vi;� ����P�<�?���������E޴,��c��ě���M+� --j��K�{��&�6	���E&d8V>���-�a�L�Э�7�U�$Ubr�=R�^����s$��N�ʻv1�8����]^Z�vjA����?nG�y�N�1��V�<lJ���M�����iׂ�ʕ�o��P���F; �M��;����NuH}�� m�H�=(�W�A���􅕍_�!qf���6_KĹ%��h~�(�U�+��Z�b�����Ǣ�b!����x`Zn���2�C��v�qF`"r
.��5��%?�Jܩ<6q)�(�	*U��g�^����:\�5�FW��.i����3+<�<�����K�}��^�k��ڦ�`JC��R��|��шA�.ww ���^H>u��A��^m������%Rˏ�@Ի�������67lȒ�p�θ� �u�,�����$f��/6IV�/�x�?[��jU��������}!�����|��2�~4���}&���=����bY��3��P�W�g��'a�~-�Ӕc|K�&^gW��ͷ����6���е�FZ퍶y�	:��vʣo�?�-��{�;��Ei|]��g��޷-{`Ի�J�
�G�a^YjN���/�Ǝ�3�-[d�{e_8n��i��7
��K�}����f���u�`��V��:�B25E1��+�N9���u�����\ `�d7���i�a�;$�P �����J,(;�ؗ:Iq���Ӭ��)����u�g��/÷��`���2�=��2���eH+��H�K(���`��)ܱ�O�;������	�-K)�rj��X��)���A������t��
��"����P�)�P�ߘ4�����߆��,��-�A�NY�l p`���a���Ц��"`"���Bo�͎�H��0��`�e		{�|&h2�A?F�����A﩮���K��ʑ�
�Eyƾ�_�~���K7G'�[m�,�a�X�P�+�nC:!	9Y�Ġ[�$�(�󇔭l$'����2�D������WA&�ِu܀;��a�.K/��v�L�B�M{yz)4h��ݻ�"J�����ɬ�d#��a�x��"�+��-b�������gv�
_���X"�.��T2��e�`߳m�K�Q+X���ͩ�ͅ-�|��kA�wF�d-�����6��N���{o�;��a1���v̎�u1CsKw�?�u�vt�l����+�,��k,�`��
5|A��[#&�"�|�E�f^p�_����nO[ͶOAlU�Ã�m��y�,ӱL�:��.~�4.��i�n8��tl���Ƃ�d%u�������])H��g��ҵM�c�A�&|�:j4㙃	�zW�A��C���y���\Ėf�:��s���2�N����`�>�ceD��5�`�-��dY��eiز_`-_\�	�{�����������Z����N��u�V���v?]K�����l�B�|�K����Ү��x�B���MQ�|KA�Rcz]%��d)yIZy!��T��	���Yã��$��z�.)��#���¡Ǝ�����
aU⤌8��ĳ����R=�^o���z]&!v`)���๝$ͼ
=>�" �F_��.�Vz��[�ةv��7�:�� �G������pxx�z8�3ҽ��h���綠�]��6�]������ к��H�3K��ۥ�=z�N��x>�z����Fэ&����I������"-��1[��a�m�Ns�Q*Ml|̛�#�K7V�6�K��B�`�;,'!|xr
+qhX�d�=:�[�Bt��J%�$$;XBt�`��`5����m�ǃ�%�#V�k����ß���߳P��a��egW�<�2�	0V�4��]����+m5����˞��ч��O�)|��gZ�S�4T�� {�t����ȣ�BwL)��X���4d��P�-b�4��#{/����/����<K�������6�T�U�^D�vh�g���~�Y���"��w��J�l�S�&�Z�m��١J�,q��E�N�g�����S��H2��JG�?��E�I�'W���S��n�cK�~���g�=�O��í��^ƕ�?�}�� "(�j�W��6�t�2_��^������M�Ы��Z��2������+I�ISN;�i��W��c6���?��g{�I݌Ďe:���������t�OO�-l�n�A��`4����խ�q#�z�ŋ�o'ܭ��������wN�`\Y���!�uE��wA����8�OA�GӱN`��x�H�l�X���xp���(	?���f�����"���c{O������ X�@�m��L��n���*<�O�i����?Q�Y���9Ú��lTD��p�R+�ܺ-�7@O�훹�H��a!O������|/�+�a(G�=}^�_���9ާ���	�4S�wwãÃ�����ˇ�?���#m���eE�m�ފ��[�:�H�`*�)[4�3F�s�LXd�*�cv��b��fc���XP����x/\���:���#�{�o0½���:"���oe3}+��x��cz��~�}��	Y�d,�$����<� W����N�O�p��س�Z���m�R"!��z�i�r&�{�:�$
7�f{����f�wP�ǰk�H��J��O�z2��Q^B��� Bc����d���:�Z�2���U�P�^6�ٛE
��do$!�Ҿ+������p)���0B�>��|��{�����mۍƮ�
�2���)"ڤ_�����w�U��ؙn��Q�bCkk嗲g���?�i�ۿ����$S}�i���K�Rr�����6�;�{�!9�����{��)O��e%�a�pR��8���*+��m3/mQ���Z�Y��[-�Ȑi2S%c1R��P�t������<|j'<��G�{2���/�1�8َ��q�\�ܕ󟝠�H#�,! 6�v�T3���O~�_�� ��o���?}~�ᙀT���0<{�w[��}��_|v�v5���������s���3���f�,�]!n�N��DM�Ul�
���8ً��lE��p{�(P�92_'���Q���
�j.nm�i	V�>�U�&�~}� rrr"��+G�G��H�R��Oh�/}�K;��s��R�j�tϬ�+=�e��	�����"\!�E��l���K9&(��j*H�2i�DB�`E����]j��J�"u�idf�qi_;�p�2�Kۦ���{�r0��?�u�>��B@��u�3�8K�mH��a#��ƺYt�b)��_W���V9��vZ�.^�)�����?��ki�"`O�L����6H�P3�tM'��g�_�?�Du �["=����x�����@�:׮� ш��/Ԕ��3�[TC���߇37�f��#�֠4n9�z�0t��[�gS=�$�Ӱ������=[�D�G��Ã>w�װI(/���<�xj���� \^�u� {���m~[�w�]$a�8L�JY�VN-[(s� 2���k+ ���j��~�lYH�M(_%�l#ZVذ���l(�f��i�v���;	�8x>��0Zڎ���Յ��v4t6�I�dd:��D��Ch�ϱ�i|� ����+�a��W�5�dN�r���@l������	�ʃN���&�D�(1z�A���'�Y�88���~���$Ev.�n��X�¥�	�
+DgV.0��~�����]���m�m�saT��ML_e2+B��"���/�h�%o~z p���~�����#�B�&H�']龖�����`nJ=�!#�Z��I���lu���ߕ�S
H�^6���|�9����7>�*�8kh�
�Z�o��36�
�R�b�~'=ec�/�������߇����V��l�:{��m���Eo��[�-��Y�RX��.v���B�6�m��?*q#�g]�|ǲ�����̣D���:�,����YP-~h�;FN�VM�^����Z3{7��S��Yel��0�lc?yz*�d����eH[���#������T��Iuif��##D2+�~��(l�B3W��NB&,��I]\?3���8���]�>w=N��/���j{Y>lG����L������3�i��>�Q���Ǔ��+��rq�¾f[�ھ{�W�|y9V���rնd_hV)�p��� ������U*-�c�����`�������0u�Z��1�ڳ�nd�?��􊏀��s.QB�̩��Y窔Q��̔`�i�����>׵�����~�� "�:�d^Ft�DV�ɓg����w��y�w�G$��a:�k�J�2K�N�3�59u���	)���~�ݶ�k��Y�����t���l��0�^T�Ḣ�~�%fg���Ǽ����
6�ʿ���1&1������o������Fz�����|͉�����{�"eA^�G��J���d�<�k+{����ׂ+�@�J������D�;�s5.��P"�٩س�y�������!_��������(�aO-�t��ԕ#8;��!н8���}�/#A0C�k���v���'��;V�H���L�q���&�0�t��N�����5�#�:#mQP�"��8��Z�ġ�xj�|����֮�r�ixV�k�w�<��h��5/ɀ�l�{���E�P4��:*����@|�M����!eFF���ϩ�U��\(RfW�h��*�cY�Z9咙�p||K�l�ސ��L��r��͎~/�Q<s��Hb�`Wy��u�aE�#�a� �`�֛߭({�Z)�w�oL�J2��5e|UHj�M^D�,�BR_ę��w��t5Tp�r*�y��g����	r�܏Fǳ5j��uǺ�I�1�k8��.�9�'w��*7x�ԛ$�_ja.��"$�H���c@YI!VQ� s3mO�=�IH�N/�J�zuO�o.�Co��������w/�G�7���H�)�����]p����+dl�cMQJ���w���Fോ	i��ҤiAC���M�L.�w'�ak��I˩G4��It#+��6�x��-�3��ƿL�#[�R�`�׽�w5x.�oM%+H2�{�$��RT��j�.�������m���8lA�{&�!r��ct�З��Y�P��P�p��&��g��n���������b��C�?Z-��&@�`���q��h�6�2��%7��y>������3G����r�Ԉ\}->7���L���.����f��B�1�!��l���j���$xv�tVˮw<��`F��-��b��=�Ov��(��%T�/����流��L�s̾�:���"�eTk��^���5���f\�}-��vlc�ALje�2�fjD���;׻T/en�дb"�U�eB	@���p��õ�ڏFЪ�
E��<K>1A7ڭ"�S��Ԭ3F"]#e���1b�i,�����[g+Ơ��,f5��ԌB
����PV���x�z�]4�F6�HX�ET�JLcV��lK�QXu�7ģ�
+����CV�R+S�#ae`��pz	tŸ�{1��@��N�l���t][
�Z�Oi�
ҪӻM}*���^OB���L*�t[�[$�=����2̆(�q�4����n��V9�������\`�ж�!���t�g`�.ŸX�O�&9�%#��5��+�,��]�����]�U�Xbʚ7]i)��Z�"�	[��d��
�E� ��*�	�2c��$0e�Xv��*^�,f,�����d%�fQ�z*Q�_��g�~��ү)붞������lJ��v�1:��4VJ�����Fb���V̔CWR�ϳ��C6�'P���F��Oa2��Pr�D�B��#���`k�@��!��f�n<_���&�`�GV�.@M���(g<��S��`��J`˩Ț�o4C9�X U�$��3_ n,-KCQ�SԈ��h���:������N�O�\*����tnѳзal�%ӣ�h*�m���Bt��=tX0�Ӵ��e|0)���L5W�B���in�<x�$���j�b��\]L����U���Q��-���@ı	ε3)ee�,d��MI9�W����reY�F�tη��؍�-&�b�Z��@e7�v-( �8_6t"��;�!wXDR�ru���'�:�)St;��!n��
������I�%�|��%�F9�k���\�=_��=�c6�����%���
cZ8��Q�A'���V���,9A�(v%�����J6#R>��6R�0k���d,�е�<��++�j)��b�����0���$'�����A���u�Uu֒Qyc��H��Ԙ����0v����ك�w�x�)�E����2�p�,�K��wE���]���o�Ǳ�Ǩ�Rn�Ti9����4��� �{��b�$��*��7�I���#��+���OF���WAB'o]�"cSiU���P�n2���	'%*�ci��T*���s	9)[h���)�|?Q��':d;�
Mw�dJ?Œ�5���ɶ0��~�g�#]�p��R��CoU�g��S-��u���G��X���B�rBh(��@���e$AѼ��2)	x��e\tC��Ԃ�!S��g.	Hp+4:�j2
����yU�)1�<#��]ƴ��B�Pb�'�{�i ʞ
���M>d+�g�S��	�7��}�岫v�6���� �����<�U�Ă�<sH�SS���p*R�n����F�F�ڛb�f~��Y�����|�{�_>{-!�˹�oUKA��)7��"� ��l�HX��K����`��,"��"��:f�������!�x�2�r�6�;wW�����ꃞ�4c1삼g�9�x�:<��Gǒ���s5�	-[S���
w��C4�q)�"���䞞7�?G\�-���:5[��~���Ŀ�u P�H�K�D��ڼu2*�ϗ��3��ԏ�X$� ���`���`AH�)���+9���~�0f��>�V�)'6������4�DT_��7�YD�VW;��j�E�]�{�Eh�>I��r%�Rj��4w��":�{0���R�y�N������ϢS�"J���)J�EK�Fg7fO��4��#!>���E�T{�	�F����y�u"���k1�� �*RʋU?�g8�.ևL�:���6ww��U���61����h��_�k������Q�����x�I�"bn���D_�b�������̉yXp��卤%�+2���-��C�[y��4�d�ha't5d��#kȡƤ0 Y'��~�*�C������H��8�,"%���2�7{�����J`�N���ҽ��y	����$���LZ���ݷ\��⢽ޭ�}"'a�<��1Ƚ�tF_h���J�KpXU��V)=�ؚGS��=�N��7N�a��?P<�X��ݎ�n��B�TT�ꊃSzVӌ*=HM�(�4���7�������a�0�}}��*d05�9��&�tC�y���麤8�����Z(4X�D95�Y[�)�0�au嵬��nc�(��(�2�j{M�9��b��i�RmN�6w�,:�@��u�y�*b's��ˆ��H�#��d�ƪ4=�����E��R_0-�FpRʅ7�����u��{���e�V�Z?J;d�G���2wmKe,�;�JA���,$�gc�3w���G� 0Q��pN��ͺ�f�u�l�<p���g��ۃ�O�n�����|����ɓ��嫫p}3�pT�l�V��7���fK~2�ŵ�������F�`oǾ����[3p谩ir�iB�5��u��xLp5�.M	��[Ǡ���N3+$��,,@�~%cSj�K���C2E�EM�弭�*{����w��/?�,Ba<�ѷhxP�� ���3���V�ᱷ���Y8�6ò?[������D2ө�{��UL�%å�� ���,R���ǅmc7�V'O�RFÝ(�C`b�%�6��/�������}t�#5��.�7��H�~���k7s�@�1T����o'ľI�W�Vڲ�]��A�0sS+&-��v�Xo����$b��j��ͪk��"�A���]�������v;ZM�����ō��,{ϭ��V�k�e+"��j���8%/��z�E,;*;��pt���mԛ�L�g��)�"�e�D�\Yk#�ѳY=-�j��Z��}�h
�y9؈��є�t�����e\;+k���#y� 0$��J���X�ۭ��m�������_�2��u�W~~��߇���4���GN�4�Rx�P�P.�kE,gǙ��=;�)�#�H��{���.�j
�}Ӟ+�nLx�-k���ڌq�g1`���L�z�U8q��K։v-ϋ�87��`��Ã�kb�q�������(fR�[ŉuc�T��� �W�ɀl��G�E�n�^��o�|�L�c?l�i{;,>:]	5�fj:�=�������;>�Ϳ�ﯪT��Q�
�ƿ��G]u��r�Ԃ�r�[YFztGSa`��F����\�ԛT���锗.~�d"<5a��Ώ9 5^��嶤(j5�k+㣤�M�Z4�es�1�Ẏ[f�2#.	�"�&�i�����!��O]�5�#����Y�Sr�=���9�-.L�H�G8m�����9�����1�'��h�t�
��I��ҕ�	����`"�U�|`�, 5MF�B�������}_=(/�f��x���f�����_2�b�e��c��Ϥ<�c���ݻz�|���������K�����Q�q����oFH�^ߵQ�y�E~�Ɍl�L`�>�>���Є�9��z{�(�������c��������){�5�t���2|��'B�.����Lۗ��m5#�^���*zl�Vl������c���;����aw�)vcg_ښ�^H�i�6{&}�+���S�B���\� 6��ϥ�v
"���!���l�Nq.�ڰ��6�i��}��Au���lk0Oj47�O�8{�.}p�^HA.պ!�����A �N�V�(��˕�B7�2&+t�K�"�
ؖ9 Z����-�x�h��d>
.c�:���*�" |����8��������͵NH	� ��L:c
�z}��_|!:;��-ǾNW���J�{�����ko�^	�KP�w��y�NB������?w%��W#��q��Ag3o���V�U҂_�\ 8>��,��I2��X�_ ��>
?��c�Ʀ�t���zHA��Ҟ�������ĬG����/�w��e�6�k�@���?Qp��8w������h]mE��7ɱk7")�Z��R@QQd?t�JL���_}>�𮐌�6i�F���R��*f�Q�-��_6�NxǍ��c��o4���6���0�5zOa�r�Az|)�e��N�:��5H.��j����b����+	
Nj��Q%}�:�h&�bi���)A��wQF�j'C���=�e
�v8�ӏS�^#o؆�K+�MN 6T:��DO�^�b�9>�h�Fp����L�x��6��|�˗/mC^j3����ܱ2��p�jW�Uu�-�W�#`��������4)��O�[����q�ܟ����u`cZ١v���9D���ۑgq�Κ�պ"�@�ՒuE{�q�Z� ��l��7~r%H�+���a�)󹞖ԫ�o7��Ah3���ǻ��mں�{�u��ۑ��e*�����X7V�b�o����R� ��᣻������n+P|!��W����C�h����w����,
�/yS�5l|���Uת5 ������������o<���ް�o����?�i�ض̪��q:����_/�S�uo�8�~���S#GȮ�i�[+%���zz�!=�����Z-��l�o��w����x��N#<xxW����9j������1J�~�0$Q3Y���h�v��Y�^�۱��Y� �G����G����o�M�4i�HA#�F4)O�t
B�뫍{�����7�b�(Sol�������o��������{�G��:z������o�t��2,������ҿ���]\l= �    IEND�B`�PK   �EXr�>�� � /   images/b24f041f-17b3-48b1-9f28-cb1f31b050cc.png�gTSk������H�o)қ�4K�
* UB0��A�J(�E�RUB'�P�I�ރ&�jh!��Z�����1��{~|�Xo����|IB訝?�v�����}�m%g̟��'�_~���p����O����s������\�����Mv�􁇬n����m���\���p������ճ��b�.��k�lTTQ�Cn?�LY�rp���M֝�VOY��u���h�~f�����y��$+e�%+��2I)��ywK�*����ƋAg�?��+t^.7�.p&��NG��wg���~I$�_��i�"�pw�e��͈�t���47w��x�[��� K��ӓ6������Pu��ʏ�/���Aa訨,��x��
3�Q�A�4�ɉ�U�5F�0`}��{:p��$�]��I�ץ"��' 5�x�!�A=���=����_�L�M�Jj��*&)�~4�Y{�o������ }@b��D���!��/�+�M��u�5!�;,Fə�@7��jv.���ɛ�++=w�-Gx6�Ǎ�'���HQNS��:����>�gE�3���Q�Dha���^�-0�[��U�����/�a7�Z�|��d佉	��޷AL ������&�`HU�9���?n�}��!_d�Y�9Ҭ�	s
<�w�Ԕt�h���Ip?���T��.���ͽ�W�:h��Ճ�P��X��o�N�^��n-Nդ{�b�/4�՟��σ���zG��`�����%�&���oX%Y�*�!)��#��J&������s¢zG4���%��(}�����GY"�G2Uץ<
Y�H�Gh4��'j��J����6�7]��	�&�!ٱ���u�����Fc�4i��4=�1Z=�0�޸�/�X�X� @�F�����Z�W�q�8��ya>pO�7R+�Щ`cc�ű��8ȹ!7�ly�<)'iQid�LRc���NaUa�7�Lړ�����#N�U/dX5M� ��5poO,��w����5o=3�奚��mm�U}4),��Y_���ܳ�ߢ�"dе�F:���㴊�z�F��U�E�0t{&����D4���M ����J�;���x�ϑ���]5SJ�7���a0�Jvc15=�or�}ʅ�Zٻ,�*���}:�Ѐk�^��~:U!�1���W�Y��cuV�`�J8^�m9���@����tЛ���8q�v��7+��8�����)2UH��P��@vE�v�Л��{��}	�%0f�H�"�9? �L����{6����n�?g�\�:�1�#�{Dt�f����g�����pI�t"��۽���d�9��H1��`F�ܪ�迫���>�E_�y�5���tz^����s>5�5�q�^�0߬n�u��k}q�*��[��к���,(�7�JɌ�V^x��a��^��MW�Pt��R��l���Z��,���e�-�I��M0�.�����۫,�c&��*�C�9G�M�;��v@(g�rw�5^9���7�҉��H$RRq:�MHF��c�?���Hy�f�X{�<�!�;��g����\z�nvj�s�ժ��*%��0��+��I�������z=F#33�����Z:�#��*�x
>]�0�������C���<g��6D�1G��f]�$��>�����K}�|��v%��O��:��L�|��r
DĤnԎ��ld�Y��맑{�����ޔ�T���Z�v��
�����2�̶�ݨqFάP�ԧY�=�܄<�|')1T�!R>���{�����0�;����K�V�����<����	rq_=]�*����n���*'=�Pg ���g�~v!�y2b=퀕.?v�ui"@P4h�z�|�j�Y�u`�xvx����<��e��GLpo��n����5���V�ꢃ:�5�U�H����O�UN:�O�_���~�)&��Cؗ��&N��.��RsQ �oe�^����h'5}�k���?AC�!���a���'n��i(D��*���H��Q^^���x��qu}w�����O[�Fsz��ir��&�/%����x-q�.��D��!�,���@���= ��|ډ�f�I�׬h�)ĂUI�\K`%�*�1?=�UL}���4\ͅ �~��N�����x@ !��)���}N��z>�e7��>D��19H��md�+����8�ſ`�A�#��#��{�CY��/���!b����[wÂ{
�,�"���د˛�dQ��x�����0�*�t挃t隒o.R ��"�WQ^�6��6���u~L��4���:V�B|KP�����55�7�#�aQ�}]ԇ#�kY=��q�R�����Fh��❷j#C7kF�, U��$�_4S�������wF����ۋ���4�G�iq�:󪲊ѽ>6h{�eF��V�XA?�^�c���^��Cʁ�F�.x� ?Yc5��2�V��C_����7�`�RX���(���Qz�����d�7�)q��S�4���GARzz:��+�����#�j���몚�%Y����a�I��*�`��1\�Y�>�Q�IM�:�U"��Bkٱ���.X��bow� �������������� 2�|��=�B�ƹ��wU�k�~�����x�������_��B��H�A�r��¹��P�%
�a�S���NN���`e
�4b���AJ����eI#,�q�;��������<�(��b#�[g��v&n���j*S��	���
;��V�ubM���w��Mi�l�2YW�:�Sc	�����~�i�}�����xN��U��ѺQ�c�mV�%�4���ƪ~=���@"�I�/Q}����
M���x�2ɡp9)
��9����TĻ�:)��(�$�W��Daa��+�M�A�	ѳ �~���ď�
�"WC�3�z��G���{��@T̷�~���}��6����JPu�C�Nܛ w0�76�:�`?�Z��x;�Ta�W���"8�#��ȉ�)D�<��uO�u���c�B�u��%���XOJʖF�g,�������*%b��>��N/��������N��HM�WA�4��M�n�H�˫��U��#%��=(>��`j�S�Dd�]4\�K;����U4J/� �6�# ��x�{ͧ�ۋ�<v�����n����vuu�ۭ^�w��v�ᴗgu#t��l؛���fұ��$~�1�ytMC��p��M�ܴտAx-��{�i��8ֵ���������B䳣G����߳�(�; �!Fft� .?��Λ5Ҕx<�y;k|s���&^R$IQ���"�������zz��"h,sn.�C)�d�����H��O��X�0 N	)=�%��d�B5?w�Y6+�N�3��I��2c�q�05Ymԭ�F�!lOR������W@�X�t�Ͷ���ۥ�U�R�X�-���B�OVL���6��ᨆ�
le<K��ӳ\�����_ZZ�RϢ�F��ue���B�<��Y���'��{QB�\��&}�Z�oա�Ǽ`�Xz���P�KZ��@�/�4S�����3azn��sd��MFg*aYD�pZ�eP���}��97��t���y5J.3߬J�P1*�k����t�0�Fadg�k�z՚}1�=tӽ�5�v��<���/�0�DH\h���ù+����*u��u� �v�	��X(=�G=�x�<�U�F�2Hu�l�L�O�{A^��@�'�i;��^���9���t�&=�cK��� W����N{���,�~���J�G��!�C���E��׵Y Vw����z������ĎVY�79�'����k6�_7,f�M�"���u�<oM����$�<�.2��Ë�l�(��J�̯��@j@5�H�DO��[���sp������_ �(z�� �?����]�=;�p��un)a:ƭj��d晴��W��̃�����R�r{�\=$qa�ȿ/�~d9�%i���6����ON�",-�<�&��ڬr�mU�7Ψ9Ց��׏�I��X���ǻ�޹�KJ�K�X�5��2 d�J��!�
F��a�moDs�*Eێz�~mL�/��w׌?����ܱ��t��1����!%�As�����5l�j��f��ڬ��>��ƌN�Ƌ�n�&bJ����W�3��[7��Q��:J��\o�-�����,5ܿ�D�m�G�Hሂ�&����I��G����(��X]�C�Y��FM��ВIzzc{�j#?	�ze�u|�{���2n5�CaZ	�*���uϞ��m;u��Vf���[!j6g\ax��1f���J bwR��iF�&��f�pd	(���a���?�.��_�Ά����{f`v�Q�3��Ī?���>Y�"�;�h!����4�}/9L(�-WHs�O�b�8���]� ��u0n�-o����g��oZ�J��x[@�i�ajJZEO��0�:�b#�����dL��Uި��"m�?#�<W��`Y�����՝��}�0x*/�ͻ�2]d�Z[C�c�/�Q#����W86�]��:�N��L۸�w^����f �7iʃ5 �.���쳳>�L&�E)���O�x��̥%R��c�N)��!d�kۛ��P�?�pt ��+G���L!��c?�U�M)Z�>�K"��@[^g#���X�iM]*k]��DD�,�ظ��!��WVt\>�I#���[�2�?+���u
}
o8<�[��S��>����m'"@�g�K.�1����B����I$���RY�|�f\᭸X7�:��WFa��(���]:�� j?���~�����G��e��^"Ϥ��? ������y2z����M�ˢ�+j��Q$ٓ�ha��b(1M��Q]�I�t;$$=�NQ�~�Z�FW��� "��QS���N�Jð�l�%�*�X)~�*�q�W����ܙ�O�q�D�$-��N�5q��dk��oV�������Y� ��|���
��G��6�!im�+;;�t���*F�="$����"��̠��6����ƶ��ĥ�ɧ�t�n� ���VR|����������J�Ϲf]�X����G���C;�G%����?�;K��O?��6|dy4���r3g�;>��f�2����$J�zՒ�M�d�-d�q��.�����!�lYi��=}��{`��v��v��(�����H;J���'<556W5����{si��駕Fn���&��/'��u��5	-�F·������?�g��`�_�g-�;�	��H��U���Q ��^5ЩE�
��/.�o����'9����>d�א�vr*�}%l���I��@�zP�rD~J37��):a����@fr��e����������w������?䖿�� ����m0��J�a4L<y�)M��qc���_'2��[�5������>	�]��j�޹P�쨙�s!�_�F�W�s.�|�����?�]v�{D�x!�N��H�)�DKK{�^�&n*N���h�=���$�g�|��ύ)7�.�������{��yQ�nY�eJ�P�TP��.U�U�g�W@K�z��z_����w܋�͛?͛��̤�[��3hzr��U�L2z9�[�Ϗ���as���Aq"�`�q��>6u>u��#5�
�2X�O��>����h�*�*�W��߻�P贆݋I�C?z�fL��X�sC}Sna��to8�8+Xɽ�A��\En�ʄ0f�gG�B���U_z<aȠ��cPs3DƮ�5�h�r�}E�{�	�ꎿޓ4�U��j���=�������?rZ�a���ѭs���iV�W�����lFDN��W
H}>��\a���`��=�I	7�x`w��_��U������뵳2L������'�+�w\�٪T�e����[����W�z��;��"�VE4%FDb��?iѮ��xC*��g��z�h�]�pn0��=o���i�{��U7�TQqq|�LJ��۽�K-ǮV���ry���o��+�u��h�D{���?���7�zo�h�j��x_�_�ϵt����~Th��Z�����ͣj��="v�H��Tq��z��k漪�<�����b4��
�w����f>h��֫~5Ȍ��g[lg�0���WOnn�>u�̵�h?x��j�o��*�C7u�f�T4xc'��/5SvcĹ�Z_�%�L������A-����,_kn�_�e�O���L�^���"�{�S\bmv��h�1͹�� �~�v���3�i1�'���l��l~z����.�nM�u��J�G@��ݏMO|���H�f�+8|�^[���K,���ӡk���1���_ھ_�!`X�.�Fh6,�(dG�G"Hx�ұ�9����C���+;+��O�""L������"z`ߎ�E�`_U���^"������u̼�B�#���鿎m�u�.[�8q@}�:=���whb�N��V7?�ɣ��N?{p�������
��(t=a��m�3�/L��}��V��(�s��"}�^�ıe����՚�PU|�ޙ��1��t���0����9��ζ����Tc=!�?Y7m�g�R�>>��fڨ���6e���r�8An3��N{�̝חr=�_yȽ�	��q��\�t���r��1+�8Ё��(��+������,a�{�X���\զ��ߎ5�8>�R�c��1���N�I��N�Ѫ<MN���D���8��.�����Шf��ǥęF�G/�!�<�̹�ǬK�6����y�
�Dպ�r�:ҍثs�֨|:��ZT�}2��-�B_ZF������Y��6!�ֹf��|g{m{fǼ����kRaN�"�n�T���f}��KZF��ֺ�����dW�����+M�)�{cm�T�7�wj�E��a?pVb߸K6
�%���u�;�u�~�Z�����-$ۉL�
7;��������u�#�g�Z9VLnt�a��+֣�T�G�s�b��c��hר��ԚZ�h�g�yç�}OU8�W�[8ȁݮZyY�e}������ރ5�V��j������U�q
�'$k�{|��N8���� N�d�����{N���z���V*�3&��j���h"QypȀ�)�]���1�l��?��{��ɤ�W�*�\U1������H�}^��XO�b�A;*��vY�V�?Z˭�fԤ���;����:I���Ѧ���V���CޫIF�ǙO�Lt]��\�
�_���a��5��Eu>��k�
ǚ��3Bj�>θ���>���J�~ϩ����k
��=L�șઝo�ǔ��|��򆖧*T|�K�Z���E}t�q�t[֮pZ_^4��'q���0��Y����G	)�
i��f��}��}��{�#��F��xb���1J�t�S+�� �{��'�h�]���������+B�t���H��`T�0����b3t\8��O����K҄�4���kw�zjD�qV�hlLsVk�Wt[~_1�B����'Zm�ȯ��;3M���y,u�yV_���8{�`���k1�Gg����ś�+�z9�ʍ�o�0�s6�N�7�ä%�z���5�BMw������r�Q��iP��\��S�q��2�� �C���Z���@��s5��aڡM����,���#�+�'�׊��:$',�?^�>ܪ���9w{���d��=���q�6����o���8�����i���U��{$�'���e��\/#{����1L��m��ð�q4S�~9ͩ[3�c092P!����ʵ7[xv-�y�Dc��k�Q�mV�3O�v��������-&��Yу ղK�����)��)��/?�z�*�щ	�_L���o������s�E\�I��ڒ8�r?�uB��XF�����J�Y�����6�te_�\�v�}5i�ت�3�YJs�p5��v51���Ho��=&	������N����,ګ�>��-v�w�T}�=)mڔ�>�$t@Ajw5-��y�|��HX�F�f����=��%n� ��z���4��[���s/-j���c�͌	��ֺm�M�F5�����g૓�/��w��n�E����WS���c����p\�S�ً�t<�/o:*��=&��v�>J���(}�b�pE���s��B�GH�Xo��l1�Kիxyy��n3�^��E�����c��_�s���N���ʹ_�.��W�Z����K�c�}]���\P�}/Z�k+�Ć
�_9�fvE]��wT�$�91ϰٍo��kj��s���<�vb��e*�&�=W�1ȟ���]-<�Ү͎�2 �Ē�5ym�Ѫo�1����_$]��c;#;?���c#6�rsp�k��i�4�-�ɵ�I��G�k�����1d�{V{5Y-k�
�`��<��)�mr�I�~Q�Be^�9�9:/�(> #*�p�p�<֋�\{eS���S�7lO'� z|�~����>3.�&"�q}6�x}���lpr��+�ڐ����Ne�U]:���gm����oNhVU�f���A���%��;>����䙵m���ck��]���S��?�Ty�漏ɷ���0��8@M�`�N��@ ��G�����{
H�9�h>KM6oV�賀����^c�����>�>a+�L|Bqр��$�������:�ɕ~uִ��9�Rآ����}�`��q���<��^K�ȴ�B��Tb7;�8�k�]'�%+��]��%�������wT�T\�'�e��L���E�J�4GD��phX����#�z �qn�{;�)qz�}�C
h=�Ɍm-)�v�Pr)��V�鑎Q���$��ȽRcG�x�枛��������k�4^�{�ve��|�_�'���"J���xj��F}^�CqV)}�M��rԛmL\ov�^�)N$���Vu����L��D��F��͜
�05]�r�����K(��|�υ���F��=�"�3��%��hi�8�ū��n���kKUp���P����ܣ�}G��.A���"�e�(,W�K� �����H�~�N�:�����S���Ee;��l��F�I�4�WO�y">��	��$| TF��yYe)�2�0т6$~3�]�I�յE��Z�o�~S��sũ��"���	���G�/W�p��}j�H��}m��~�Q�i�x/"��j�䨯e�Ϭ�.���)%F:����rk��֬�&��r���m�ĂP"h^�e�?�f}�|� L���M4Oymg
**�l�;�V�L����IeqZp�gX��%�l��)��47��}i�����4�,�S���>i�>m�>e��-���$���*D�hAk��g+��rh
�m��~d��M��rѕ�j�5�����L�55Uj�/n��P�%�\X׉�Ѳ6��'��/%NY�������E��=�~�`iڢww����L��W�|�B�j�_OR\1�P��G�����?�>�?����Q%3�S�2NB{���!��4q��Rо��[�3R:g�<�_�P%�~��������������b�~RK������A6��iD޺W�/�r�ѿ��%�F�W��3`��3�y�ݯՋ+1�
Sу�꓿n)��H��
չB����BS <��q�J������M����K��l4����I3h	��re״b�X�ۼ��ü�3�tU�ա=�,&/�з��.:��b���f���ѾA2aS)h�s ���C�J���Bű&��ا���"T�2A	
��i�-�4�-���zJ>_����m���9��'L���8��@�^��xk�i(% m���V�=b��jٲ�%�D-q��Ep���g������f5�Z��ĳL ^_�<|����,s.�R����Q�%;z����aht����ě�E[���5�K�K�W�s<���!r>�s���GV����o�]�v��fwC4{��\�w� cH��X ���Ĳ�Am8�{�<�(ThU���ڰ�����˭���7�;�r�x቎�%�Ez�����*vU���'Zv���aw�Gp���^ʆ�O��k����^�<��
T�D�_V�S�~}���{����)�j����K�:7M�1�5m �P�&��-�`�ok��rv~�"�!?��h�l�:���B8�­�/ʤҪ'��լ_�i	P��8���D�%Gb�L�&OZq-4?��3M��V��t�K����cW�E�
"ӗsiH޹ɶv�H�˱��c��^bɞ5iw$=o5R޼=��"{�bIa��*
�29���x#?2�(��;� "�t�M�nĈ(N����$������Uΰ���Qx� �f߿�oh7�V1ov����G�!��Ŗm)0�fS�E(�E�.Gp"�5��=;m4ڇ�c(Tq�s��t1�2���R������Ae|����ĭ�~��ms?p\���Ӱ�4V˛oq�r	����u�>Bˆ�~ey��k7}��7��0��@(��ߌLA�pf�?���2< o�P��gB��P�[�Io>������d��c0�̵�H{㸟��Q�W�n�_���e�n�5�5�9��Diw!��9R��SMM�ԣ��X>znfn���|�d�;Ϩt� �v3��n{ad�ɽ���.B���4�-,,�)}�}�V����R���G��&�Xz���-r}ru��"�2�����O�C*#�ڿ�S� � ����.�LS?�|�fzc��W��pe�]n��m�4OJ#��P&��ֺ��%?�����^����dKtNSIȂq��m4+#&oχu���C~��i�@��oF���|a�4���'ٷ�L��.�pf˘�mݯ��Y��u�7��b�s��.�'wYsp�(3&��)@1ނ���T2��P�C�̧�:˨����.ny?	������aϣ
c<��w��R�2����m��m��)O�����~X?G����]�#��+�|���%��������e�����}����o���[���ږ#X#tP��+ƫ�M�KmF]u�M������&z
8��&��6�]y黓�R{L��<.:�PM**]ˁP�ڽ؏�vC���r;�|C-�5o8�u��Z[|!��w��� ��ڧl�'�5���$�d��o�S�� 3ŝ�[��Ͳ�n�'�~Aj5NR�ʂ�x�<HA���W� ȧQ��]�w1^���IX�G�7��0Xզ��n��~󼖘:a_�
�Q�/W$���'�T�*�`T��x���u�g���͋p�:�߭.��Ŏj�����Sh��ҷ��e5�y�)��:�0n3)�O�
	_��J$�(�Z��_�����$LXd�$��5;�R0X c��m�&�23�7p�P� ʦ����e���"V���?��%�V б�L���5K��^�Z�ȕw���s�NRy�5A/�`�̭{�"fХ�H�v��ﯥ�J�j�9��r+9�7�ŒR~zN7=�C�,f 9򞻬%}��x+ܓ��D��65U���f�r���oxC�8�> �NE&�t�	#�<��|�g��X_/�ޣ5�M��	r�G�#vc.��ME�%ht��_�2-��N��|�Ԙ���\�,�:���Nl	-@�p�S��R��v	�
��� EF��� ���<�
����n�3E����WH��'ld���.#m���x�}�J<<��؂�O�/K�~jy����tP�_;0���L	���b@7����Ylӕ��<]���iSa�:V~���u��^�*��4א��B=�y�q���]9a@�F�в��{eܕ���%�7!2��J�:=�h�/_��D���u��x�h���G߈��Dו����N�Xo���(U�|f��VK &�7��%�IcN$͗K�p���x�"G�JO�v�s���Ş=K��Ƽ	\�sY�-���>����U\�;���,)JM�a��`��
xg����u�\~ $&��+.2��n�O4i��#4Ǭ!Y� |����7Z��d�3*6��!�o,�.���̕�� ����#Ϸ����̕bC����<0��6	��h�~�吻�/ۙ��I. �5��ȂzB�!�ky	��L���珺�@�V���I�#�B�3�_-����,>�?�������g6�zV�D��p��'�l�3hj��]k�T��i�W�4e�n�m~��|�Q��2���T�S�]~jX׫!T&���P��[�3��8]xk9'	�&(Z�m��0k�P�ԩ��o8��⫑��#��1�N��/�KT>��@7��#�)[)>�8#v�$�L���DPl�	�d?MEY����6�q���i|kԫJ�s	o��B��?'Fz�|u�x[[�Jh�9�
��oM���DT�� ��5��=��7���\��Xjm�.G���H�.�Z� ��#��)��	���z��1<N��hN���m*k��>yZ�P3:�wܦ�ޱ����͠º�}n��	]>pb%	�`�w��@ܝ��~��~�
֛Y�G���P���̳Q8�+��s�8�o�$v<=kW�9�Q~���b�n�x����Q^ z8Ʈ_/덈�.��u��N#�gxK����Ӌ��������ȷ�x� �d����ӿ�m��%�|��n'�qyK�h��A�n|Y?̜);��L�tX#��%8H)�W%L�fyS'P�s�odQ�|�eD+A*�ۀ=�[�������y��Z��}�������vD���� �� ���Xw�@Bޱ�p�����s�&'�._�B�&72LEZ�Vs���*�"�?B [ n�F��
4a �c��Л������?.��wj����Wc�;�Ŗ��r~\P̶�n~[>V���cR�I��R���� ;zPa����i,�.M�"���s��}4�x�)F��g��*Z�)u���);�E�r�kG�ͳ���Y&d���� �[(�������6�X@8M��ID��9'M"��+��G�s�H�9���s+��;눏o�[�� ���7G��*H��7l7d�S�y�����_�����*��vw;[=�(eNT����#y	+@����7O�� �� �����"T:�f`��Ҩ�2�ĨC*�N�0�/�kC��kna����D�Ȕ��d:",��z$6��'�t�q]�Kp�F:�j�(�:xd��v,tQ��f#�G�Z�k-$4��X�b���Z��daO����sT;FB	a1�^$ԣ'$����G�r�.b�v��mQe�ơ�e�<󏾻�S���Q��m�*/��J�4
�@%�3Y0|�O�T��5Tf�?�\�C����Z�"��ݩ�U�2;�	����s����ui�{:�Z���ɕ\��ʅ���u�-�
�����y�LMx+@�l8�=�E�Mx����Fj�j�����h����w����@��3���S�6T�@53���p��2�*y���K+�ۓ�*KH�$�@�0�)S�1����X��~*�	n�˪�{]��Q�9t.�g�V[�0��������j��۰7�O��\A�UPg�=_^�3��j�hDl$N��k���f��>�8
 Y�fZ���` `��I��t��0uўzr0i3�5��Y[*���>(�0�-���0�q"i��=|�Pц4#3��nW��c���gJ�L2;��\�I���P�>�y(Lƺ������V�qSۻ��0�a�`�r}�(#� Ʋs���g5p��k@l����g��X�n�"fٓ�'_���0���}M%�s[�y�����j��Թ���2R;�S4�{��HTlĨOΞx���Yx��6w�Z@t�Dv�aQT+)=���i֓�pC�%����8����D�����	b&\�=�l�U�ð@uܷ��uM@h�ܽ�Ǹ%M��g�����s^�@�mZ�_�yY.7�5lݼ�q����	��Y��M3;s�'�d�FN�/��s�ܢ7�T�A9O}�&
���\�@]�d7��bsR��w�9�C��&i�݇O��.4���VH��L2T�~ �fY��\�2���L�&�R=fL$��_��|��w�-�ԡ�(�������v��Q7��`�5́L3߅�@�f`�1&^�#S�x�w���a4��m�	�{�����<K��Xw��מsR%&��7�w%��u:�tXF?wn�Sҍ�J�aC70�A��͆f�hDE�<�����G���|�/~SI�E�l�U�K�u�*q��m�>*� ����CQbu��u�I3�C#�N`F��Љ����Dm�sм��( ����~ �o(����W*���\X�t2���4�tQ���kb��6gl�Z ������[h�*���_�H�Du�e�&�% 	�:��w���M��~��OԏtƔ˙���_��x���]� ��=�@̱�hȄP�t���5�I��{],@�����U�q�k�`k���G��Tx>u���R�+��R�.��l�����EB�?17j����om^kdRI�T�k0fQ0��5>���@yl��e�1�V���1")����v��K�h'���TW�|ŐG�w�XΩ�`ϑ�2�j�?�JMx5�
=Ӷvʭ\:�N:������g�|�7�H ޴n�u8�p���7x]� �^# �l`�^���;(���o��'�Or���%���pVj�-~�m�7h�{��M|�1|Rh�R[��`xi�L�Ӡ�4hC�=2�F������֐�֜�~avi�d`G� ��H!x�$g>���>�唋�
s�/���
��djMQMؓ���&��9�lfi	9�����DKrݜk��]ǥ*�0��ubhw�E	�i���*�p�&K`X�3PI,"=��?C��dŌˤnn�ܣ(t
n�� ���aKm5 4�q]jW��K�aM�|�1�7  ZPF ��|~��5g̻WB��P�����}�≘���O|F\_Z'�Y��:�(�a,"ah�5	;�������_��� C*ҭ�`#��$���?�c�[��R!~�hS>�=���M�f�����(�	[�z�/��dL:���� U�g�|e�`�ª��(W=�Ђ�r�둎4 �����/VuA���Z0��U��P��J��Ե�@P��砡>e��W�T���tZݫ����z��Q��I'�=�I.�ɋ�Ϝ�RNh�]��;�����P��g��l��������3��7¸M��l�#��eE��^H����!M���'s>��6,v��uߢDE����O a.
-��'sR�M�Ō�x�i[P��|�G�e�b�tC��4B�&~䪗r/�pR[�q���]�[?�bƕ<�$��+���5��:�Dy
��w-�֛K\t�������s��:�ˡ��w%j��?�!�s��G���ں/I�Z�`%��0�f5^L�LhG�f�f5�� �o�y����j�A��4h���x	Y� =F�2���q$��hK�>T;I (dsN�3C{M���%� $O7m�{��2������p�S�4C���J�	��Az�!�+��Ǯ>ZA��kBk�p`�@���La��T`�r�L�qC��@�rĔ=���QVd��׊����G+ �<Ǿ�۝��;������JLK�`X�j�= �h�(�d�{�@��s��#/O! 9ۡ����C�r�l�_<�����g�0z�&]�l�Ǆ� �%�7Y|+.�T!�TU����~����NL\6_<Zu|�R���r�r�_�퀷_֓�'�z�2׶�V�1��L�U.7\��������b[�tȅi����sL�;G�u,|ɢv�2{U�vOL�e�<���$_�}��U�%�C/@��� 5�2��ÇOⳅ�#b��^S%�
?L�o�h|��A�Y<4�,,XUU���m	���04�5��c�Ix��|�\׸*/Mw	�5ι~c�|o�� )��·��)F�&����o�+:fїO����w̢{$��ZR
B��[���+ܯ|�t��ظ�m⽃#��J�	�͒����و��j]b�	�"�5�N�G	nu�������v�<����D���]�����*6�]�70�|��W_a�w8_�����(���V]��ݩS����nvdI$�|���m/M�E�o��y���t���}����J��0��[6)�{`ĸ��0-��F7?>����c�ASQY����3z'�{�3V���#��^�8lk5�7gh���{AE�����V��8b�K'ݓ�����{]w����T>�#��L:�
¿�U����4gO�$V�8�\"dciJ#N華;��ӕ߹�T��;$�Tn�i��ԗ�l���9Κ�gۜ����|Y�1�C��h�^�S�4�dU�C����ۊ���%���m����@��7 ������X5�)^��#t�1�B{ř�D���g�V��3��l=Zc��'����ԕJm��N��m�U��u�=�tAo��g��_Eq�H�gX�����j��tu����8�ؓi�=2��%�;���t�z>e:5�n�L�Y����j��*�5�RL�3�ڟ����g���|={������%_�r��j�	�M�x&s��}pM�ʧ�֕Q�=��˳�\�x十͏�rW�',,����U
�̳AG�OU7ߟ�u�]��b��<2��E,��l'�lf���췌�n��F���ò�y%L�&�H�e�3�OT�i*)�������'�f��o�G��߅V��H	�O��t�sa�FfN�fZ6�ę���J�=G�q[ �s����)|)��]��K ��S�<�W�؝u@��N݅����m�%��ʱ�4c�^�[Zh[g; <_]6-�}�9ݤ��N���-����h�(w�7�y�zxU�~�'���o�yԴ�m��A���|^�<��Fџ��E�[�'T�W��U�-��W+,+��ˈ)�k�{�e�7�:î������6�Q[�$��{��@�J̆G{b��-ĵ���Ŀ�ߌx�t
�3�y�s3�g5�Ry��J��Pw�{=�p�th�WO*��H_�{����'����e�$��͏������M���h&zS��Kz����2���uU~{���`�N�ML.m�:|U�g?�A��������
l�/T�1�h*鵷�Րcfӑ����g'҂��N����5�����2w3��"�ThF�]�������T�;S��u�a�&����f=��V�,��)���rV���P}K{��~�`��E��#��9�O��:Έ;�Qe���l}wr|D募��=M��_W ���$�9���ad9��cs�#��8�����S0⯆\�\��ȋ�9]Ǟ�bj'�X�����w*�`w��Cd�Wu��PZ��畭����]�<j�n���)(0����_�'�̰T`{x���5S��v�L%�T�ۦ�</���̥mx���e�a���N�)���-lrm�$�^�H��T�-^�z%D���ǿ��w/��>V�{�t����L�w��BT�C�������/��SQ=!0P��d0_�~y��0u��p�M{E���5:Q��%:QCt���V��^�GQ�wV�{���,+���x���~�����{�k����ϵ�0��m5� ��D&Ja��=��Y�TT�Sx�Y��z�
~ω�9��t�!w��C�������,��������JJ�/��V*#�����-d����ǵ�ֶ*W��7�ҁ#�{��u��%2e^�q
�gW��'�5��Ƭ7�J����+������4��?�g��^Y� z����@M���3����6�`�)z5��9&����
��m�6��G�*�NO�󂤣E�M�K���;p:��Ԋ���[�e��q4�x����>ə\�Y��@��v��,�\H�<�e�!>���=���C=R�V�+��"�mzC���.�ّ�;ZS�V�o}�$m��pV��A8D� �9N'F�Oz�e
$��Hw�~�I1��'��v�H�J]V�|�C]����::J��q�V�����	4|��L�)��J��:M�0� ޟ%�=�nɚNJ��|�ְE��J�?>�*�LS1�M�.�y���(��E����C%�4;7�;B߭�&���:ۋ)�0Y�K��a��ގm�k���~�ݫ���?������a�����#qA�K¹,�[�\��� :�9���#��� ����M��̀�[͎��t�{��o�Î�R>Г����ҹ �R-���tK���R0�ߺ���w�YA9:Vs����5�Q�7mM�^&||zcTk6:�a��q�LO�4*�b��W�v�R�<]W=+̹K��M7('�!��Li��z��Y�2�`�T�t�/�t�̑�z��iV)��"����2;Y i�ÿG`�FI'PX��J�����=r�u4������&Ǯ�cBLL�
X�g�Y>L/=k��`:���'�'HN�����y%�ǫ�@�m_�8'm����e84m�Ͷ�/���V`m��I�<�]�l`W�+�e}��2p��Q9�N�=�����<0�w�Kϊ�����3\$	�R���/��)�BG��<^=`}�6? �Dz����+�ط���o����/P������3t;�XТ҇�W�[�k?��-�I'X����9��8s_�|��g��sݤ���t�a�]a���{����<�xF_p!�D���b� �5��?�ը3�����6>�H���?9��_�Vכ�ݧ�2/���qR~�?-5Ld�hh�=��k:�Q���#)m	��8�C�	��G![���h��(_\�Mk��ݧ��K��3X�?K:��~��,3+\�5�V�q�0P�J߈����d�ȴ�tO}�۩*����ܱ1����Y묐�D�j뷯]�!��8�*d<r8�>d��G��/���I�Lm �R/���w�Cע��7�.9�b��#�������:�X� ����������+_� )��9��A�)��l9�_�a;����*@iS���2����T`T����X���kR�q��Cic�e;��|� ��1_������)_��!4��è����)濽��9����:=7��s�1��a�y�	��9���n+�G�M���E�5��;��(����m�|��8�`i�5�Nk�*��4�
 _�M�	�>���[�a��t̍������ۉ��b|�0e��G"�\Z���a�R-���z�<+H0^@v�e0~�r|dT��q��˹�����aR�kࠤF������>�DpΔ� W��f'��"1�9$�q�ҲG�����3�����3d�SR���UQ���2��A�1dboS�X5���FbS���](�ȁ"�� +��.���ϳ�|���r��k�f��>�CF�+�ЭP"+����tq�Y�-_�*рY�5�?l,���)�h�c�U��ẏ�3��u�&��o=���B产��9�#'&�:l�M���u83�RQ�]V!���h=�4�վb��Y��V_�����^�=4Y/���j7�dK/�f8y�tB��D�#=�� � I��DC����u��O����������t4�j�(i�o��s�=��k��xJ�cj$�W�h�N/�xP6s@��z�q����^Ced�Zg�F�(U%�}``��2���a�[U��#F7�Z���=��ŚNb鞹;cQo��*8"�ޢ��V�(��t�ݙ�PN�VJ��d�y��%����Y�2����M���[��U���_=�����ѺCF�����u#H4C��������Rn���H��e�yGf���H`ml4�ƀ~a L�w��_�\w���D�K�/֤�֋�O��N��l����2��k�s�y?I.s�ek��?�ʾ�I"n��5��q"dn�u$h�z�i��o����w�rms���s]ANSD� ���a�������q��/[m�P����}����ZW?`z���WU���%X��~Ne�y�!I8�y�.�JƜbM��+��妌P��l�s��'*�[ُ��f��2��rM�uuS��׾	 r��s��
�)��PpA�|b���,�Q#]����M��\qC��g|?@?�����;g�l�W6�B�،�W����"}O�[��U���b�(CĜ�;_=�v��T���8�M�	B��2�ݰ�Y�_����K����8
-���m�_����.�奐��s8�G��E�1��z�υ�8#q�S١{c���ϗʝp�ҍ���p2o�I�f~�[�(�����`�%�e
)V3�<>(ǉa�l�	���SH�Xͱ�^��G������7�W�W"S����[!��#ް;p�H����L9�=�;����)!6M���3��suRL��^�r�&�F|!�@J|pEsx�؟�IB�h [�I^CBv��E{뷻z[��塅 �@Et�����w<:%6����'����"܌萸a�d%m��������Pc��B���P�n֨
���ʗ�f���Ǐ0tvf����N�Fϥ�俆�Z���Շn�p9�&���C�_��|�H?�A�]�Ob{٫5&,�����*.4P��s�0�*W!
qwG=�#Ry/������7�%K�����!��?�~U~�xp�#����*��齊uE\*&����Ё��C�ҭw�԰3J��g�����i(����bn�Zy#D?HӅ�|����D���om�.D��X&˚�mH��U�>X�=�+.Gw:��<K�8���)�w�U��W��5�J*���+'��8w	����S���6&��P�v������J�����S�Ĥy�eb��א"/�TV�.׾�9���Y~���E�}���ܖI�:۲4��<� n�8��MHպ�0]s���Q�Ϧ����v�|���E~������P(T~x���t�;�TBE�n�@�6o��Tv#6�ԥ�z�����QJ AH��.�C"�2�-��S\������\HR.��)�#���o�6�#{�`�e���c��=�����X3�@px�Pt@D�Ǎ�.�.b���soұ�*��@ݛ	�K�Ƹu�mA��������X��qt?Ӆ�Oށ@���/W�>�A�?�^�t� D�D���)=�Ó��T}kL$��ާQ&#�ZVs��Ѷ's��܉��Sw�MS֥g\-�?A�._��!ߑ���gP1��S��|�+�Ӗt l���M�$��/AA�ö�L�6�	1���Wm���U#x�ˀl�
�2;��@�C�S��)�.7����R��w��W��������@m?���&�o� z�F��B/j��k}:by�T, O�y�]W<�1��k��$j�s"F�'���sl=t�#a�޸����
����4�M�E�	�n=�`sQ\Z���tH�3n|g���[> DCP�l�
_QM����_�dB^��6��ɉ�z��aelv�"m�SCH��+M�N�K�np��T4��"�����O_����ASL����<H���#!�A��jTn��dP�!���4N����^��{M_�Lͫ�{����N7o�a�)��*z蛎	���`,>5x~��!�@�6���:�Z޾<v�I�[�
h7���,\*��N�yUۚkF�o��� �9�ٹL�u�o\���x���7�c�����P!�,�U���W�g�C}9�N�g��+׬L��FT/$𓈕L�@{��v7ӓ���v�[d�0�ǎ.�����:,bl��z
�X�0i9N�,�U�����@a��DX�@d��� p'c%~X�n[|�h#���Cl�{������A������jvZ��*��EW���԰</�[�3�=d������,Om�zA��j���E~Q?D�s|���dl:Ǧ�p�Na�k��P�������x!~@!\�����Q�}�����W�~?�!�����1 	z�R"=�3�$nZP�A�d�*�ѯ@��ۆT󭛖��h_�c,��o�(��|��r��r^Ώ7��0^�}���bO�1�B�b�	k4!0L�D#&����n���=��D�j�!='l�%�y�(F��2�=��U����5��{���N΋-ז:ˑ+�'��j�{#��(��0���	����E�g&���i���?p�gaT�DZ(�y������5��%��Q	v��z������x�������-P8�-r�pgU<o�h}�є-�r�,�VF�`n�R�^J:/�Ĵ��*q؈��m�٧�jj�bKΒ���O��I~!Eek�<J+R��*��|Z��/7��,�����"�('�tT�ʌ�����gA����OWq��=-}��\]�!�&�([���^G��
GM�/��־��3z��Zt��ȱ8q;�i�5T�����u=��A��O�O��]����ⱁ�e��������9�rL�����H��Ʀ��+1~I �n��CS�'Fg/Y~�s=�ػفZ�"����΅ḃP����X����&�8�_�K�ח[?&utej�Yގq ���W>-3K#P��dϦR��]���]�ժ5�J��a�a�����!#���!��q�S�F	fye���u��@F���-(J�0��+ܱ�\ԛO���XL��&������.@G,Y�u�[���94�<�C!\��h)�]p�s�	��u�4_��o�2�[��_�+�)1.�o�,S��5Z���D$c�=��}{�oȟ<���o1	���&�͍ն4�4���W$��x{a�v�[�OXڻa�"K�����[BCM�4(۠?�!����}M���/�/-�)�C?��� ���6���j`sh�G�-җJ�_�fo����z,'<�
��\�$�Hг�	'����mcx�bmtY�y��`�_���-qk�p���z/��O�"�!~�G8����.S���e�U�����Ĵ��L��ӿVC4�:uU%�+���#�^vf���]x�8#�ɥ4��m��?~⯘�ts���䯍aH|+���bV�98��
���?E5�����d4����_��ɜ�b�?�j
�e�B�;��,����:^�mL뚷��p�j-�C��6��B��`N�d��|������(.�H"PFmR|�ֶz�a{(D)_yG����{"C��k�mڛ<��l5�&�NKBΫ4���,c���WN4�����G#�\n�0�տ:�=�*mΥ�����?_���2�����ML��,�Q#1�jU��֐،�~�~z_�Սy����6�o�)�E��.�v<�h�zZ�����޸�YSn�>J+�}9���O��}}��w���ɀ?7�oS-rM}�#H��%JP6X;��&�:	=�δ*.I��`�i�d�2N�.bH;���c:[�1��k�v��`��⑲u9q��#h��V$%�o�i	�4�e#��m�;|\*`ٳ�e�e�a?Hc|Tý���%p=�/ ��Zp��'ް���΋�#c�=��8O)���{�	݅�ԗ�o�a�Jes%/fef����'�]�m���Ǯ���mY��s��6'!�a�$�I�oHd
�V2�O[K6��|���h����Sh�iş=Y'Ɩ�f�<�22�|�G-�����?Ά�f��%����!�*A��U�{V��ey~�vq�����GDG(�~Wo�9��F�����j� Y�?�v8�cK�L��7�L�6qoY�.�j��I���^�t
י�s���X�À��2�V=��B(`��v&|��r�1ϫ�n+�{]���
�r�b�u<U�>I̘��Ѧ�������l)�tD����ٗ��s��:`ߝ�JMaIPkcn������Oρ�E�R�dt0�c�S9��غ��9eA�P��c�҇�u��YB;NB��`�YOM�]�K�i����'�ϼ�^��I�b=B�������8�im��[��	�颂r����r{Ͻ��J�@��8ĸ������v�5�e58�۶Pa��t�G-R�x.R���*N��Ө�ǿM5�q�jѹ��,J���;WeGC,�gt��H�ǉ���Q�\�/�2p/�����[&�:?��(��ړ������n�%
���B��I+����K;�靺-��\Ƣ���y�v�s���Mr��������X7e����9*������rc��W����(����~�^�2��qqJ
4��o쓇v7�õ��E��j��D�2r����U���Ï_��I�?�B�jE e[��Y�+��#>6OZU�B	��
��a���d^�`�/�ۺ@���{}aL_����O�����_l��G�+���YO����λ�'u�dC�����)9i��i�u�7N��U�G���%p�?�~ׅ��Z����]I�(�y�PPC���)�%�mlm���u�ͣG���.�e1-����zd�\X�^��c����:��a뿞���@�+�p�x�����*w��Ԍ+l�e2�F4P2���@LJBAn0����T׎������N�=��h�R�h�_����s���QE;��S!��3�/��Ϫ��փJ{�s�|��Y=�:����^V˱ʦ-2��~�Ky��Q��Dlg���Uv%8`[��o�e=y�Wa~w�g4hɸ� �3��5�/�qT6a!��a��p����"z���W�OL��*"Y���w.J���^�Hv��%a��$d��ě��e �_'�!ߜzN"-}��T�{Y�D*Tx'H��\�3/&�)_���[��L�^\OtD:���.?����^�q�p�17���U�X�8arüOT�l���& �4��miR�����[�9C/��>�8��r0��ꇡӯTN���o5��C��ױ���T1.��*{l����6�ۤ�п�s�en�wK�m`t����d�o��Y�����ܟf���Os�j\ݫz@���~�7�w�BIE�Y�y?Ƕ��=�ION&�0EG���}�GG�M��e���;*A''`��ޭw���`����'л�D��2�0-�,���_ndO���f���;���4����嘆��gq ������P��9&�P��I7�̫ˤ�*�>\�|0cgV]����8`����^�4g�ٲ>���~������ER36�6�&G�d ofe�6���L�oR=m��L/��!B�N�K�۷��T�y��o�`�Bf��Ns���l���r;��,�$%w8��`��ڌR�����hl��������(O+�c�i#�F����������/<����V�{�_9r�K�70a�~�p���˧1mb��|�se�0jU?{�xo�Yc�7'�X�4	W�B�n��\\cDp�c^9IL��q���E��p`�!�����,�4W���*�`�w�Y��6["4��,ö�J]e�A�؟|� e�$�m�1�gۋ�r J;�s���9_�ߢ��_"W�@��wUp3o���Uk@Ė#�g+Rb�>+��-_����:a��_�Դ�!�* jmȚ��5I|!�ICT;0|���Dy�
�oV#���@7��q�b�5|4,t"9���Wv8��ĥgz�bY{�뽁����M bJ\�CV�����А�訤O������Ы�X�T�w���ȓNX����S��4���Br1ǒg6K.�N�O�����W��1�n��L���&BQ���RO�%=?��5
2[��g�ldh��b&}���f?v��{1��v�Zw��u�hs��bF27VO;ω4��X�G�]�KT���D�}.���/��0I����`'i:j��sC{�W�����c�%����+k+U�Ob&g4�Se���/��A�8�������QA�K��2�.	'�pjBrb拟�p�L�N��gp<��B���Zeyۄ�v��t���RO�Q}
F��+'Y�g�'��F���N��X��W�D68
�;J��9V�"?�?�"��Yw��p ��txh�4u��E���Ds�����K����V���(� ��XϏ��ݪ��Y\��f�bï���'
��ܷ���B⪣�$Y]�]���0jf�z�d.�%:c��Q���.�>T�-L����,}��� N���.�bn�7���]'���v��7���ީ'���Â �*����bR���}����#����R�UG�,��b�1��#��N� `-��}i�t�u<�ܲ�.��0$Q�����y6���C׿����g�ge�XC�	�4�c�E�����&_-��-�D���5W�F�1��w�;"�ۢ�𡎤Q\7����йd��_HSk�|�_��U7g�!�[d*.7m��&��;p�.P
��r?6a�/�A;��R��l�S�A��-�tD�p�U*f��C��wY`�>�fN�H̰Rll�~�o�'��3ko��O͛c�w;��"�������x�Ɔ�D ���1u�����տ�(C����'ۅZ58���Ż��k�u���-𡒻��bt@�����'2��B��FF��������R����x,f��_;��z'O���W�!�汎��K�:����7��(�}�&�ŭ����wsx`����iDP�[ 슺��/c��Z�e����y��a�D�>���z�o5se<�o֊�'����-�������Y�)�p������߮�8�Gg�pe$ݛ��^[�[�Mw���|���>_�޹��'��[�]M��/~��G���d�"M�4��5Or��OV(���=[�D�0_Y���m�~�`����*�T��1�lX�.0�prX(<�^�������Htu�=	�v�uRY��E�0
'�G�5��?O0}��[��jJ�5"&�P~�F:J�G.a�?l,�����jk�A�� Ir;�s&y�й�ɾ���_ù[��t9�:�w"=�}/��RăT®�"��_���g5»���-xᯁ�1�h��O]��EBy�<�X�
L;�{:�4Z�H�n{���E�F�GBM4LvA����y0ܩ���d�C�T�贐/�bYē���L�	nu�5�Mپ��%@�M%F.����׾tl��r��S�j�0��+��~8�$em�y!w͕��`*���%�&=�����A�B����؛��jU(����ׇ��T���]ӿ8�3��;�pz�ss��OP6�O[�2����tLz�J;�?7 ����io����[{�O@������m��wS��~}ie!�/O|�1���gu�� �,X��\\�IŒg�O9F4;�ǿ�d�@J���SPބ��W�zx1L�m�7��Ɛ4�;>�b�J�=s�̿���ҝ&��eP�q�o|R�K�*)a���nC�����wY�����T;N4gj�a%>�sLh�t�=5���)M5��|��B8��f���h,2e��k�O��+�l
��Y����Ox��fmŦ���x�W��'bS+��J)s�#~�`��}ԃN2"�Ǜ�ő�E�d&�kH�x)U�nL���Y����Or3���C�/�,��Z���T!`�~�P��R+P�oM�����¢Uw��E�3R��U�)~�<1���Ga/���9\��weQ&�~�����E�k;�X��Xn\�).��J>^��X	?�LXM�� t��iӘO�œ�����{Y (���n��CӘ���w	��RE��c���c���s�o\�D�4�m���w�!���&���Ӛ'�M�L��UU俻�@�����_�a�F�#��ӫמ�Ŷ�πՋ,�!��4t,e�q_@s�M�4 ��+)}/�	�u�9�!��̾���A(:JR_�;�۫���=0 ��"}SJ���Qc�6�BJIs��+��� �S�«�^{��B�=z=�uq��l��<ŠA}_0�%���Ì�;�)��z.I8yǌTlZL�,'��ȁ,�3G��ע¸vj��<�I�����v�y����sB%բ:1e�@�@Q���g�'�U6Dh	E�Ov�A��1�O-Ͻ�兺$��c#�.��c!M��'��K���ʸc�+&����zK�j�I	X�6@gR=<���_��h}����^��X��hw�"pN�i��:}����qhڀ++�;BP4���i^��*�}n=�O��1鲡K�Ew��GG�h��6@�f�i�:�]�s�^�\�RJ�4�²s�5�E�A�f].EWen�3�#������8]R�R�9��KT�:��PZ�`1�h����wO���B��-U�(��l�Y��6�֥u�S�	?��y��_��n��{e=j�4�fc,�Y<;-�8�,�[�'����d#2ׂ���=�/�e�v<�o��X��8���)��W6j�O��s:�P�lg2���%���b���מk��x�|��Q�A��Mz��m~R}-���)ب��{��揝/`�%�׈8�ܣ_�8����<L|��W?Kp����*#b���Mc�y䒆 -p�� 5��`��uoK��T��034dHZAs�p �
J)���'�����O.Ȟ��MV�%��9F#_��J�r��{Q��Q���w�^XZmh��֚�ߑ�\��������6.���	�c�1G/�����=[�e�p���Ad�Q���{E��R���h�й��3�&��j��d1�`U��'-���G��z� -��C�/[����5�m�{�r{���ϕ�Ir�\C`z,�x��,�$W|�;)z~C	W��v�{_�ycx�>�D�_)����=86����,�;�xFAp6{W��F���]q��ࢱGYid��A�,E"ˇ^,�-�)�w �7ɏ�k���$�B�'���Bs�#3��Y�_҉���:�f-yv�`�����$�Na�*�:g��r��pN��������Y֤����b�L�h�P}-�����y�c�aRe�?��Wo�[]����ZS�����0g=ʁ6G�PK�K F�=%v3�,��HKCŊ�O�y�|2Ԡ7� ��8��>K*^L�+Q�����ʵ��'}�J�|cQ18��<n��bښ�
�{8L��|���|[��މ��p�֙V#y�5���&ACҮ�!��_�ŋ�	W��yVd�4{�u�aD�Lh�T��:��96Q��Ю��'� Նl(�V7�%�n��-�Vz�#�zX5@A�������ӦV���p	�!J��d����	%2^v�}mlQ���Nl8(�(��� @�Nd���;W1��k���O͟/����u��t�B��s�g��1u$a-�����o��v�0�8ZZn�I�ȪL ��}��+Z��d�ϗ�5��H<�yc��yiY�����5{&�{ޭ^�nD�]6[���W�q"Q9v���ٿ&���G�_P���"�ڎ��E���h���}mk�b���TYQ�#V�[�ƀ��W�O���_x���v�BK"�-#�>@�x�W���;�%;�@B�1B?a��)���_�������s �9��ƌ���9�Y^�������K��z�4����h:���B�?�%͕�ȁ�,{63��H�D2VK�	���1�td>�ybAz��'����x99��N"vjP=T��?�H��[Z�Hg!g��L�Q61=�������b^��.�	<nk���XRZW2n�$E����LW�ӫl~H�crJ���WQ��x[���Tel�j��	���9S*�����*Zz	R��8�/�pl�����%%�W�֜���\�F锂Q�q���2�d�k�4v+)h�����y� m���Nk�����&) NE�ӎ�����S�X�x��BȻ?�]Ε?7;q�3�<�gIm-� F&-�(��ݫǽ��$�@�?X��,���s�$�kt��j������d��_FD�R>_*絊����Z�޾-���2U�h�dN�Ҁ?z%��K����ٵͪ��Rj v�l�9�ߵ5;���p�1�����o�`K>5����g-�H�ITrLQa�9�I������o_�wϗ�<�mX�	zx<uIO�XÝ�����I&����1Ԙ�k�G�%
x�t�V�R�z�x�����N�~2�� �g�߮ʻY�Z��CǾ��j}�����6j/�ʊƭv&`�it��q蝜BT�s�<?�w�x�b�{��7�> ���}�Mw�6����0r�W��h���g�[5>%�*Z�EKd�kF��7P~��5.J|:�F�x��$����>�|�]Aw�w:�d���Ŀ�����F��<S��sL��W��n<�f�(��/ߋ�g�pP)v���i^�Y.K ���i��g�!u�UD;��/�ұ� �g�
$=�㇈[a��B��VX���S�x�y����m{�H+t<d��~� `�G)j����d�U�@������wp�F5n��pW����s���o������h|j�:�of��$��t|�<~���Az�5�k�vcWU�q_Ѡ��l^8��kg#�n3�5�к���2s�_�����r;7�!֨�uPO���'RQ=�����������i�m��$���ڍ����v���=�����u����M���#���v�agd����45P]FCp��3?�\�&?�p�-�+o����r��s��7�{��pPn���Zc���g�V.��/ǜ�#3��(�N���}h\��[����3>��x'���f����LHX��k�:2<p���%c�c�TO8����|	�ahA1�V�� ؼK]���v1�ی�X���~}���k�x|+�E)(��G}N�H��75�T�n:d�눕�h �n�D�G�V�gmc��!4�v3�>�l���"�>nB��v:I��$����>����Bi\���.������]1k�F�V���ѺT�zB��tY�P�>b�������:9����}*b ��;iY�9�1wwm��QrƮi�c�5?�Vl/��I�0��E�[#���-=^������_y��x���
 +M�J�-	�
���'X�e���3�?/�z��`�
G޿Tg4��=��үO	��db
�Ek�K�C���8�������黭����n*����Ĺ?ƿ�6TF.?�P�4}{�K��yhJ�{,o�E%���r;�wO�Y�hl�v�$r^	ډ��Ɉ�y �.�
�#��2��̚�\��҈��'��7��vV���0��ڤ�����* K¹b�+�w��7�][q\'g�)�A��ޫ�)��T$�=b� �۔.��q4QU�3�0X�p�E�P<s����&圹`����� Du�Lv�M5�)�V���=n�q:>i�gW��ՅU(���Bf���~̭i��%)Q��;�@)�B���|��k���O�Fɻ`�I��V�S�Fo�������y�G��!��L�C�5���o����G~�r?,8��K!tTG�G�8���Z��(��̖=�|x�lG��y�#�R]Bv�G��WFb/a!�yQ?�V*�����n��95�A �GS��j��w�3��r�viü���߈^��g��#$τ�Z�י$�٭� G[-��:a�r��3�����&�W�@���Γ?����qS���k�>�������֣th�����D=�%�ɢ@p���֥L�У��R_��q����E&�o@n��BOԏ����'�?"I�`&쇪�_������\�v1�H[Ӵ�8	ƜGPWh�K��`+P�\
g���Vx���~"�lܦ-P��ݺv���LB��@��~�$*���)F��	=��#�rb-�1Ѧ�
?Ͳ�^k�����u�7��XG="	�;z�DЛ�
pq�h�f����V����_�}��ߊ;Gǭ/8J%�!8�-^��A*��~�Z٧+��|Գ��gԒQ�ł6I2�Ж�$ž��4Nd�����I��������sܔP�k����<_1�`(�U�7���@8�Xߛ���V��8���e������o���Ï�oi���_D�i?1*t�KYk�W�v?���� ��>���,�ԣ�B�uݪ��s�2�o����S�,������6ŷ�e����*�97�D���g���֪��i��xT�T���c;�!ז�_	�MB�@�	�_Й�$����Q}��JH�ۖІ2ⓥ��K�c�;m�)csO�Y�u���;�2��>��2��N?�B��ZeQ�<ǭ�r K��U|����6��v����Ye��ſ�p ��9C;�R�k�����n��EI�]h�b�pb����?�16�����l�����P�ۛ^p ~"�HU��z�r��K�w����l<�ol��6Uy�X�SSj��)5t1/��I��.�N�S�.���3���/㼩�?�~���L�l<!_k�x�F���k�ppI�9iQ,�)N�v��˾�٪$7��9�);������NHJbs��cp;?��g~,)����F�j�mG�<\�2fv����+�*�v��c� ������'�n�j���l|�d�T�G3�ҧ#}VI�$��&�K�l׋F i(n��\lh�  0�\L�JQ\KD���w�U�>�yNNN�O��k��`�~�����Х��Vƕ2��6t�Q�N�~�l���gCw|$	�NO�:�'i	8�u��A^��Gѽ���DL�.�w$ *�4sw1>/�r�-�L��G��>:���:o��~���@-h�뚸^[92�a蟭E���m�C����U�`�fHj�7t�Pd�)��@�<Yw�Q7��	 �'B�>�Qv�9�ʷQ�7�<д{�U�z��/(2��ʼ��?0$?E�7�Vcm��|V���ۃ�"j���0��	a�\ E�|��1IK�r���d����h���j�m� �f ;OY��Sf@Q��vj�H߷��a ��(f�Z�g]��}+&���N��%!Z��t��`-���2N��t��#�f��_=�fq�̣��zrώs����|M�n �L46ن�L�t����T���Ye�&����ʀ`i����{�!e<D�&�^6�.�]�"���� z`蹅eÂ�r�z��ѵ�E���A߆k�j����kp���X����c������d���2��{��0���@'�q�M���/g�L�2>P�g���<zK�%��춋��($
��Cf^�X��<ۣ���u��G��cZ�MZ�[Ϗ�z��h ~^�z;1�Y���F���{U���x��*̯_T����|j�_0�D5��;b�>'�h�,s��������p���w�����+�i�[7!����|廛!�]�j�ޒ�s�����ͷ���̟4P�^}(�ܴT�7ݬ��!A�I��,����N) �k���%f�A�G9^�zT�ҁy~������u����:���>�k�1�0֠���1���yv�JTC���IeDS��xVo�f-Z����BX�����2�����'iF���s��|ѧ5?r.�2~�/Ap�1�~��=H'�u`�ze&���U�r��C},�����IV6�y�M��f)���w�fDY���2���EF�����wE�v�Q��Ժ��k�����9����*G؉�b$G+U�yρY �(;�D��D8� ��G��O֎�����X>����k��7Z�kFj�hcӅ����S�>,R�d������2��m߷�ye�ks�zk�;��c���E��T,Fx�.�?.��9�:�=������ad����u���9C@[�B�g�ސ���*�������J���@��9���5X+���.D�v���)��g^����e��������W©�'����O[38�5�hK��ZCr�1�����3�40�B$�6�a������#�% �\��\��eM�yk��a�ge�w
8u\A1ډ>�sV.��V�g�)���=.�9��.�/'�B��)� )(�J��\�/9ߵ���*�7�B��!��w���ĝ���J~���0 �l�5�Rc��F�@�M���V9/�a�ٲ��U�)�����=�~^��Ë��X��aC|�����N'g�� ��ؗHmuWݞuYd���ϞFy���^�$���{�vݯϖ��#���zP������������@���F&���))Ο�u��+��]��!G�cwE��
/9k*$�[k+�E�j�u57��_�s�Q� �(��ׄʓ������p��������o�/coF��JJ
�E�
�S�>��оߝnr/�>!!�L�1����t�>�\A��@֚� i�L�3�b������Vq15�P�}��,oF}|�fǔ4Qw��#��k����bnZ[���L}4Ҍ*�a�B~���V���Do�\��OqeƔ��Ӽ����|��ײZ|}��J�Ƨ�(����7���s���7�ᘭU6��i�!�v48���׻�O���uh�´�A��3�64�F��A��C�	���N��o|�����^�k����9�Z��x1�OQ�[�.�Xk(A����,e��]֌F'�[�ÝbS/�#�?��*��}D�"eЈ��H�tyQ@�;�E:�NE��.�J��E������ ����׺��������}���=�#DX~L6�Ng�eY�K���B�j ϯ�6����I/�\2~�|�cp�j�/�ܝ����-z�vIm&#�{7��sWR��82��IFq�,���\�ZJ��Ӷn� u�q�w!����!�)îO�M���JJ�8Bx��H�aC\�Q5��%U�$�Ga���<�[XIg��J!t���y�<�pzvT[,�^���4�T���z��j�$���d����!H���R�9��N,t5�o�c���3�����KɳMd16��P�p����>7�����lӛ�N�<�28���H���N'��_�Q-�?2��u�f�y�x�9�\�iB��У-//հ���|����/Oy�t�4ڗ��Bfre������0�l��}$�\2-gh|�%��荆	�0-���j'}~{�b|{.?�a�	_q�ϢH��1:k��t��̎��^��]"x�[Y�S��E���D��U�Cl�wm��u�U#.5�_H�ܽ�oU��i�)yI���(W��lƦU��Ky��0�.n��$�D��c��ݑ�5��D��9���)JVI�6�Y/g��Q;�g�l���-����W���խjww}������-��$x�϶a!�ې�>h���ߊF�a��TdM����}�Օ6n�>4졸����ȼ��9�8�j����^��7�S03���]��U���ͮU$���`c�<`�?~z��r㻘��6��XW�{i��V�|O�Ӓ�'ۿh� �*�[�L��=.�D��@�w�R�#��VJ����������ӿS�]�N1��E+&�f��͂��N�i�ٖ��m�8��%��E�Ců������_����؛-�v���YB�vZ}q���/rQ��>����q�@ާG��c
�S*ٛ����%�g�I����kn����Ţ4�$*�_��J����G�[6�F_�d���WٷwQ�W::Of��p�9��.���/s���gou�WEh�--����d�C��j������6p3$	�C1T	�u~)�k��\i�˳&�g���t�b�h	/)N��1pu�@r���F���0y���BC�����?��,�/U��ZZ��(KW��b�O�g�6I�:CƷ���{��1�aʑ+Z���]4���>D.�_����gD�谏�/�l0�'�x����G�A�#�xg7�{
�O�[Y{���M��[����#P"$ـ������a���o�uT5��vS���,68U��6��m��Ƞ{0�Yrj43 �]��,�^��rA��p#�k�;�����Kg�	¬pD\W�Gw@Ȯ��+Yk����0��.G�"�s���~���=�?�`�	R��k�
#�:DEv�(��G�~��/ə�ND��.��(4�ӓ[��U�m،��P@����j=<��ks��R��h@�VO����i�HDE�T-��;v����r��c�J�U�/�9��	+i=+ M���bYsv���k�zT�!�뙈vz�6��5ѭ��v��]_[4���W�jz�t!�G��T��k� Lۑ
��I���d ����zK@���g�LD4��n��
�6}�3��}�['"��v5j��Ug��_B�ڹ���D1�3u{.͓�^j+T-�/]�RV�Zd�웟�V�����c�L�c_�6s��ׯ�"۸�Hz��uU@����K�]������j�.�P]�'�V��N7�ga�<�O��ӒK�X�/3lg��5�±���*�cd��BVul�5�d�l
=�K�f�mzyr���L�
���ZZ��h�Rj.��nl8���҅g�+��.�ޝ����u[��.�gu�g�x�S�6]���ߩl���� �n�l�o�~="T���ùR�'��?�rú݄�Δ�o��!pm�'�����,���� 8�q�l���Qa���յ[�nȱރ�X��t)S�-�nbk7yKF�*�s=P��Q��z��4�h�����`��|����pd��(ӲD'��߯�m����D�x�����@����&>����P<��,�1F���3}�����Л"����#X�������'���JG�j̜я�K>^� \-\�=,������b��.8���3'�mt��8�{�ޘ.-'���uWƍJ�ˆĥV��md��@"k���h�u1��K��Ef������V��v�p�f|lRn x��5<�QW*��K'�@�@�ՙ���j��	1F:%�C9����wPt��{���R�,yW� ���͝w`d�<)w�LÊ���k�9�օ���ԩ�U����U�z(A�q4:X��1u?7	$����	r$�0�^��!��t�S'�)}���e�WZt�����O�5�CO.ѧD^U�KJ˯a���j���8c���cQ��u=��p@���J��w��S禊a����n��w�5�bu�]N6��ҁvs�Z�f�yt��`��X��:����vU���+6�|6CE�O�կ�v�y�Աn�5�g��S״L=h�Y�%5��c5�g�+0�߈�"f]vFz��V���̝:�4��6�^*���	��&�}Z��8o�����v!�f���S����^�'��؋�(��uB�����,݌WF�"�J� %L���Iv�h�v���Q���08�h�T��%^N������VW���"���9�2X�s|����f~:��+��e��/.(���Lɛ�Q��`N�x%�v,_�7qf~�����Cl��'���2l����I��)�+���ԩ"�D>$�h�i؝�]ĭ���t&M}²o�*v�Q^��\����׀����j
�>-PCp�<��������q������H�O:��l��x�X0]��y��a���m��=XH[��<�jtqW-]&EF���g��ATp�,/�݀n���3-Z���;��n4kZ�TP.�(��]����?��A��4k���Fk�o�<�"�3HC1�F� �a鄙��Q�(��[���}��,�5�	����Q����4��g��ͤ[yӑ�@�k;]�.��-�t?7��J��Zf�N>�jF)ƴ��}���~��<����Q���֬	"'��mѝ彩����²�P%�ən�G�,h��K����@"3���Mlq��i|,�/l�anj��@����E���VY�uW��:�J�̡4�S�S?�P���%��l[�g�k������ڴn�z%����/��N���o<��ɪ�[
��J�+ 8� ���-�Bm���QKwoծ��du����$���F������%�� `\�]�XkN	�ߩ$ ���G��}%޹�
凷S�}�Y����O?:ڵ�9V���N���X�>Md���f��2����s��hx�����E;���=�Oċ��^�^�g_���w-���H�g������uy�a"�K�t���BF2���Ҟs"S�p3^�\�ǁ��6$&'V2}�5��\�I&�+�YȊ\�E�]�:�d"���%m���>W��t�@�R�j�>Y^Ȏ��Jli�fw��K��=jS��K���;�Ư:쌑x���#^G_�8�Dt��3��#G�@D��>	�%1*�+�U?B_,�^.R�NvxгH����?%�r�{�I����3o=e�l�48ݵ����ۢ7��oĬ���aO��N%*���(z�R���Dm<d�4M)z��ۧ^�K�)7W�J��>f��c���kX���o�lRx߸/JV��g��Y���Z}�E��=a��-��:)�V
ɾ؏�j8��朒�l.���5����d�> �f�/]�o����q���&�|k�!�W�<�����ʷb�l8�P��u��W����
��1n|�J�韨���S�݆�`ś���>��u�}6�թ�xN��`��q6����w�|Z�%/��C�mۓ�W�?v�U=��鉜r�A~�Ø
��Z�bU@��ji���}I�`��6�q�/�0if�MlX�]��??���Q�6��<�h"��k�W�5\�b�o���-M�6��A[��׾�w�����*�Te���D����2+_NKw��VVzIQ�;-���
��9T�&aSi��K�rZlM��c ��XN���XF��e�Y����Rbb�����O����f�U]�)�)��:�'���T39ߑ+-O�v]��IB��2��u�h��.!����G�&�����q
լ#Ў��i��j�u��"�Զ��o�1qI��S�s]vX��4�g}�����q��K	���S�t�5�����������"U�L��ri��/�<�raq�{Y5f�d&�i� F���OL��Z5�-��
�7��VZ��нJ�V͇�	%*Zwqn���H'������	O�:g/7�d ��N�ݲ�����6{~���̫���8c�"Y\^O���]8������F_���g����E����^n��2nT̔��������j�I-+1K^�1���홿\O���RO���W��^��y��I��?$�3<���KΙY�n�ꗧl#B�XM�pKhUG��^�t�Q�����h�t���˕���n��as�-��#�`���i�C�ua`(�p
���C(�Ȱ�5�%n\x+  ��O�#gj\�Ej���K�Ԓ+	��M堥�~�`��e}�V��U�j�����䰿�y���OjT+���Eڱ3*p�/�tdӉc��$r)(��6 ގ@�4T_}ڽ�'��jў&��7�D��?ۦ]�j�m��%իh�-V%�������}�¿|D:ǟrgNƦ���z;��3��E"Ζ�q�/����0:К���TN�6�3���������>�u���!�{��F�L��n���`�� ����U����v-�5r� l46r�ؘK;z�b]4�*!�r``�(�1գ�i܄_n�U��U�i�}�0�4��/���r��I���ԗ���G|�h{�+=�M�b���E�*�Q4�y�{Ұvݪ���f�	���0ϵs0Zya���tu�q���&��qIC���T�($.������H��3N�_킊�*�v�g����Gu��\3�����Wx���J`���Τ��Q�֗+B���.wY��6���0�v�Y��S{�� (M%��n��Y��+���`�E=�$��e��Eö���Y��e����q�5�YUo��?��Y�l��8\�+�C��x�:2�}א���(�Z�?~Z�}ja�Y>��ϏJ��y�f�����5N�n��^��@$�_�	���:�T3P�(ċ𺫰}O��wk�����ᩩ��t��`Qgcfу@f��rm�bn}T�/�4%8��o��7�5�t-۹_}�JD��������O�M����v����]��u�V����w�(f=|9�|Fn��s�(��$�T���!�g}��+Q�^"�xܷo���k�m�%\�T�M��� ��8I��W�&��}U>E����+Fw�,�����5��';�@:�:q�m����Ł	��/�.�讕�Y4�(f-�1q��ƫ�}.�n��v�J���+�S��t��~$�!����Ŕ7-�qAF\��i����;vk]�8�879�V�/��.��q���zx�j�f���q�y�j�ԣ�t�G��3K����M�t��n�'P=Bf�A�[�}�Xm��(d���O�R�����S��P�	{H��(��x�����C�=1ګY�G$��fW��ɧ���!�$��w��FڅQ%��o�x��\���e�vp�>�r��s>TS�B���Q�3��I5�^7,TRL�|{u��m0�1�l{y��Z�y��?��dĬU���Ԯ>/u:�ɒ̔��^�j� �ퟌl��p1�^
x�ޝ����i�8.�=О���O���{5������0�ʼ��KALOEBOMq�""���*�b�,ed�m����G|o����j)slW�Nh���L��Oy������\���~��w��r��~M2SsU��;j���^K;�XZ������u�"����ޚ=�e��U��}�8�.���+;J���X�� \�^����[��kF���b���KB�k��q0�6�P}۵Y5�5��l�6��▱t-�eG��5�l���ژ}�\����}LҬ��V�E9&��m?)>}�(��Uƣ�;��b�'���gW�:�qՓn��/��!l\ܣ�3
�Y�����[���+x�Ys��;q�\g�Q��"��}��)Ib�Iqa��&Ȁ;�����H?��{C�Ϟ���Τ[�j��6-w�����V(����u>��� pE��ܞ���\ }���68s�p��8!��m1f�m��:[d�0�p��}ei��=m֩5�4?���v`6<:��j�^ߙ��	q���6�g��!a�@�p	{�O�Q|8�#*���	�U�����z�6h$�1�z��mC���������E��>�7����9�����G�Al���?m��G`��S���Ye௵Ƒ�Ы�m>�:�31Ia2�߳��w.?���ڥ�r��k�qqU_����{B|���(����j�8�K��1u�~o��o�W��3�w�	}f \iL��l� P�y���x7t�(�X�s�J�=j3��
�S�-ksg޷�4�A��p��-�0�ʎ*O( ���K�R��Y۝��j�F���3�dk&�Zt��t�ӣ������j%J0e�v��w���������U��s@��Y�z�6*@��=�z �ѳx� '$����z�k9-����M�TcA��52��h�"1�9y��6X�jQ��SG�"�E�!�_@��^C��u�_D+$bjͥv��^��M��i�1-�i���5
Yq�#�(�V�䁈�P��l���\�gVc�u��S9�%3hMf��
;d�d�UG�SM��x��<��1��Y)�eĬ0���G����S�5��[Ѓ�i��l���h��3���Q:�]�Q
>r��&shn�b���	Ki�"s�]�rx������[�0&�qxG���_���5�z8`�w�3`cU��g�ɫ���[�	2�X:k�.(c��s�ܔ��-�p��h��* ��+ҡaV�Xº��Q|�ފ���fr�eN1Fw%#~o�[����_��R�[�5�㆝�>�@�(pcd�G�(�3t�H�m���#@�u\����=���D�|D���dݪ�"#fl�b!��]_U���a!�Ƣ1Y^��a�)!��c+��:��p�c{mKne$\�B쳸��5���-b��mxJ
6��l县�*�A���|-R���Cycږ	�n�G9fC�s i}���#�$z��}�ad��c;R��QCr3.fq]�6tm�U;>��rt;�;�"�G@�?�,п���@�w!���c�X,e?���򉨛T�f�jN��T>�����V����?Ct�*.ʬ+k�����aU 8<Aِ?���İ�W�]�wl��5�����5� `��*̲�a#�s��<4o�x�s�d�Ѐ�엎�����M�}�`L��9Q�~ܕ��ePA7��*R��g��& �.�!G���?����]=������S˂7a�A��!�?�!�� "2:�De���C����J��P������{9~��ʣ�<ގ�@'�?Z3�Ya���X�ݶ���ڟքH��(m�&S���9���l�fLH,],��P�?����n�$WJ�ʑC��O��ח��;�<�A~~t@�Г��q�w�?N�
*�T���]��M�P�3Ф��E�E�_0�[���؁�=�������Æ��J6���)�%8Rt��:ݫȑ���|=���R��߽��x��ޟ�ͳQ]>���#�|�CnZ���H�c���aoy�6'�L���t<���!�F���T��.�aň�}�m3��v�t����}菺��ށK�Vo������hZj�\������|��a����� ��D�4iaE�v�f�ĘD�����+�!�Y��: �V(�kb�4�����XA�b��_��L�K'ܐZ�wF�����H�ʿ�*�r�4�hl��M�_yÿ���v�g��SZ���e%;MNe !��A�x�q�:�4���׌\���[e�&�@��I�4�VC�lK��a=3�.�7�E�N&.�E**|ˑ��`[���o��T�\��s���;o�Z-0�(���&s�\�H�ge$�+�f��@@�$&��g��U5�f�A��e�1���;1�6ĿO�� �ޡ�+����ˋ�XX�Yl���u��:�E"q���0�R�-����m�b�ӫ��}l�!�����g�ܚj*T��HUz�N ���~������Փ�ak5:x���y�I�ߠ@i�Af�.6r>}�w��l,���'�h��}c8��K��ܵ����i���]�oq�3+/Md�$��}�[||��,��.���u�S}�b�Ȫ���g� Z>����m�;������z���n)�w��V�]��t^Wut�O9Qs����N��s����C`�=����CD�����Y�#��Fk�Q>#8���������N&���S�J�/<��fr�g�?��l'�c������m�$���_�sٳ|����8����f4�ʼ���V��G����W����5���;B��{2�L�t���������e��\*�2Z� ֔M�"�)Y�?����$jv�F6����3�Z�p5'��}V�'��*�(dd��� �+y�JG��E�:���;DR[�%�@��n@��kc�����r����A.��1XZ�d;��f��O�^6��xM<��D����xlG�e5h��R�E����*�A�h�'}צ�`z�-�%��H�m�*��u�(W�v�ddzC%�wq�9*���V"�̭N�c�}��*�gxU�.<z.��^>g��	J(5Ѽ�ǉ��H�YNY�Y�XT��h���D���"�k�+��8� ����F="�ڋ�1t|q�Y����a,�5㸟E+�u>�3r=A;���"���l����|	Ød�ёƫ'�_����d5�F��g�<J��+ϗ�`r�?؟ECB#�u]k�d�,lbpt�k�އl��첄�ʘ���p�Lz�[�~ؼ�p�?�w'GLϊ�]��e�b��+�\1K"�^�:B&���{�>� �PRS�2�0��**����<v&YG{Sŭ,��cr�P.5�qW�E�c2(z P����NuGܗE��@<�3�4K�߱��1������߹)Y_���[�c��V��RY��̞9[�Y��H��m��X�¾���=�mV�gs:��cԛ��5�����'�iÔ����(WNz�����]!�s����6�{r��ߙ����d �,#������
7��#��;*u�z�GC��HE�U5�8+�awf�`�y��i*��nT��ǡ�~��O�����E��>��V �'��6�L���Å����W��0����xZE(#jd��lf�פ���M{�����P��>n�#-��X+V���Y����1�����(|����?��o����L�'ƨ�b���"��II}6y���EM	��&�k��_	7���"� �l7{P4gA��xw{{5?���&�]�^�#��nG���G�͠q����3*puxݳj�H�<�7���O��12Z4� ���i�Kzt�6�
_6N�h�z���9t#Ȫ*�� �
f�Pڭ
�PZ;�E��
)��l�!|B}@U�F]�w��J;��c������{��aBj��$�(�2�V]����{�FW�l�G����ʧ	��a+߳?h����+��g_��<�����7���GO��.��f �H�þ:]d��1��x�gc��5�R�Y�^�v4L��O�,�l�д8隗3�E|_'m\���[�7n�}Y�u"�J<;60�B9y��jß��v�A}L`�Й�E+��_ڶ �]g�H�����Na���������s�WR%1�A͎�h#��x ��V.Z"^"�X��v�*�a��P��S��S�9�> i�۔����>"U>����ᓣ���=_EW��Q����פ��,�sC@�O=�]������:�X%�f@�V�7���.<���'PU���)uIJ���ŭ)V���g�`V���	�d[��ˎ��"��O���&�r�6.��E�dP �s��h��ֲ�:������h`&�Aѯp�yd|&C9T�w�M ]~�c97\����g�n58�������)�z��w���B�қ*<?�yn�&
�]�wQ�#�ƴ�i&��u��^�ezѵ�5?�V��u3ࣶ����޶O�.�a��g-꼅����:Ì�߻�Ρ�ye$9�ށ�> ;j���`S�4��s�w74ˈ��"+7�(�ny1z)�	7�h�d���S�7f��|��z�k��l4���? 2:�?�&��4N���ox^�N?�ͤ�q�8cd,+fD\��;'vA+y�Ť��/N�{k�p:@G�ס- ��t�U+����]�y����x8��Ø.����`�|]�J�Y�~gNR@iW�J�Sv]GeĈܙAܨ0{��i���f��y|Є�@�ޑĤ��T�1e�E�6�U�T���H?~�ȴ�r@P�(��>*0����o��y��〼��m�r���A|���@�eu��kY��`4_����D>�aJ0�}wc�!�����q�I*@�Zz�mꏠ�`��4������$����N�rS�H��޺n�o�O�ܿ�.f����,�������@�l�K�5y��}��~�* WЄ2�~�~6��I� �������Z
P2G��(Q��7>���J�PA�����OGn�*�������Xej�������Mp[�>h�[�L�E�-�_���f[�S�
��E���?��)�7{B�6��0U�n ��;X�2�5N�<�M馓W7$��  �NC���B)��b����k����7]1���X0�߉%�`���ߓ����D��1`�r
�4�:W��?�w����G\��{o�~ ���F%Y?��H�<{�ccW@�� �W���8,:����$/�p5p����le̦zx_g��{x3����CV`� Z�πx'����f@�BZ���_�c�B���݉4f�[����@�����,��O�>"�����?P r��{����/���-�w�<���9���AAq�	�Y�[���sO8��M�!W�~� ���c|t���xFm��LɊ�2����{n(�Pޣ�<�Q�H2
�H��}���y����jϞ|��u��s��WD�{�*�C�Y�D�B����X�<���tS]���ׯ���s��M�����O��y������Gm�l-�Q1H�e�_���K�TB��E\��D*%�Z�l}�w�"���8���ȯ�Ro opt�y�箣?�{{T���E��,�r��-T|��Ro��1�is�V�yK59���n�n���B�r�Y��? ��.i1Hj�'�]��g�f/p)�PT^|���:��wlF�Km�w��w�$�b��P�9�ȕը�AXo婎E���C�@G����=�D���T���w��/!�T,����ӕ2a�L�w�����I�;i�P)Uݽ�{��(�|��̷yRP���"~�с�`��2�%/����Z�XVD³[|;�� Es+���)? �Z/C��q�'oo��X-�a�4 �n��I��`�	����BXP>#؈�9rZ�R+���w-I��D�^p!]���#��J ' '�ga7��܈��'<Ac���|�͑�UF��-��w�b��4��.v,�Z.�X���0z�g +n��g�3~;G�I�v�^!��F�2�$�.f��0�*I����"f:�:xU�'T�8@3J ڤT!���J�P�v=P���������	u��p�\F������i�:�A>�ug=a��]z�V��?7���Ř���BxR��g�YInA��I��a��)rL����s�]�Vh�$�t% nD�w#�;(��a�������t�$%��T|�խ��Wjl-�G��g�PM�_��ڥ���-����NoJ3r�j���S�冦ş�\#e��:�Z�ny�so�J_*�Z�,���t
����ߪ��T�Ya%E����T;u�s�B��׷�qq�����
�]Pu��߼�?��?��9�0,8��M�r�쩕�g��߄I�x��9 ?u+�w�S�G@E�,S� ��|JG�	�#�i��f�3-odY=��c�R�0������zӷ/��-é��щ�����G�<]�1�SC�P
U�;\lv����V�
Hb�O���<С��P=�5Q��P��@�bi�xW=���<�U������*�:��~���VZ�gb��F���Z�Ã�V�AFIO��iD_�a^y��$��Ն(/;���H�ar��ۢ�󳝡�-Q������{��Q�1@	q7�1�[O�\TN���%��n����W���I�i��j���G��Z�;�������\� Ϧ�THd��W��WD�Wr����W�p�����ԱaG��+� �vP��e�z����tK�]��Oh!w��s<t�Y�z� $��R��1`K�[�-!<N�"���׮s��r��N����@���*�Z�Ƹ���;�Jr��R�Y��".����{�] G�)�Y�&�3�ݣ��\���y�I���l�j;X�K�_`АǏZ7��S���%ɪ@|ו&Y}����T-�>�*����#��t��jԄ�2(��<h�pj�j~ew�<�X��N�Ը{��A�?���N������rzs�\��]�.ݽŮ��� ��ĎY�@ދ���=d�dV�DB�w"E�x�;��b�m�>��Ȕ�wk�����\<\V������e�8��+9ۀ�]1 �>`.5Bvc�yz��t��(����� �/�oB=׬��K�z�DH���!-��d e����H�q��KK�^nw�8(8�D jM��MU����UKݴZf���}GCY��oDmq�F�+諚�">��$E5@猞�̇:���V T&�s&1 ��2��Ͻr �;�wd�o�<��x��{�t�[ؙw���)�Cc�?jƣG�q����q����1�K"(1ea��?g��\�Q����e�3��_�e{]��''�j;�޺�r�3��^a�o�$׋��A�L'�������@��j��M�	�&f=�g��A�2��c�21��<f�,�݊G��_�R��evå���5��<`�� �b��]�u��[�E��$�Ý��48j�ӌˇ	ر��x�&a��2��?fղQ��� d.M��tE���*��#��>ޅ�Z�\�3p��cVՀ�o�� �	���X�Do����i�W�,+&̮toڹ�f���hC��8�dBT�D���UbP���t;Hέ%́l)"V;���NTH#�`qHgݼXT�P�9b�L��Ru�3�&�-X�*���R��|W y�fG6��A����vD�.��wa�#"o���P��`�G�Eq���\7^q(�2�l:�m�"H��S�[��g��u�;�񅽉�� �,���t��D�E����tMrk����q��F J�_��p�8Q���L�@��L�(�k=�X�4ÐA�aҡ�#����{��"[8aQ*�?��^�k�p�r
?��ަ�71T����O�o{�+AJL�hMUz��zh��`Hx���XT�;W�.JH	�2���>RR�Y6)2����b�8�
X6��(k]V:�˴١������J����˰�����E�FI#�nmӰ{��93�1��M�"��K��:v1��Y�j4R
U3�X���jى:�gN?�뾞s��Obe�SH�M`3���k��JR\�_`����d_o����GF�a #OV�K	�'�	������_7`�. ��E��@^z����:��c]rx�K��,����P
��?J]��a2Gw= ��kY�{B\/L9'����Ï�OaNx�Ն��Ʉ׻�Wl[�@�d���H���IS��k��ٕ��/B_Q½�J:�N�a(����+��fR�\��Q��� ����Շ.�@�����)�i�Y)`�'U6Z��OX�	�J�*Oj:�a���ɧ �<��.|	�1���>rPT��
�#4s7C2�H���7����b��%�V��ّ��}�z �����J }��L)dC��9m�br>
FF�N���[����?��L<�%��t�O?���@�{`i���� ����Z��2ɾF�w8�ֿzv�-dpWJe���!���^���q�q��c�Z�6�ڀ�%�JΎ�LA����dRO��Iry���&�ѭ���Q���r���ddAd�畡����0W��4�y��k:�Ķ�Y��r"�n*��C䅵�Ha�¦�C��7��Fo�<���N���9����,} ~v�I�[�f2���Yu^�����wö�J\t� o��4��R��o. m����P�w��_b��3�n��tH��ݡ���?���Fn��\��sN��8���C�v�%��������凿�����Ѣ��Hb�ݏ����LE�'���պenn-]x����/(dO�}C��e��X�O�Z[�4��@�#�Âm�T�y�Z[l�vcn�	���؇$c^du,V[�{��2ΐ��{$Ve�3&p�l�ǥ���3�� ?�۰ԃ�3.\��օ+�(���:O��,:��,e�������-^e��Zk��-��k�]�<K���i�S3�s6�|!����%�Ǿ��K�Q�-�~��4�0�Wzg�Ik��I���aZ��g2γw��R@�ĮA,������;Cw���q�\���?n��%�C�}�y��X!t�٥x�Q�SN�j��*o��D��]g��r�8ӭ�oH+f�+�
.<;d��{12?��0\m܌���]�(֏�V̗x@���?@0��,ծm�5�,�Qs��'e"�0>u���Kf.�P����\7�J;:dHk��7l%��"y|�ݩܿ��ي��l�,��Ud ��7��{�+��	'?�1��Lsi���",W[�FX^w�s��v�ƺ�嶺�,�n7��Qx:Q5c������0��[��P1� N�Y�o$4��n�yd���2��=�rm�� �S{!!>�L�$�Y��}�l��������]�aq��!�I�R��>����Z|�o�W�Xﴂ3���SSC��e�֗�]��9�D|��f���ʧ�Q󹴥,ΗS��x	r>�z����=���3��E5k�?�d�f՜�~�a'�o�H[l���9Dr���4=��*��x g���t�M����j?�z1�:���)���|�5��}}.?�����FZ(�K7�O1t��2�?��'`������O�����h˘�T%�Z� �e�ϖ���:���I��D9�,�-��'>R�G��Br�����#��X�Dh6RDp���RF^@���M�Y��CO����߼�j,]E��@�)*,���*��0���S�z�1`@ح����{ǆP쾩c C��t�ܝx�%T��<֭+]�0��7qz�q}>�+S	��\��ю�z��q�1?R��1|L��P�cK��W`0��H{?n5���`�"S3W^"��")~���UO����n;�m-C�W6��e��-�3=�p46�޿1��/��xz{հ]<�w��3�@^gY�nh�۔��ME���۬�eex��;s�>R��Uc2�c|�#��L�3�_D�n�
>����Wݵ�9�x�+�'����9��#]MC8�����\�<wq�I�|Lc�b@D�p��v�W��B�,¶��ǯ�6~e/��O=w͆��1�� L��k	��&�hS����Tyk���~)G/S8*�R3���a� 	�R-�^.�� �#�0G����Q�0���ٞ�y99�Hd��-��]���^��r��n����HV�	��B��Fy�Y��G�8͎,���q���e�k�J(A��^�_�L�uv�X]�
���@P���Knd�F+ڑ��(՞Y�W��68W�!�\�H�������,����������5�隓um� �<q[���C��d�,@M�} �S]���u��l]x��^jJJ�g��4�W�����{�mq�	���;�����I[c�T�_T� b	G��`�b2�i"p��O�E�k$��!7ʍ��
u3εRǸ$�|��:�`O�`i�SK�E,{~2�)�+C���٪v�m����l�n��Nf�C�����g�������}��fz�P ���|�1��+D��G�S�un&�~����5-#P��E�\�m
 `��;~<b]�����t5������]K����"�<�&Fc����
�郷;b)L�$D�uE[I���������I�Ӆ�7���e��3E�`�K�H9�ۅ+�z����n�y��:\�mOس�^��'H�ޅ��G7�_��&�6`P�/_��J+/�Su��M��M���;�݄J��py�����^�l�9`���F�}��[��/��Ӱ�5�YG!�W	3��nB�}�L�י�ȭ�$e�֣S��BZB�=��~�
�̥�C̍kn��G?f�Y���zt�����`��5��J!��\����Eu^�����0�TE���<&Q��!r�M)�����]azS���N�;��"��H����`�\77�#�r���3Fq�<���*ЎE7���_LŌ #�Ǹ&Wy�W�QȳԘӀ�)}[�W<�ӟ��Pm�~=JWn�$�27��+��ȳ�$7�U����N�$A]r�CSBF�&w ���T�O[Q���E��=��=�#a��NRN����B��I��8O�P���l������
c�1x�t�~jR��/�oB�c��s�҈�4�����۰p����S��l�P�h��]��s� ������6�>��O��k��y� ᫘����_q8���')?J2�|i������}%̺?n1q����f�}��K�������7�Pڗ8R��m��+_�D�b��}IFp���}��Xe�/Q�?⎙��-��X��1W��E 5��_o�vi 	~Bk���7�#�X{�RV�S����7|.z3Z^��%���~k��\���G�`�&ːPc��LA_E躂G}��b�d��Pγ���Z��g+Za�D��$LҤ�3F#�}����fܒT�����K�cc+�������q	&�����2gyC��B	&�I�g��|z#7-��;�+���l�Jy'�P��x���1-z��������I=�[]��c���3V�Z���452��k��{'C`��S_��E;���t"�(��2�t���t��HJH3t�Hw�Hww	C�t�{��{��2g��g�Zk�{fƜ`j���k�9�)�稴�fC <��{��I)h��f�g��Y�=�!g�,F�t _�6��pko��$X���b,=z"����ԯnf��R�<_�yM�<�a���z��bT�~��2Z^�h�twS�E`R	���T�����r��${6bŇ��Z�i�S[jR@(s�8G�+??�2!�7W��֋��/$��ކ��ߖ�GoP��� ֊�+wc]�i�.��5���q&�b�e_��d��"'�i7��:B �-��H�@�P�_0t�0 �J�����	�s�lwu�6<>����v~��8M�{��'J]Y�.��_�Kw#�C�?�oai9�U9����"4^");��ݝ�~�b'UN��	�ĕ��<��)�m��0X����$H{u�\��������
d��Bw�QF�6��V��>�Rw����Y�\a����=��l�ͤE!��Wn��ڵ�`�1#��k�1�y��cP����&�����Fy��n_�����4HKF ��VC=�K�np>L���j9�ȩ"5�C/�6Ө����0��Ð��p&�f�S*!�ک���Њ��ϖzE������E Mv\��MĴk����+t����$����]��7ֆ�S�U�9��c�6��xG��|'\Ѝ*=(�u{'C`�Uk��~Q;���=�t?���D�x�ǻ�T<�{ƭ{S�5�1��ce����D��|n�k�rQ��Qn����/	�`E!`ŔV#Λ R�@����v�����O5���P�p���Ȅ@\���V�7���o�YJV���I����l��8Ј�\f.�Q%�6|����u	{�Gn�n�r����g~
u����呥���f���M��1)ۂ���o�V#��W�0����ߢ�}��^�L+t��54��/��xA",ŗ������f��o�+�<��^}�W������2 ��|}�e��L���l�Kh#&�7����6�����O\G�#d�'`�ԋ��ZG�G�&+X�����8��;�M�.`E��A.q[�&�Oj��E�[Nw��^%,��j(A��-&�,��,P�j���83T��4��C9y<u�'�C�'.�$�XM�����g�2�|�N��Ab�Ƶ:7Tmł�$��dy�u�˒�L���<?�o�K��ƭw~�	�O`G|Ά��g+k�k��ۚ��E��/��쬔��s��CYڣ�E�_����a����nS��Ae��2���	b�6�n0��-k�r��HT�bɤ����aθ�j�%BI�Zp����C�:��(��~��T���뼏Y��@��
��,��pqk���� 3	�r�������D9�{fʴ�#�Z�K'yU�h7�_�hR���k�H��_s��ǜ,�+��k>�B��~��A/��ԩ)�$>t�,YxK���}�z?��E�ӃIinp%�J�c��{�t�G.��kcy��3e�A�|�!��� J,�կ+ތ�Q=�`W��@:�z����y���\�]�9�~N���m�ڪ�N�*OEA3�Y��;��o#���H�S�|׀ד\������-T�4;�Ş�`~��e��FZXN&���Z���%'�S���+l�g���=����t�<��G]�B�dA
��/��>�h��4Acz��Nr~��=�g||u�^��g��?`��P���������#��i��x����qCU��U0r�\��U���tq��xəf���^btH@�u{�t"�%��5��?9����<��fW�l��R�����7dT���+!ұ?�%���>� ��j��0]�ei���أ%��r&�|�Fք��H�mO�� ٹ��w���?�]�&����$Oa@	J��O��r\2V�X:&��(�����i�5��K犯7ʍ�Q��D�
k�k�z�k�_Y��kW�%����r�aap���'jȈ�Y�噁���<oW�H��7�nk���b�=t�S�h��Q]�����VE�t�V�Y�s	y�P.�t��q����@�Oy�'�b�V��o87=�'3\�
�5�'���[�u��M|O�uV���|r�Өx�}y�C����g��ڐt��!��cŞi[����9�ᴯ�k�`�rS��I<',/�d6��6WP:3����Jz1W	��`p�L�v^XX��SN�V�)�!�&�f[��ezC�T���3'�`6%)����^�eQ��	']q���X�Ǥ��O�Yu`qsT�����\�12&�=?^�i`�QW��=��3�C^��Wi/��QbKmϞ�S�n~�g�s��=>���?t.A�CiX8�t��Y�h�|���n�����ᓸk�{����H��O}Լ�{j�GU;O����-�30���g�gW����^�N�"3#hW�|�~�
�H�Z��s����(]��{��ǖKY[+�Su�p3F��<��A@�����=��3�����D�t5N��b��6�Nc�~�d�N���h��g��u�����}r��xNJ���v=j{0���7�u|���D���P��q�.|}�j�L9�������
�_�jb�'F�$W������oŞƩ�q��mw�� ��.���8�����]�Ac�eT����	��Z��GSl�s�r��%������lug[�Z�N�����%l���I����gb���h%�n���D�=��y.~��W��<��#=��#!��q��&��n{�l �_S���1O����]򬞚���O/5���[��o�*�V!Y�E�x���%�=��o-;�6�VD �=��n��œ�fH�&����z�$_��Fosf��ص��I\j�4*�C��������\���E��&)� ��bvCds�zj)��WD�k	^I~���ye7�
�:ś�[ݎk�H��%��Q�^8c��� 3������5V�'b��9`,���#��3��[ޤ�5���҃ˏ�/N�g���U��kE��b�F��)�e�D�$y+,8QVo/�~�a��ۀ����E��Gz(��{�B��"('A�����^����d#���R�g�j��D�"�i/����V�9�4����D5,�o�< �|��F�� �!��H/�aO#�&$QiMe���*;�&C����a�oJ�	]��K����q�^��2�B7E������J���Q(����y76��3����y2�f�\ ���#�V�Y�]9zN��g#�k��06&g�z~Q�o���P1ٸ߆��Q��}	�:�wQ���1&���(���$������}I����K�X��KFQ���W[b�O�볯��?���F��<&a�喞�]"U�a�I�&�L��`	�$�=�Y|jڪ�|D�������{�zǳJGT3�'� Ւi;V�ƚ�X�� )��9���<�z���2���9��a9���#�C�5m8�35R?d���1���j8�ga�!QP��Ѵ�!&tk:�*���8�al���n��I��~�9<����mq����վ�ϵ\�z�C�8�HH�s�`�E!m�mB�����1�����@cT+	�O���30 ô�q��P�Ȫ��ﲥ�&}CN����|2D��l�?M�]n���h��k�2@Ȣ�W������rm{O ٚ�0�'/���R0��*8�3��WE�m�zJ������7EX�?7��g{���ҙ}��4����%Xu]Sy��ԡ��P��`0�9�_~��}&֟#OS��>��񸯤�{��ዶy^ZE�D�1z���e�>v�E�P9�
y��xg�ys|1+nw;����^$����7�}7��2��0�������Ͽ
W��Hٺfi�E�9���Y��2.�}5Y�T��־�P�y�����>�;������o��;o�G���i@"��3�Pl�1�9>���Ԉ�ܮ��3�b�,�>?����ҟͨ[h	�v��0ۏ��HR����He���檌l*O7:��]�R�u?�9�} ��r8�tչ�d�~��x]��Wө�x%�-_m)�|�C�����9�$m�Q^Pa�*���%�����I������qɣ͊Co�³����]����p[����D����|��$$�ҭV�|������w%���:c�25/��@<ёF=�:��j�c:#�Q0�����a��H��_-����!�ji�-�j'����?�����d�wݥ�������l;�j��[��oa�˼����:�Il���d_%in9y8J����Js����9ʠG��pX*�s���y�!���IL
��}�4�r#_@kh�L�����V��$_B��+���62���t��n���������2��l!���bx�I�z�H��n�_���M���/�)��*��Bٓ��渼�ʯi��J{{�[�[��r���M��n��?bO��A����VA.�"��wy��g�d������{�HYf����a��U˧�ǒ.VJ���~G�4�w����G�ڏU?��{bv0k}%ګ��#
	����(/�r�]�_)�?�,��>���ϣEdf<�қ���0es!����U�.�M�Q�)��]^9k�b��L�6X�zU4�r�� ���?[��X�|k��2w��ɟ���~�IC.�#��7v���Jq�WvT悥�
�घC��
�'kT�-Ё����E���,�ݓx�gg�t������Y���i��oB��efi  �����蹬t���R�-+��NՏ#�
s����=����ܸ�;P6d��YNVrhĈPI���pO���Kvc�Ȥ�UX&�w@_s����p�{^ׁ�H�H2N����C��ēƔb�z.��f��F�N��z�\n�'�CJ���3��s��ݭ�����Lv�Ή�h��q��y	���=l��K+AKn��2!p���jn�� �@Dx]�d}_Y-u��m��2��Z��Qǵ멟��eM v˩�����*��͉���(v�y �6��Zf� �r+��:wk�+��
B������t��%�U����Ђȹe�W�C x�'k3�kXJ
D�ii 7�%@eg���ʥ�
�!n�;�0\��!�$OF������{��N�7/�ޫ���A�H�3`٩�BG��M�����
&9���l��ZG�	hlm1z|����/Un�Ԯ�Y��ݝ߸�p�8Q/P"jg2픛�5���f63��:��7-�n����B.�k�9�\�u�d77�8coz�[뚨hWC�VU1Ӎ�bdv���U����WTHFw]#�`�/�����N�ߤe3���>[;L��ai�R�?�����������ۣ^&�琗��笫�DT��=Y��2jz�&N���H3i�=�'M�.q�����$�$Q����:;w�&ߴT��j�kM��Kz�Ǹ5"a�ܬ@94"pg׳������OK���wA��5�B�x�rX7J ���!g����&A���I�i���|�{M�a��\��H�Z�<gd8����ϻ4 �w�J���-�߾[�P%�@H�ۈQ䘶�GD��v������D�����e2��3������Y%H�)%��a0�yTwr&S�76 \z<���
U����xt4���O��C7Bؠ6w�Z��?���[ֱkw�{�G�����o+׆��뀠�������!���/�C`}:, �v*��Έ���D���h>�c]Nt��(H��,�ͰO���Ԙ�ID�n.4��՟��[��C<[}P�^���ӈ�� �:��+m>!q��$�v�U��C��#���si�?�����o<�ˢ���)��\�/t�ux�f}��ֹ{�I�@�Q!'Hj�F�
[��M�>�q��/Ƚ!-Y��[���]�o�z���,���aj��QȻ��m���|;c_���@R����/ϟ甐��4 ��F0��À��,��p�/{S�L��8X$�?u�~����5CQNN˨ڴ�p5�bx�3�='����K�Xx$�0N�G[9��¬S"��~�\+�<�R�c�x��; �>�(`��66��9ڱ(���'S>�q4Oc��eN�,�f�w.�gy������z�6���~#9��Bɬ12�Mͦ���*]%�E��h�;E{A����cBnɻ6�fGϰ*Q	i �F[�?=�8F�-�	;���]�_��h������n���I�O���Pp���ogT+�~�����ݺ�e
�L�^M!�.�"���)��5��q-�qG��$��hL���<�A�H���3�a֨�R�>\����3����nz��,��E��,#�^t�=u�, �!T��m#F���@f�]�;��*pd�F2s�{�x��"�2Zf�g����Q�|�v���IuN{y�Ϙ'�Ȟ��?M ۑO�5C������2^�aJ*��vߠ�Jh*[�P��Y���������A�#�k�t�ce��2�R�� ވ�;���� HUx8Gwq�]���W׋�vL��9��NU�T�f/l�u��u����Ң�jG�]���KG�-e��r�?F��;�5���W���B��5X����[��b�x��?r�l��kG��䦖���çi��74�0�U��C�\�?�F�h�k&b^���S
 � ]�Ǹo���~r��@������ D��׮��5��t=�洘��Y{c�U�b	�apnmE>�F�c"�}M�Z2�WU]鑫�*$ �A ~w�X���ujr������j� w
�|�֠~{�m�H٠�<o�h>�g���Ex��j|(ݖp�]��4�������ϸ�Y�1n�}�T�)]k��Z(-!�@LmR��~f�/oHٗ;�B�&NϹ��U(^���xY���kV��Eer��X���� f�m��xAz��e�AW��W`��Ů�́ـ����c/�2�Й�>1��K�z2�6� �D�uj�sg�n1�o�%6��8��ZWo��̏�*��'
�>��͊�RՀPwT/ZOF��8�,�|��@��Xh��6�K���CR�#���h�[sdFĻg� ��(���^4�� p�z��z���8�R۵7?�!ꯡV���@@�n>/�!!�O������И�C�K���[K��<�3�"�TOc>�����iql	m�oo=�j����|��pė{@W T?�����A��� /<a�	Xp�G�d���X�E-�"b��G�䂊
��:�����~w%�q7����6���"v�~�,Jr�j}�#���;L�V��q��2��q���Q߽Kb����i{�Q��@4u�z�����'��'*���ATYy�vp�M �*��e�,��H0QZ�Xu�!Bg?�@R���2�X6\�(/��k����B,�j1R�N�$7o?j:���Wxq�&F`�7�y՜��]��Fy!�2�ڃ���@��y�oot�_��?( �������yt�F����3�6�4��f�O�����A�h��,���:Vj@�A���Y�f��Ϭ���y����l�h4���uX��s�����n1[-�jA�l�"�r �rwG�I@��I$r^����&ށ���~���EJ��Aa-9�ÄV*]7�q:�}��N��v4(G!P9�B6n;������x�mzȪiIp7��Z~�OT)ڜ�3�uʔ�6<s�w<g�:���x�"n��0����7��u����-5Ek�d��]���ˣӌn��h��Ϥ-,(iSt����%��������ap�˻��el�2o�����@��it�/��w3<��F9!
���%��n��@a@�:@���R����R�<�yڀ�k�\:3��@k�<̰��A�����rǤ�374��~q��z��8e�"�F�vG��݇0P�~��
�$��THI�S��"8���4F�� ��rk6�I�v�S�ӨC�j`��/P������nO����$rs�p�>?(��%�:�w��6�8P����/��L}�;�#I�L�w��L؞���<�D��i����|�T�,�ż�M�nh�g\"y�4�b�G�%F!"��g���\��	�/,����6Sx��\c����`3,Z�َ҅�iTl�#7BT3�q�DUm��Y+
	�bF��U�0�0�5((t���w�`x�p/KG`�����S�W�-��/��YG'���L�������^y@���fk�".Nw���{З�j}ܺ41�Y}4����㍫������x��V�����8�~[T���d��o�f�cB��ܲ�}���-c	�b�ka%?4�������󭍏�і��@�l>R��&��t)ǯOh�!�&���2�0�� �N�������`:��?���p;��0�0;�����Z���u�?�_�BL0���f�v�_���OM��\%$ȳ�S�zQj�<�sA�ę���ֵ3���|�r�1,��@%���'\��6ʟT����?m���3��ښ,ѷb�q��^�AǎARmv�_L�O�ne���nn�B䚍����C��q�= ��#ϔ�6��������C1c�F�R�	R1����e%G�V�H�)���GSd�h�5�3H�n�|z�5�kC���E��C�='����h�v�w�K�r�o��)0c���"�ΰ�T�|���`(����\2�%�vڍˮ/���W@�L�?�|�h>9����:��ׇ�]�G%����.��x�6_�H�����Y��&b�Ƴ�@��)*i�T���j
鑈�O���<}Y�>[X uL�<�Hr�o�|�i��|LƢyO+��ɜ�]:f���^����kGwzY��_�I|( �۶�w��j@���їvRc<�l�ltk�)_���t'7��.9�;������^ߛ}����+;�zP5�LJ ����>|b��R�h��,��v��4r#t�a%Q���� �X�qGڼ~��Yj���DR��i+�41�MQ�t��٨#ԕ��>jO�Yw�#I.Pg�u%*����{����L�ȈQ!�و�����;j�ӌ9���8Dߚ�,��j�BҖ�ܺv+X �B�1_Z}�[vvs"&:J�h�����r/RQK���UNA�3 ;Z���o��lL쉏eJ2^�zO=�,�5�{j���%����� N�����O�4��{�&�؋��q�@l�#/���DNw����>��%�T�=�u��g�6N�4��f B1��"Gv���*	�瀣A�Ayj�� M&g!�;{Φ��i�F9���������|������X�f�z%�2�(<( pʌL�pt����w�*��H?{��V�=�5V@z!t�Kz�]�a$���1�[x�v�q�w��EA��AH$�=��B����N�s�)��(-^��;���^�_ qG;��a�𭨤i���[?�^`�D�a~mW�o���9�c#W����P��7�f���E5�ʍm��{��P>�xg/�ӂ?+?���%��T�|q4v�������]�x��.crܙz��5Y����sUG+:M�k7�����5�x��ʯ��:���	���ܕ���ԣ���� u,-S������V���6�C%��&��@"�-�X�[��'z���O�`�$7�:{1��zNRAΪٷ�&��Iy��]AoX��d0=�ϩ&2�p�EVU��u��Kнy7f9�vU�g{��ƑJ�,�����:��N~*d�<N�RW���{���~A�o�ΐ��y9��Y�UCE�ج���a{	�c`��x�F��?F\#�@Jޗ���X�)o��v���L����'�q���u���>�n�N���)^��q�TAYh.��l2�Iz)
Q�${n_Tv�Q��+�ϊ)��y~���Q��$v�.�uȾ����%Ewy��/�a)> ��լ�l��z(��oTb℁��1� ����qT-�����Hv�%W %d�zg�2����bV��x�Ǜ�O��ú�NR��h�<�[p%Um�
#��h'P��'������l?�GP(x�i�A�T[F�	�*����u_C�D:E���ߏ�Ph�y+0�q����ְl�o�!������V���s���M6ӛ���[��ꋣ=��^#��3�$�F�s_�����x�5<��z$�I�P���8CG��n��s��9���TLX�.�硁�'L6��eN~#���u�	�91��-�.���\0Ӷ_ǥ���x�9�ůhH��<�A����m�H��p�8:B��p�hۣ�=��^o
�⿸���[���.x�-�Qq7�K���r����3��Ѩ�S��zz��.3>t�/eZ�u�م��خLI@���p!�F��6�Z���K4Odx O=���t���=�<`�|O����1�ln�	��U� d/���a�D.�A���^)�D���ɰ�����9��Gdi�#���}g�ʼ��9΁ȹ� ��	K79�u�R0}�D�2h���X�H,�Z��a ���A�3PzR�&��v�y�G�y��mEM�z�q�zLpX=�~���ћT��}B� ��+�<]u��}5������8�i���{�g��Y�k{�����)2~�摶5�� �H$�:�)!�ҝ�S�ed���=
��x�J����"O3K�D3;v�M�� ;�ϳ�^0\:48��LvV�c���$������[۫�GW���[ �/����B�]��~E�SZ��t1	�稟�m�﬜����̛q47����oZ����5���y�f1}2p�������j��a�T�(��)?�E�oԢۤ�3<R[zK'lID6�CI��
F�$���%,Ny�~xT�[��&�6MRV��N�H��i\~W�3��~�'��� I��8񇔔Ժ�_MH���9�]��� :%%'��2_�Z���)�a|Lֺx6�h�->�,X3^�߲*
=S���ix]����a�ZI�CP�i^n����?�����3>��c�H����N�c})X7�+d��6�	���Z{�9��%�����\�(��JG42Q|w�aJ=����`ũ�B�ˣ���Fv����+��	�W3���G��ОQk�W��R޾7��h4ߕ�xf�m\C!�m���-��|�YuP%�V�0|/Z�����O��U��^8��d�����3jb���ڇe�p9�c���n	����D+�C�lF�|����&W����f�J�=o���4���z	D�)�VZ]t�C���-��;uƮ���;q �^}�2m9J܊���>Y��9� �A[�a*�H6@š2��V)�(4�zr2u_�1�����x>j��y��}�t��ʣ����u�9�1���A��o�X�|9~��1�'���fQ�P�Q�z<z�O�P���YWz=�/;A��z�/�<�hi��I�1W�y�:�w�Ŀ�o����ٽ��LoԚuj�t�_Wy��ئg[��X�6�<C�D� ����l��*I�� 'a��ʝS�v��/���P *ވ*����.��o����;�D�1D��_���늗�+Ƴ�^����n�2Mڀ�}|�3�]��")�Z�����7�u����ޕ�=0[��W%1�&n�!������c�cV8Z�����:s����Y��!ro��or)X��(`N�o��0�Y&Of��MZ�qN�C�������m,G�w4�Q���	���!Gs>�3ݓ=~��76�g�s��И�=�U��o���Ã��5ї�L��E���tܧy� &��=��`����F��5^v�����n�(^��1TK�F��o�}��#u����*����ArϩQ!oȩG�.�I�j ؘ�8��u)��Wɂ��D0<��Tڋ<�Z�0w��8��].W,��}�X��um��Ǵ�֑i��Fe^^\
U��?&�
H����4b������-?�")�N��b����R���o�����{�1������z
FW���x�䠉m�J�#߫bI4�ɢ���f�
	�ZgS�5�|Q�~5�%��=M�Eju�W�b.,��]%��:�w��i�!�8��y�f�D�-@��y�l2L�J�~�M�p������Qȕ����� .��8���@�3@zA�-"Хğn�XH�m\u4�Q����*�a]�Ml�ʇ�Z�\<��������6K�Ʀ�+%�P�S`��&?;J���S��d�u����m�J����qO���b��b4B
۟ �� ��ܛ��z������3�����h��0��[#��K�E2���B;�����|wޗRr{|�~�ۑ9�z��3Ƭ����#���~|�v]�o�hb&�IE�{?��D"��aE����`mf߂y+��ލu��S�ʵ�}5kņ}=�Phd�N#��Ff���Ov�ٜ�ͧ��G�Y�?R��f��N;,���(<pܚ���kr�z�Z����?����Y��M ��f�Q���&��� �U9���'� /�qj#�h((K&I�V G��n�vm���S��}���hWME��9ޠa  |a'p��>kR�.��O���t�.�>>���D1��m'���Z�]��?��B�͵�܁���at$M�7'�����2��*��9.xsnF��Pa�'+��7�"T8=��裨/ˎO2��u`��fs#���8SSa���6����.w���	}����f���eg���$\L4��a΅��m����*�z�>���=�n���*J"+���)d��M����U`P�zb�>��v��~����ʺ�}��>}�A�⛑c���{�E����w�M"���/�X�v�_�Y�U���s���Wˋ�
�u:(��&���q�K7�n˒�^���fdVEţg<�! dd@ί=e>;�b``�U��yٱz���'�ms���%7>>$P�-�f���j�gF�>��\�/�C椊���t�YC5 ��7e�6��m<��W�&eߝ���<�'���m�����i�4(�C}"jj>���/>h�Z�:�n='[M��ų�Jp�n�,�*���f�scʋJ��<m�x�re��]�x�X��!���!�5c�=��@x�����_��`��Rsm��S���޵;s��%[�f��� J���aK6�@A���=�,�����6p�%��yX�s:���}0cN����O�7--
�ccszT�@u�q�P�����ٴ�,gF�߳���S��Q�6�G�[p(J5���ȳ�9m˾�d�\��y��ܗ�.[��)M#+��Gр),<]c�����e����U�(t�mJ����}�ŧ���<ER[����p��Os�1�c/����Xm��=CW��Ã�P�5�^l<ؙu~�.|��<#:/����P����8����fQtgk��gv����D���8�������`�Hj1�lqnZN�ZR�1W�Zm���"��|I"!�N]P�E�OY4��~��b�2�!�?E���ֺ�H�2 3X��ރ�����贸
2�����l���d(�8��2��O�q�G�_���m�:B�/GT=�fYH�n��o1����(v�O���Ne2��	v�Ǟ�er�@n��Y�;JH	BI}2�ҢikPwk ��?���S�P�	s��!|�u���wn�;<�KI�
��?��i0��-%X�vM:��������?��<���z<��D��퍎��9:�ܴ�l�;�SfI�D���F���L�v��a|8�K,�:��iWZ�K�o�`V�Kf��h��%�qJ����"����~��:Ӕ�.+kC��\��A�i[*��*\8��BE�0�}&� Z;��֝�UTa������� �_hɔ�08��P��1&.ePT���Y���O�wr�)�OҥY�KR�RRe`^�( �2g)�;�f/��$��O��^L�W!h&H��� 煐(�Z���}4���rS��K��`�	���x�"�DCq/v�~�02_U�G,�Ѫ�YN`���ak!BJ#���)�Rt;������k]�������Y^:>�fX �h���t|��s5ش<沈8e�8��rP����K�O=Iϖ�85.�3�.t�i�	�<��������v���CƖ��/�~�e��gu��̜�#��Y�<��d��Zz킺]����)�3̇$[��3k;_����Y���!J�Q�K5O1��M��q�e3v��U�>��8���-��yGn�uN�D��υ�E`8�
��dj�8�F/x�:nAoJʟ�Ҏ䘒�.�:��Ƈ�c5�jh����X��q��'ץ. c�K�?� ��b�����95%#n��j-	u��V�Ұ�+Q�g��T���|kiA��>�5�ʆ��O�|��s~c몕H����<��4|I��8ʓZ���=s��t�G�	�L	�z�%�$��ᠷ��K6t���;���M"^����s�Θ����]�ͥ�?�����qfY_�u��=�b.!~$O����Bo��!7��hW� �p�l��
l.#1z�"�G���)"�6�s
��"U![���{=5���eUyR�r�?��+U��h��DB�!<���a�|���/x���v%����X�[u�U���N����U#�z�e��'�+!Ƹ���9��XA���ގ�*���}���W��D�5�:q杒#�q�Φ&ӃY����/I��@��[��c+�05�tOM���q�y���i8��	+|@�߮	��	f���)"��kkk�-�/�M�ab�@MpX~x��t�$z�(�G�f�g�棌�(}�Îu9���$L��>f����9E������S�cO<��t��"�(�S��s}ˉȥ#ɺ�`�����U%J�y�#o�Mʃ� �R@���:�R&5�<�z����麬hO]u��$�oK"�����3��c��k�%������1yb�*�G�CWBA���w��z���=o)suu���ZHu'��٫olw��Kٶ�-��o2��E)�����~�v0���;S��ym%4Qc�Œ?r�m��|��ӭ�|!$!�����7�n
�?"�z���,�!���!.$��$���j�.�J�uix8��@�_GLœޡwI�,v�,Z\/vD`��O4"N׃$�Iv��sLw��0��C��?�4�� ������̺be�r����y s����)$M���1%��y6��BPa�;a�}������a�ү�J�^�`��E�#p����z���V�76�̱9T5�\���6��0{��e��H��5E�ddM3�b��F���ri���>��B,�ⰍF��	�������[�^�:c����E9�:�kq�h��r?ry���� �Ϊ�/tl:�5��&�)�`��F�o��9�bq��p������ jT@���ø_q��͘�9�&�\������]�3��Ƞ�����HI��xC,x�x��!P���#�y{'!�~^���Q����<Z��*��;�r�_���t�Qci}V�����˞P�(쀘_s����=K�~��Z)����Q7���RI�����;�+!�9=�	p>߆�BZ�.��ׅ�eo+��n��d���F�U��:�.�11��w�;����~x4?�AT�u.�5��ف>i�aI����ヂ�h��sa[%�t�r�H[��W�]�%	�m����Vb��$�&a(�UTw���e�Urn8��
<}Ϛ�6)!5������%�&o7�%��;�;s|Q]%�C^Ĭ�U�f��;F����zؾ���#�v3�42n� 9�q)đ6��(�0��Wp�;��&l�|������*�<�y^�1 �,�蠗4�������7)��p�9�w��B)5���c��0j_@��(��V��ńu��� 8/�)
����YT���y$)��KM=�mMz��r�B�V�\tDI����<%��i'��@�V�y檜���z��a2�"�.~�<��aS�,n�Z<=����PE��vƶ��dd��o�"�L�蛏i���]=J��>2f��	6���W�;�_<�ij���۬�XsrB�F�m���Q׃����-�������xϋ�c!# �[��O�k��!�^�W�[A���.�":ۃF�� �+�*�~Kr����
���.J��ˀ>\�4�����,�I.D0^ `Tߌ~�DR��%��)pǭ��T}&{�ܶ����؄�&���ڐ"�k�_&8�x%��#�:s�Q$�h�i�k���CV�QC�K����S��m:U훖�jd��<ajƭ����!fneݜF�定�15�'�'�bǔ���)� >����P/������#m��_�;���L�j�I.2ԭ`̟lO��3{<@EMM���r�xF{N���:��՚q���-!�����9��M�~+%�T�W=||�쪝< ��m�_7�̲�e!���а��}S��F��A�B	� ���R�����)��du3��2�yw�֞9ק$��weh�]>Q��[��Lx���{�Fg��An�Up�I�O���h����a�����'ĤHv�}�t��U�f+�sƐz������2�-�vs9�)� �
��O
������*0|ȒH:e9��E!q.c�?��P�\��0�����"7�U`p �f�p�9��t�?L�갟��.C+�u��,���b�cKG��.6�U���9�W�/�6X*���k�4�NL�B%z]=�p�a�Id�[�f��;��J��"�.�$�'��f�:pUsW?�ޑ�N� �|Mn&�ZuO��z,ӵU�	q����:j�aB�G���&�=��^�n�$AM�ğ���i��Ȁ���gql7^�%)�n`�o��H�=�(�wCė���=_yW7�����H9�C���Er#$"����Ԋ����i(�X��6��o�l���Ё=��zf�1���r,L����*���Č�r��L<(U��/S[��>�>q�QI��V%va�}�SKF꛾��$��G���CZ#�(�=\zNX�w�dε7[B5�1�=`��@:�

=�)${/����
���7SU[ܽ�%��W:�g���A��?.�P�����}��o��#]����+�7���)�t�c�*�c��t�)��4[ZE#�2�ƚ�]���4P�Wc6���](;��^���~~ÿY���0-���{�aA�Cqȃ�Sψ��z���.lXDA@@���S�[�D�D�d`hP@J@@��n�����c��?��|����֚5�a�����}]׾��>\�u��Z���Vu�T��u�8������!���+/�������j'ea<���NKuN���S�#7=�̲��V� ��		�C-p<�ʒފ�B��?�aG3hb��������U�=_��}����P�l*!,W��#
$�,o���i@B����L=I�٘�V5_�ϫYU�Ze��*s{�rCq��3���R�gdCKcfw���//VA~�˿i�9�!��>��qc~ dJ�y?��]���U�&������I$�-�@x��[6S��Z6�:cTTԄ���BlJ�(��ar(Z~�*q�rvF�j�a=�4�;X�xxYJ��k��2�V.�,J�$���fDE�$N�.�$��DP;�hŵ3�/~}<�:�ɱ���LgX�}�;&��$��l�+"�\��Q8�.���K�k:[��#>����$�O��R��Mk�������D�A�뫍��!F�H��*��8x�cԂW�x .���y_��GלU����恟f�C'*�g��˽�����=l��C��B����ؼ��l��`�L�& r?�	�S�s$�\k�$�m5S��pui�Io7�˙�5TW��v�&�J�������LE�斥Mf��?^�n���p�]�9��<�V�<8?	+ϧ�ST�U����J��Q��vf�*�Wܒ�P�zȅ��������� :!��i|�p��hy��Z�5��=a1�<_������>k��,�⿄��|o�������N&�z��N��ʯ)�D��L���tq�ϐ^7�^Z���;�u�ퟑFsv�ݯ񪟪\��"����/����hꡖ���'�g���
)|����z������UB ��\<�-�����oa�0�q���U
�m����X�}�d39qo7;�acIr�����X���{����1��]�D�'B�qٗåa�73�C�b`�`���D����~mǡ��������̠vT�YK��t��5S�&Q�K��q��}Z���s'�I��t#=.(���N'�A+�X��S�٩�Sφ%a���F4.>K\�g���˧Uj,'z�1B�H�Ȇ���ug�I|L��G�R��k�{G?�  ꝶD�����ձ�9�ޓ- �]) #��\T:��	�oϮmG��O���.4����8�1����NS�d�:���[��Y�E7�v
�c�ц��,����B��;�/�[W�8�G�;�:Ri��l\%�KRa����w��4x	p4�&q�֭�U����
$)*����6�Ӎ;5�� ��do�94؇9y���q�^��e}�^C�q�f�����E$\T�^
��y�I���̢�gf.*�韇\�vX�a�/!`��J���
�:1� �2+ţ��2�C��znNO�y��s�kf8������H	Z��裫�	��Q̣�=���UU�&~9��	`/�u�h���ck�]���N���-�xA�Q�d�ϒ�	���z{T���Lu�V�pE�ֿrV���ok�!e���Ob#��_�����v�!A�M_w.��	�8�3枙%g��C����m�-�cF�dN(�\?M��7D=�@�e;'��
V���a����`�7�Z��%O��i��{�qv�L�H�1� ǌ>����-�'|�XۣϿZ&L�k��@�ud�ݚ�0 ?�08��W��3�Hw"��6tUM�@V�By�/)D9B��ab��<�*�[�.0� �� �'aM���&�z��K��L�L�VxVh�N*��vŔ?�����m�󥹐o؊��{�'�'������]�O�������w��%}�v����j�l ՝��)� �n�uE��r�ߑ��?nK�Ӣ����Z�a��_�46�@�dr�hS&��:/�D)܆i������O3����CwIy�89�MSe'h�+����*v�������I��@�')j�^���gڴq�`����bҡ�ݩ���K����a|D�(֋d1�7	���a�* �j��DM���l��Av�D	OI~��r��>/���JbA�5�W�ܔ�gA�@J����4�S2�7��YQ�ӝ��LaJ�*g�g��~4?Z$.�U��|�`��{͇%'���U/��>�W�v�?���T�`�ZH�H"Lh�T=����Y��e��f,��VWL��(���9:ύ{��5�n����j�3������M�W��(�	�ff�te*�z�e������Wh�C7�CPz�{�D�+���׾1A��`n�"��[��<Jsח���xw�/�X�r�IU��4�i���N�8#'\W�J^9Y��1FK�Z��<�7�P\e.>,��g�a��?��M��I%���cv�|^����,����%���T��#a'����ka�{��~���s���Rf�K�����J?��q��#��
¥e������!��x��eg����8��LW�.W�(	�FU��5��3�K���*`Y�g���޵�J	湸��>��ez@X=1��>n�����Zŀ�0�ڃh���?�e����, �^���u�Չ/F�(���i�q �MO*Ĵ���2�r�j���j�@���
�}��k��� &�ﲷyr�KI{T�M�Rg>+��y�C�)'�Ѽ;Odǉ��LN���m�P"�D��a���X�ϲ#�tZ�	E�c6�%��w��?Y�R?�k�����G�����`uv�e+���8T�-7eV���,�K�R���c��$#��)Y�L:��m��NK�#�f���k�;G,Օ��*�o'���29HԶ��^�@>��\�)����N���#yW240R�'k�B����ym��ƟqJ�+��?����-�_�,6��]��>�����3�Z;:[b�~������aWr�t3�=��r&����ԋo�Rj���ݥ}���4��¾/ofo�D��G�|n�l
�a[Ź��ݬv�7��x.f7�vȢO����LU��K�	STL�dmfA�C��+rȖO<�*����l-:���c�f�%�QPb�0�}���fZ��F%����}3h��V��K0�t;%�-L;�E��� JM�M�4࿧4@��h8���Iq�?��ɑd�������!��;���3��o��r�Ӱ�!�cMr�.b^R0�;m��q`���~Ba�,[�g��JKѸ'�̺8�
�7�����m��p�w)��?E�ΌÍn�p�>-�����|��[֧�@�W�xJY��q���z����F�WX�@�Ym�e582�J��s�7��{�y���*q� ~vQv#�li����b�7�K
,�abwW^(�D>L�������������u� ճ���Ez;�F[�K�1F+�4b2��iiAU,ݹϧs�.���F)�1�
�x[a Uя_H0��+p�@�/������N�[/x�����
Z�ֻH�@�8�o� /Ltw�C���ծH�M)�����'�:�	�$��d�/�3 �H7� 4D�vTQs�M9��Hs���2�z_i�-�gFb!���d��O��2��P����=}�z�oFh�b�]2�ﾪf.	93�>�����b(y�ғ�*,�RF}sв�>������-�{Rϻ�-�#ذf(�}d�2&ל�s3��_�D�����K�%���y�A2<z,�o�1�D����Y�/e�eA2<db�=�gu����|�οظq������T��/.�E4�֔1v�kiV��eD�I_�� ���A�M��p���"�'��-��*����Y�d���N�� K�3���ܾI�i��v鰏%>�Z_���?19<���!,��㲜@���y�s���
M#F��7��_��2�+�NT�͉��8*�5s�ι�}+f�0�r�R>���-��������D]*O1�F��f�Fj	�I{_��A�C5���\��ɭ˴߮�w~�֕J>Oؤ�>1��%��<e�4��O���?+��tV��c����� Տ[}������YC�e���}�T�W�n,��w�AmR�j���<����Iҗ�A��=D�G:�a�a�c����Nʧ�=���l�a$�!�����Y�L%�8� �O}�Â>�+:�F3L^収?;��ev��H���_=��Ind�O�mr^�v=s1�뫰��p-��M�Xő%�F�t��y׃cY��aY��O�}��� �E6b�G����A�5�d� A����M�_�fw�2R�9�_Kk�{�:���5Y�������U��R��!y%^
@��36���6y42��̃v�(JU�l�[0���B�5���y�R�G������)տ�,�?�GXZ��4�G��|�촌��������!3#���p����A����],y܏ |���Z�G)Dg+��͔r�1��gvw��ر�G�unu�D�B��������hƊU���`J�J2<�؛U�9���]*�Q]�sw1Ox�|�����tSm��Ʊ�,���
�3��a�Ȗ�K�ڣc���U�7�!�?B;��*���tvX��ې����W>��F�nN�ŠN��������ytx =�IM̀��"p����-�?h`��mJI8�1@�<9&����)�~�ظLǌY�$���3}�#Xq�Q����LU����,%�x��a�`ύ����:�s�z֬�k~E��p:��d*)�`�AM�i�xBm���
L�a*����~6��l� Sˇ���� 1{�M�Zj5���F#�+���*nulFw�ƛ�����H���� ��r��L󣏖I�kqm�w�7?���^�[��̡e
o����;LPLi�oG�@�ڛ���&���N����gR�vN�Z{.����� `�g����?�c�?���Y�Σ�jM�x��y���JD�fZQB�y?�9��B��F��S{��߮�����j0�J����dn�$o�W:�kw��"�B��Rq�&n�Ҙ�{��&JT�� ��|�CS��)*��H���._:h� *��5f���"@�\h�"��M����8|����˷b9r�v��+��"�:%��^�r����	�\�(�������,�t&���z �j7�r��$ڤ�b|L|�~�������LB!aN	�z]JPm�s�h��x�]m�S
��cG�W�ҳ��?�+��:�����&���8����R�4?ِ�uNqJ��~z�i�P[#O����n������v�ܦ@����.��Ô�4Y�����d��U�t�d���[�:*�Ѹ��v����Z��=մKDIj��+ZHi�˅^��
e��-7?8;;����U�Zw����cK�Er/�#��E���;<MF������k�<
4��ܕ�sC<E-����RL����K����F笧�4:^�zza>)��̏#�oɴ{�X̐ikj�b�����io}���ύ��Q��b����9�0����P���+7���t|+[rD9�64/�C׉oOlw�}_T�Rg,-[��p�9�<��g�d�+>�Ķ0�#��N�A��40��v�ދ���Y��F��s�S7�d���nߕe�Yƽ���}�d�)
ox[�6�o��c_7�3P`!�+����k�B�m|#�I�|����W��e���|� Z�S���Px�	�f�a�0����'��;��joD}�4LE�	i��Tf�p����hX�!������}�<��;�[2<�=q�I���e��x��Q���&�Y�U���Ȟ\ncd4����*�����^t��|����:`B��]Je���Z�$�*��/����ՆӁ�g�K��&�]]<���ˊ�--#\o;�7���&ja���u,�f'_��#�Ϯh����.x��������������L��,��tN���b}�iWN-`�lzB�n��~����E�j��b�P?�Ι��.��OW$y��!�^o��{ܵb+WY��K���V�5�� ��k�)Ka��΀���� j䕳'�C�zB�]�K[W�-�H���A��)�tXa�ȷ��N-d�%�J�ؑ���O�b�6'�@��D�U��	j*���v9�<�5.�	��K̐o�.����-�����Y3F;�CaYJ��o��e���;�&���7���>N�)�@�[�ע�ʜ�;�J�t�[��
�:d��>��{�I��>Ȯ�.[
Knۛ9����X�� �����ج���v�t�-T-_YĽ��Ut��~�fw<@���;
ø��
׿3�.7~�}~��u�7+�A��W�K�f���E��'evb�z���DF?Ye�_=��#a.��[4�a�;�3W;d9vO���k5&�NRNC�o@7�3�;��asj��������ڛ��~�����V*���I>�u��g��)��Ll�;�h�:��u��oY��z&RL���;�ø�ӆ�'5��4�NkL���h�0���gY{Rc�C=${�DK��p#�!	�޷8nb륄ֶ�_�FIZ���i��P��e�KG�.��j9B3��"�ګ�o�攴`n�2�P7�=Q�����Y��Ҡ2�n~��dwس�6�bY��3U�FX5>T��ǟ\H�m"��0_��CV�A�=Ƕv8�a틍'W�d�/�i��7�_�(I<r�6W2l�I{�yB�O��\�Ҫ<t�.]$m�9��~�J���Gz�C�H���F{IO��=��2P6^�ɤ�9�A0А�*�!-M
����޵��?� !�YI�{��f�U���p�ulJ�Tȶ�]N����x=G\�1[/.xK�ˢ�>y���NS0�%�)��O��c��r|d�������X�!�5�(���s��Kj����}�h=͠��[��5Z�+���w@D6���l���qHj,W�M�V���u�x&�/�x����~-0S���Kz-��T������N�����t5���&�j��W����2O^jp�w~�_�8�m"�t�Z��C����1r��^+�Z�VtaӸ�lԉ�Z۵�$��D��S����7HED���Im��<N��'M#��\�#]�U�|����	�:��e)�)Pp�M*A+�$G$�"��	}�~ja���2�d��
?������m�@1/O!�3�bҩG��a���b���R`�ֲQ1���%tDs�����Ki@�u�d�k�n�xQρ��`���a���0�Y�������a���t�}�x�1���ʌ�
��*�~��?�W/Ϣ�An>웮��g�D!.!H9aG��_6�`��
��,7<���z��i&�{�����zZ� ����ŉ�����Ҽ"D�.]�zc#yG<�,a��z�����x@�i9/�('��A���2h���a���Jɕ ��,��"�{��A��l���s�[tA�+BjǃY�pNԣ�0W�G�f�$�{����ߌ� �:,�4cC{�K&�lz.���%<��n�C+f��k)���:}Z�^8�:F�����CY�J�q���<S��w�����I����4E� �8#5&�Z����E�t$"E���P;=�q�<�� o���ă��3�
o����eAYg%?<O
'J�[J�3�n����
M�4˒����3U���O�,�iٙ���v�?]�B��}�c���Y�?�p�ԗ��UJ��6�`,�=kˊ��C�6j��e,�u���y[���ȣ�[֪d�w�cs_^'��eM����ia%��՚qpc�:͘��p����`W:�t#i�����@
j��h�u����C�F��(�{�֙�6��ɸz�|���B����a.I�j6J�_��|I~��U7�`��E���*p+�ퟠ��5���Y�RLzj���7�@��K=���ٳ0�qױ�4��X�
�B�������?0@+��J&�F�W��܂1�X�� "8�\.�Ʌ��>^R7af�̨�
����]��~����T��ـ��K�	���Uy���}��]�x�u&PS��FDVivZ �uJ�?���E_�� (�w�'4�03����|��,F}������L�rk��?�Z/���g|�S��2,���Y��=i��Xe�=��G����̯��-b�����"�g�/b�f�Ee��B6�g��#.K�(���B�lG�b��7�UV�,B��ܥ�Q���ݔt���=��7��������h��Ւ���ߋ�7@ �Q�}2� q3~��~���KB]U�q�?T:z��1�ao%�I"��TF���Ό{���	����s"��b�3%I������!F@mpbȾ3��Ikwt$I��W�������xz��}M���R7��S���B��l��@B�/�l������X�s$����4o��0����������0¸���ͨ���ER+�{j�����qL�1xѠ�|(c.�{�=���1~�G0VV��ɩ���FBT8�jޱ���>rt#�X�����c�=�Ҫ��,m�ԛ��OFA ys{-J�Z���r
(�Ek��~�l=I�Zi)��W|�H�b JbKN@ڶ���XsC�*܋ޫ�1�_��[���O�
�O�gLm�A�<UKc��h��l^���
�g]Ӕ����?�$�^s	U|NG��Z��>$�5�I�����5b4��������\b�d���$Lq0������.!Lk0|�lD�ѐp!Oc��K�~_�{D=M�L�����R) �����LR+�������<�{��0��kP�V��] &:^��umGC�3r������Ȟ��w��zb�E�4]��~ �?��a$���bG���+��.�yx/��WwE� �V�j�NW�=��9ߍ�W��o���۹ā:Yy�� };����jv����Yf��h���D�����n�bAC����٘�0B���F+��QD@�d�4��:�ykX� ����S�l�M]������m���}�H!e��̑�"Rd��c��#�vc��cCq��5�Qc!B���J��F�)��<���-�����~x��u�=���J�MM� P�{���[�G1��3$y�� �.����>�E��(_Y����v9���N \-� �$1�����7�L
k5uܺ�/���$"�Ne��F�=,7���3��I�d����R���#�߲n����p�g����l����Ѫ�C�Zl�(����ʞ)����~�;����E߫��|�n��t��Q�+���.kl���D�Թ��Rz����1���upYu	��X;@��إ9���nd�=�<�8&g���(���'�%�a�ҪbK���H@�����t���p��%左�za뾓��F�>X#,U>:1��,���&O:��C�*�Թ�i���������3g
[��p��.��8�k�������X^}dfl���R���<q,v�\-��@�(������������>�c�V�@�M�k��A ��#߷w㛾��Q4���+	uB�W��Dw����y��O������oc̥�p� e1�cU���2Kp®;bћ6��k�h��֎��Q&��s�D 8*���DMӖ�"�QC�ߠ6�Q7��o�1�� �F������Kq�G��GmrT���d�L>jY�GtTj|c��6�.�EP���^��0�b�U%���_�ƚ�iHY���x���� �� �4u��}�ʳ�\�Qp�s��'���#ٜ�>�;i���|��y�>��2������,��e.�ï(&��"�i��(����5v��u�����]��� �zc�u�o�nh��2�F55�ZҎ*���N$ꬷ����SҜ/|m1����I���~0W��9%/���������I���4�`�h���g/Ŕ��=zKP�f�Y��S�'&�6�:ab��Wll����N�2�ND�.4(I�ʳ�v-�NP��-�?���XS5���ǃ�6(��M�|�Q'�6��$�J�P�6�+cxk��Rh���w&���Bΰ�������/�~�#�'����&A����l�0M�CD����7^�,��1;����(%]J�dN��
	K���w��)n���%z�?��ŕ]����oxh�3�i3,���]�Ҵ��K%6B��<����82{d(b��j�qP�T�AF��N��VQN���'VJ��?=*D�$yyG�_�.�8v�2cQq �'n6��g�I�N0�}�q,�?Ʒw��1A��k�F�ly�@��ZG����jޢ��ڈ�?G��T��ΑeJ�O��=��M�L��?~�H��?@-��5�砕�L&�;�=�"F�dҋ�w�B&�%xG3ކ�NZ:�_9�Gif����;]$a
E���>��Y�(�*"���p?�Hy�԰�p߉dv�0b$@�_�ŕ��[���U$φ@6d�G$���ўN(��Ƥ7_i��
�;�t��(�[K�@c� �v+�"T�'k���C���E��	��o�ҥ�n�n���0����Q�]�k��~��2N*��y�-��Z�8�8�Ɲ��?�	I�im�����}����ߋ�tW���H���p1f�  �͋5���}�֍��[v�kKZ�7��&����ν+]���Ͼ��`2qJ��0��Q%w��ѐ��R���0b`����ͮMd'3��}���w­�CQpŀQ{|�k�:Z��;<����	�_}�~���Ƒ�4!���_f>3[(4�5��cb�3k�s�K_k�M�M\����'��F�2��%�,(��̛�TS؊6��^2��ꐅR�J�hW0!$�['��-+��E��{@J�>�����p�BY����|�9��a~tB��AR����입\�5�'Ի`�P���]\����8s$��ތ�����\�hkb�/��ͺ�3xRS�[A��\�	��gfV��?S
?��������O��(�9���{̜ɇ.q{0����Qw)s�:�g�	7F\4u��+���>ľ>f��)..j{Fn�"�Eu�c �����RB�)�D�v�R^A�r�D(�8����/�l8��<HRƭӋ�Q�N�����k}�����P�o+4H��r5��V09�}R�m�Ra����Bv�6� �pe��gGp��{��y{6|6f{;KI�R��>�.��Iw����Dg�T���a��(�i��e�Q�挲��/�3�7�do��.1�͎-P��wY���	��s.v�1/��	�׎����W�a�ũ{�{���{^�ںۯMzx��V|��f�-ݳ+D�?u���RӮF���?^��֯���z1��o�L�Wq�M��́��ף��9�d���\싶?I7J�ҭ�4O��6
���+��S�$�2���������3埭q���ߊI�ޞ�
ܢ|n�oT�Bm�6®]�����hZ^rw���#۴!�ȫ-�������)��+�p��:q;�&;��j�(�4�;�ţ��@���f�DH�����x�>�R�r2�$�~"�P����C0B�J�4�&vT�
>4B������:���G�y�FeQ��W2���(���%rqS�w6�;6��]Rէ�����Mh?L�j��6W�����P�Th����O|�C�2Fė�f��V���	�QV�����F�G�[�Jy��y[3��-Ȼ���?��N��r�e}a�Wsԍ���#hb3�� ��'����$o6/~6�/T�毹,lm�f�T�۽m��UG�����arI�9�I�ӑw��.��qф�ඓ@��o(tM䈨� �4KL�v	�7��	S�{���ܚ��y�A�OG�b�n�[��Mه�����0@����W��9��5��[EU'gn���,�o�'�eU��*��|oj�gr��������~MZ�YD8@���W�ǳ��Y
l��� `�u�"W0*2�6��2.��_Ǟ��yO~��������8�nV����n�i�L_��L:��␢��פ[1�����lu���wSwzx�}c��69P6��J%�L�8a��	z7 d��5�~'y�N%O6�'�p[P�:�*��B8�vL�6Yn-�I7�T�u�:Ex7[TL��\��Bo��
�t�JZ_8���j2�+>�9��$�J��Et�a2�$��@s���-���2�	v,��}PO���.5�̅�X�XR/��/g��VzYP�ye�-��}yl�.@��B�\[_��G�R�L5�{�<��[��i�<=���y�m�7�4�[�6�[s4 u�Ng���5�[�wDhmU5t�*�v���L��{�ee��]�ȷ3ȕ=g�ZD��_	���jx��p�d����"[?O�ܘ���O+�9���G���U�]������my�K��9������D�QFm��NxyC��,�rk����u_�Yw�q���n�U%@��7}l��_�Q���K�ں:��V�،n�u�ȡ�h���(˽{�d�4>��w�(��Y�ֳ7�.��Y���|.HUl��a��V�խdA�P�Sm��	����L�Q����
W�y�6|B��v�i+w���;v PD�������o�ڦ�����JH��P9��ͣ��@�ml2�w-EJ�'>�p��i�T��K���1/�9�!� R�� Vz��¨^��0d{{Ga��°�r&á@��w�x���}P@��P�����sRֈ�[k����U�ơ��>���2n����9ݪ���Y��P��|�{�����x �S�ɼ��&�-Y|#(���R��y�E�gM�j�)-��B�a�P�n��n��~,���u�!�*4WlwV�q�/���Q;iE�u@&ؽ�^��[!�q;W�+F����F�a��	����aB���$�Ӏ�㠅�Q�_����j��7@ 3 �nR9�������A��]���#�o�k��{����h?f���
���}���Ө�H�	��6��tZ^zZ�8�ۙ����Oe1T����c3������O
/�e��׵o9l�"i���n�י�gmX���"KȩqeS0G	-�ڔ��e"eou-P��%mӓ�Xk��=�0���f1��cVe+��3�y�n=�����?khMq��V��s�86�/}���T[����K��6��d��wa�wađA��n_�����#���Q_@:�7,`4��x����Y:.x5KO޺@���Q95|��;� <����ݾ�ys|b5��zD|`f�3+��	�(jN`^*>����!­>���8�6�"d�y1��i]���>;�ύ{�9GJ��*P����n��1+$U�@@�8��0����V�M�x����ހ�H�#:��c/DZ}Wq�y��� x/$��������U�����5L;���SA;��俅��$\;˿��*�b��$z��~0�F��f��B|�y�}cR&%��:� ����$���R�{�%���6���m��9�����q않�����KR����TC�>ݛ��1�մ��ʠ[e��.�z��
�L�ƛ���Mĸ��<���tkT�g��髉)�l���Z!�0�r4�u�L�
��Nn�3�Ye3�?~��.��vÌi��kz�
�p�YvL���9�U*lI�-2`T|�P�z,������۠��g�Ac���>����x�m�{�~��L-���<�c�K6��h�!0B���L"l٪��*�Ei�.nR��h�������������I�x�К���:���q/Gq-��/)�q��Ї�+�B�.�[H��#�1лP
�Me��QV)�\��d�
�a��8��[9y�{:k��͘R��<g��yb���K�^U�H����Z����y<��.�P��{f�o^��s�~|���u/�~�F3n�\�=���N!$��\u�Y���� �T��+�<G N[̃��C;q{����y��l���Ak�4����&ų��o���#䠎Y!&��.�Wޝ�
����isM-Ƃ�*��nN��u�3��s�V�G/��6�"vR��1�A]z|��g�m�oȼ�9��:nyC��EL���@�U��iR]\�8ؼ�~ ���b�Ɨd�Sy��_=�;37��v�'=��=k�U%E��)�De�~�,DLRh3�
��f��A��=]C�*��a�Q���rz�p�{�Z�p
Tz��[z��!�mmE"�r�&���ɸ#�l����p�$������ɬ���,���G+���?��76����1F;Q��9Lނ�xl7��{���xzn�8f��VFf�����X���U:p�Q�A��Ȍ���4�_#�y!� x�Dܮv�Ǩ�whR�
g#�V!�<�Em����a���m�I�Y����a.����v��aZ� ��)�I���q�%-h;e��Fj?)��5���+.��M�vu_����Ҡ������̞���X�a�AiX��ݝ�T} UV�7�a�Za��&���z �߹C��vi�԰����k�9��'���.mq}íct�)���VG�9x��Q*q3�l�]��jL J��G;GZ�	��f�����e��O�,�y���xO�+O�hx�ژ.;�[q�*����#rF��2%jf^a[D�w׺4Nw�W����\��Eeaa����y�U�{)��}��z���貳y���xs,�^�µ�����u&�(a��"D�W��-/��)��	$DZ�"[�|��i�����la�R&���o��
��VRX!�ҡ,��~��JM�N� d�j�<ލ���2v`��6-gp���L�5�y_ի����kn�!��V�]�n#w�G�k�Ľ��4�X"��O��(�]b�2�#;=��ǎ�b�a޸��!R�`�RM9��F�R�z+�»'����>3�}�4s}��+��ă���Ԭnnj�����&2`f?��dՂ;��v��sg�V�����6�}������%">G�\u��@N�V���]ڷ�ۮ���&�ʿxT��������.���@��gE��~�Nk6�ۉ���xUڹ!�~�w�(#*=�(�7մIEM�yk�~�V�B�)���ֈ)<��/ﺇ��1T?�@7[�����|x��@K��;�'i�&�a�nM�
_k�SO��4抩)8*k����g�nyp�3�4��.��4��9����BT�ۼ7zD
���D!`,���3Em ��+\�q��w%�d�&�m���*�/� ��PO�� �`���Ѓk�!L��=0�8zGV,�G�n�a���a'���D���5��*�zC:�^-9S�l_�ȿU1g+-�-/��܄4�Ȧ��Q)�&�7��
m7���������L4�0-�P���ޭ����� <6��a�d�C��v�n{�C�P�
�=4��N3{�m�4�H?��	�{tz����;�Ba]�(��W|� �4*p�� u^��]�Z�׎�/��¹�����7Ą���XŰݠh����_�N�� �`���Q�.��>�x1eT={SA��������\�U:@;�k2�	��,셧�	3����l��k�'��y�<��YNt����{� ���jNjɿ{E���=�얫�ʲ�9�n������Z�e��k"#��tE	�\ݎ�L�� ?�3����dk.��2�ħ�&�R�u�u�й�M��(��ƿk�E���<_�Ќ,��۷+e;��N6f�����S�yl[�99z<?<~һ��9��kN�0�rXr��f&�26���hŎ\;o�7F����!�A�p�O�I֧��=���6H�T̆���� ���:٬pכp~���o�RD�6�9�K���#$b���j}8q��Q��E�7��f{IE���*m�t��ǘ�V.��d��y���E�J����
����	}��O�&[/_v:��F�����n���)�&B�E�s��7��Y���:�`;�K/@�E3f�j8�8,��"�[\3�F�@=ke��@8����8v��d���"ȜOJb�Q���ٽ�N>]rA%:_t�����fx���$``�}a&B秘�	�A�����L�"�J)nYE���ws��tr9���o�H��Z����m��*b��ښz ��V���������L���Jr<;�ħvZ��S3�h��cox2���f����P��8[���HpD�9Ӿ�(�{�ҵ�=�&��Ēۄ���gq�s�Ө�|I�K�&G��$�����.Ѫ��ݟC� �A/Uu��fp}J���g��[���"c�%�baq[��w+���#��I���x����7��ª6�s���ޕ�Dě�c�J�*��n*�d8��>�p'�L�y��������F��Q�M	���
od�BNLֵp?j��Dy�����hjWt�̀�&���m�HLs����#MB� Q"��BL� 9"e\v���ջ�Ν�#�7M����=�V���qS¤��Й׶�����.۾��s��j�+�o��Ć����6vN�G��l�?���u|.k��PRQ��M@��Ae}��������E{q��K
����ƣ��&&�JJF?�z_Ś��
��߄չH������Ø��szF|^@�l�j��u�����yV�-ٿ"zs�Υw�C���JM�O��u�<da�r�}mj^P*z,���$��GQbM��r��76
��+�k���Cע9�拋G���r���&�>�b-t9��!�f' '�G����7z��:�V���jE�/!����=�5]�bc�3��l�VkeUpM��O-���+,[��$R2����R��v���*�[���ۯ
X���
�.bߍ�z�￧s�+"2�~�(❷�W����z��o��T�d�P���V8���\�V�N�$�n��8-J>Rn�i֮U_��)~7���cT����C�3
�0���X@ c�s���䆟b� �o;���h�s~�J�>�[x�e�La�i�c L]E�}�����{G5�u�Q��Y�-�H�#]:�j�)UzWB�	���M:��� ��J��[h�J�p���~�;�;�=㌓12�h��,Ϝ�y�z����MZ����,0�񠜖G.`ʡ鹽������}�g��g��"�LQ�
5-[��aF�Z��vp��q�uxz����;�B�2��5k٥͟2�o'�!����8D~n+�P'݀��5���c����_���O�N<6�35�hv21z鉔���ؒ��mN~���f�Q���!�4���vת7���c�O�!�ͽK
���ό���6�.k�(&IHxm����M���-(��S6&�����ՠ�v� ����,4I��
��0���qЭr[0���s�#F���q��ژE��L��Q4Pa�����b��g�&�>��[����,!�����'*��n@�K"�#�{�\�#E�Q�=l�B\���Q�U�ςK������C�lj*�L�.yk�����M�	����"ǻ�EK���A"7E3�bKNInmP��=dٓ�O�1����Ј$��Y�Q�l�	���[)$M�/����Z��g��vlzrV=͙J�i��x�,>��Q�F��E�|cRq�M�D����}d������X��o��Z����2��lR�b�gZ��b:�B�yD�������"�L\�b3�m���<dǺ|g�0�$�E5��2�&�S�?WT�=n�8BȖ���/	���XW�M�5�LQ�j������K��p�^�oI(a>��G$���D�7��Ǒ�V��4�4�	�H5f녌��:%�����	̹�Ug�6�A��y�h���򥫶�\F���8��ښ�Ι�/ݣeӆ��@ꂶ&�,�4��v�=�c��s�؋�Tvםb	�}�S�2IB¡�o�O��2*mQ���3ffajT�"�{��)�	�8��̕�꧉z'/����	�b���t���t���L]|*��d����-e��˖� Ex�&ս���nؿ#���x��BC޾O�k	��ur�����l�x3Y� �Q+lbiawD���`��(�T_�M�s!U���͘/4���Y��fh�Q�J�&X����~�0/�?X�����O?������y��	� 8���ʽJ���1�ܬ9��G(�XZ���I_P�7%�*jjr��l-?�7�����W�O�Lѭ'��k��YaL;	�����ڮd���O����h�0����Asa9������?�2�����w��":Q�b�Fb���G��tT]�/xl�!�����s��O*�Fx�����~�c͖���)����Cc���k/щl�H$~��ô����ҋR�Ts|>�N�_@��ii:�=�J��/Gس;�o,��z�+I�SL ����c3�.�t�]�k�>KE�
!BCo�Ѡ����	*����%I9�?Fi+]uǕ�.
���qf�������ڸK�� 5B���u�Ĥ�	ӇqO�.��퇊<W�'�|�^!��g��75mthB�:�����਼����#��B�˵k�W�ʖ��F�Ћ�R�F��[N�����,�
��Yh$,�s�^�P���3��:7�zW?�싡r.�i;������:�|�;�h��FPk���A����|�;�����2;�u�Ȱ����C����ܳ"t�ֺ����C�:)�m(ܼ6��9��Ĵǧz���<>fl������:$U�I��Vb��4g���%���p3S4_;�8PN��X���g_&�6S��lc��X���C{{�{�}	�E�x���Y-)�4|�'��0S`�
��K���xH�<�%Or��s8�� 7�[��tX��bT`1"������-�l��*Vܹ�DZ�=z<Gu��(s�Z�4{�甯iG#��|#a��8ޣțGE8���9��L>�g h�����?EG]���7�_f;�L���u��pN��oG�������Z�o��B�EW�fT�nj�K+��vJ�:��/#3E����)	���	�&��o�����<WL�7��r�t���M�=�(m�W���������kU�`�ѕ{m�Y?�[y�Ŝ�Z�[}��F������V#��ֺƈ�z��gOY�`6����BPnO�L��3�^���Dp)V�93vY�}�>.����@@���jȭ�-�hV�A�2,�Ň��=���O�����=d��7�pD49�5��~�S����������斳]#�b��\KNV�u��HC,g����T��6U#]�%*�ʹ��^��!�D'*qg�NТ$�D����z/�!�c���[�OzD�
���^-ұ^��w��,�v(�@;|�yY`kՉ�������6fX�v��$�λuI�.;=mނ�9T�ѣЖb�D��=�[Ȃ�6g����q>Ŋ�(ӫ
�hf�ց��DQ�Ѱ�{{o<��9���=���f~*n�D�C}������h���9NI�����$�##qUȄ��;�)q���h�A`|�/]���V�� �+"�Z�1»g<�7+0�u*1�7�����<�ˍ��ա{�=Eb�[�����Ң���.O���l� �*L���:������V���"3�+�~t�k4�#23s���� ��_��������耒� ��c��`W�,�H8��2�x��!st4�+So�+~�<��#�py](�����(K�5��NK&)�.��9l�Q9�8��O�73#�T�^���*2�*+w�Y�Jt^<+�xF���kdx\�wn��c�u��{C7���cV����)�!I���XE�|Q
<[����EKs*���������Th��U���q��NB"s��2��P�퐽�Z7Dn��	�v?���*�~���X�^��R�7�"��A:P2`�=w�?cwy)�A�PMucfT������)'�gN��\�ϝx���m��ls�u�H�u^�`L�V3�'���r�)�CF�?x>�Jl�"�z���Ō>�4��ZWc܏4,%f�������~���ѷǗ֯!�L7`�z�#�u���o�!�$�?ʴ@��(_��y�\+����L�#�V�oGC�/ߝ�$%P�����ld:m�ҊeF�:[W��J�I[cC�;!߿�d���7��z�%#4�u��s]n�zS�)%�����!��d��r��Us�@&_�EO��~l J�a�pd.��:F���y������&�.��	(���i#��Ԝ�$n�����=����[�����P�1�L�PX,u�O�V2�H�%��.+o�1����\�B�Zw��Jt����L��B��F���ƚQ�aX*�d���_k�M\�M>Tڴ�"4��:�mP�c�����_.]�\eQ������A�ts�&�o�d;jLga9	�\��>�b9��Lֶ4�Jg'O�W�<P���8(S�K��d�H;vʡJ1�� �yؤ=�r�˕$�Ŀ����0�G��>VW5*��ۗIB�r㸱�K97�?�&:����^ Ħ�h��o����7�E۳Lk���͎��#� ��T�W�[y�y}�j[|$�4���;m[�����N�)��b��"��*_�6W�qf��&�N�<�^������; ��XND�@��tK�����Eq���?Ǥj�Ǐdx���N��a����kU�.f&���:�Y��.�6~@���PF7�/'M��G?iX�s��%h���*�n#�(19��wX�B,�0����J쭂��AM�[�i��Bȝ�99�0���)�CGQ�h����G�Sj�T̼Q�0ÉW��w]���Ff��F^E���~�R�V+σ�G���葃ھ��|@DW����Ն�k���/銶���,�´��Ŝ��/Id?4R'��pn��o�]����s[&&c����&t�����T��sv,)�:�:ĳ�q�'�[�'���4U�����0��g-����sҾdf�[AG���g��]�̍{�ڦ����c9-�M��\]jrM�3�z`=p����_z�8��B�ɳ�h�+�\���G@��+X8ZM&�����:@��<��(�m�x�_�������$vG�:X��$�y(�4���2%����]�j6QȺ�c����9�3'%��t���@s���jF�ӵ���o�iB}�F�����u�U����j�md08#	#�Ԍ����t��%gE�D�rx�9i%�(��[՟*=���V��n�}�\��5GB�:����J0SG����gp���!ƀ�'��
�����A��yc��ŋ���DI��$v���4�c:�Sԫ�}}�W���a��0�������.tO��V���pn!�w�κ�FQ��"6��$�KY!�ysl����_���r1^�[K4M�0�6�-������x����c/�Y�ùɬ�6����e2R'������9mJ�ݷ�QTMN�=����}�ﴷ�Ѩymڂ�_�=[�Xx������w��y�"%?��b�T�P9�I�q@J�V�uGJ���X���^����yOz1I��>.,�=l��:F��K/�s���7�m�#"�����1��ߗb_ M<�L_V�G��*�ε�̡��}���ɐ���W�u���n`�F�/?�,�1�3����13���511�����ǐ8^�J�([O���ٷ埵�5��t8fe~%�j���!i�S~Oy��]g��W�V�(�d*��S��$�(w����m�x�5�P�a�O
��J��k���R�8XnX��6$hpD�m%+P��T�u������2c�4L�zVV�c���8\}�����w!�UO�кy�RjVê#��4��b� �2L�C'��tZoU������śƻ���Ֆ9����E��ME�w�d��S��K��#e,c��ɷ|W�Я�=�W�?,j.n�o!�@.��%.�{����!���͐�x5�:V�W��[%nCŅ��:�q>sQ���Z�8�y|]�x]e��=�m:�)I��:�n������RTj�v��m��F�^�����"�9���h�/�M�3�jR���4a�lw��8kt�5�86C��#���[��V|��?�2�ݜ��P���)�mЋ��S��Nq�|��r�GnYn�2�W��i��U����$F��#�y�i�OOO�d���[k�����k��fq�nf3t��S��H�B0#�|��	�0�~�F�8��N�>y&�̓�*���r$k��F)���
H����y����u�o�\�Մb�Q�l����ߘ��������V������� $Fg�<\�-m�| �Q`KnۙG�ai�)�?�u�z�,eec��zc�"��D.zUs@�5��h�5���c�mq]%��P��|��d�#�:3N�9�\��g�J#G���u���@G�x�B4�as�bV�����
ɬ�Q/��Ԣ_/�[�%���ɖ����2�zJ �j����\u���\��Ź��i�+q%�:�%�Y���?�:̜q%o|o�ƺik~&3�K�,��|��㬗niW�躱�g�����X�T��w��T3���� (�:��j���������p�歕%�)���x����EU�؀oߍ�r+���}~��|���58�&��*�#�r��ߐ\(
96�7Z�9Z��3s�� �`5��[��+��k���n�ےf�G�Ȟ��ėS�
���DUFE�NɌk��^�^x���?�;�H �U"pխ|������,�J���7J�5˰����;0ڟ�;=�"I�W�# �;�ż�bۂc�HCVO����y�z�����y�5N�H�!j2��o�^��(�-3�M$��ғ�����b��+�v�h��n����u��֣���N�|�2m�t�g�Q`e���]�b����H�g�Z9Y����!Y��XֹM�o�iЭ�TP펯�_l`��
��l�l+B��q~���ىOR�mH3�RZW�WU�W���x�r+���+�#�Ϭ�nq�}���P�rUx���}�Z��Y��Ӿ���*��;�@�1�繢x&]��uO7��7���fu����"�����l��Ap��9ށP��X��+|��n��40;a�ף!�=~������/Q_1_���B���5ҋl����}��6׵�oJ��)w��l���g��Ew�(���Q�D~������T�y��5,����C�cI�;E��]C|����sf�'���Y��3��0�y�(1��HN��s/���.٨���S�w�P�Gn�\��yge�;�!Z�=C�$q������X��o�M�����GXֆ����GY�󜄃P�Bq�*N�D�sؐ�_Z�~��GQt�Ⱥ��o	r�0�:�
�qr{;G�j*o�Fd��m��_��]v6�0c(�{�.�bضV�b�ڬ6�9��~3��m��.p`��������W��9�y=ƚ�E�_O��6��+h�^�`�8�c��%���k���uc9X1��a���5K�΁r��`�����hϗ�6�_=!�1y�G֊Y��a� PW߅)g��~�_����e]��7q>��=Օ%���v�`kQ�Z�1-���-�}VQ�kn}Ͳ�)/�e-T�̈�U��p� Wd\l)���	�Q=�j�;�p��1݌�>�Ǖ�~��v��w�{�����y��q�9�6u�21���+\˼W�EW���{Q?&�q�ZY� C���zp����Ĥ؈d�O�yψF�u�g�U�=�a-A���#�ޢw���q4�j]�"��Z�����zm!^�U�V�e�н���X�7LI5v!g�yl�eԙ��ۂ�2��75�rl{�q�Y^�l�;��A����x*���*4����.�}�^��,::�nw�ӰԃU淪"���J?rUrR�Z�A�<�� 1��Dα�D}4	�(e��L��z�u����cs�0��-.�lDu��:��w�W
��Z4��T�� U�k����xs''Pf������gX�$��]D�<�K���Vl�P_,@�mK���\�0Z��#{ �Cd�9l���S�g>�e�9�X�C�Y�6@��nYd�"�2��NO9R��o�쬿f��%�^A�sت.�A��/��m�MU�uu/=�y��tku��PRPi%YJY\���_�ȷ�![Ȥ/6�8}Je8T�@o�`�*�'�q����|3"�j�-`���Z�j�]�2Qw��nǲ���+ Zv�g���@� �ur ��IX���C�F��x��M2qT?���`��S�F�!��r�����jҾ)Z�뜏+�kv'�D�!Fٗ�ڗ#xM q��%ܐVQ��O%����K05h揊a��PQ��߉�T��{͸��NL{�MM$K��pZ�zc�Fϖ��@�uYATŵ���>H�%:�Ȯ��ch�_�0I`���յ�I��mF]�q�!�d���R��iM�.J����(5����{�m�E%�{W�����w�L �E��vs��N�ߦ��l{q��o`9kӰ�eN�<G�_����G���� ���Gc�aIq�S���UaSP��q�h���L�
��Q[k� �?,)/�������&K��t �� ��y"�|��@_B��uu{T���4H0�i�9,�<W��w�_������� �9[\��bDt��o ��_j7��{�*�1d��X��oXx/�k�t��'6z���s���ck�[����@��,��a�J�AMTFw'ݬ�O�'���9k5�c�*�05�|��H(U�	!�,�o�ھ���_���E�
�+Nk?�p���b��HT�M���*��~ -_@�U�A0���O?�mc���ڐ����:�0���A���#}FW ��3B��6���refAR�:]��L�4N�{�m��NՔ�S���=������x��dz�!n�����5tg}�!���b/Xf��*�l�]�!b�����s�كq����\ܒ7���GB�5��x�Q���S_������-/���@|P�f4*�m
��)��j�k7��h� ����Nͩ/wR+	�F�a����~M�_�V���� �>�,-��l�Sk���;��HY��ܳxڃ��]"�����+�mv_���U�T"�� ��y.֚zh�	���z�mzj�a ����&����Y�k�xQA������Y�Y����A�W�\a����� ��dr�4���zU�bNe�˧�M�>�+�`�vzU�PJ� ���z��pl���& �y�Cj�BZ}^���:s q�:��Ζ��蛄�h�q�RЗ^�	G�i�Olr�Ag��i�}��@u����V��7�� �+�so��7c�Ά����Ɩ[7�sFs�󹦭�-7eH����K�;u�i���Ǯ5��/\�����m=�#�A��@�L�[���A?9H~���J�v����)�*5�3������*�=f�qEbq�t����N�p+KH������:»�i��������3�6��Ⱦ7{V�?���B"���Mt2[A&��J�Qm�_z���EY�e7٤��#���\B��:&o���-Ӟ�K0��4��	����|a����n�t��=�܀�
|��^��9���Z��Ux[�^Er����m���I�.�����A^ ܎B浟\Z�&���a���EO?���z\Q@��t�/+:�'�i�cQOa[;�ޟU�g�r:	���@������>�!�ϔ�����҄�q�ޙNR,�eVDV��~�|_�Z��ԲUR�z�v���M�uD�&h0Q�z��u��h����<t� ���	�|9<]u�;]ޠ��e)�d@_-sr��w����T1�t�V����e"=��/�U7�{!�% �d����y��P�A��?��.�ʟO4����ȳ�v��O\ʭJ�b�$Y�b��#�޸�`�+��]|�@O:Yؽ{+���x%�b�ͯ�
,��Q;�Y6�?Ы+ˬ'+�Va�wԋB��O�����r��(C��>���&hJ�ben��'�s?~�`���K�l�mvO�vz����]"�[����'���>y ������p� �y�B�����`�G�!zUJ�o�i��$�Mܣ��`���poOF���M��Vc��4RCrC�5�Cr��4�8����8?�ǘiվߵ��*����?.���:�`��F|C�wo�>|�(��ߺ�S���b��U>Q������5��-���;��3LI��;)��7k��v�R$��dM��"j���f��VT�V��Sy��lH��ҽ��S��oiI+��p��rE5�+�XN��Z�������x~IOS�l����J�tI�鲽�~�Go�&) �W�zm�^�<ր�����Q��-�E~spZU�@T���Ȏ!3�}�Jc�H*�<o��T�2+4(�����aJ�������&��V��:C�+�����U���oA��� ���e�.#���g�zf6��U}_�0�3$p`���{�st�`�؋�?0w����a����-�ϏO�jd�E���|�����]�lX�Չ�Il��G�ɗh+I@P�-q��9��NTO�a�Ǉ��O/���Ԉ82����霵GZ���A�`[��N�?��e6N�T���)Q:�r��C/!��bN+햆���g��h��0��[��:���S���/~M
��H;��}1vw�sv�:���ry����%���2����^��u�|0¨�nS��J}�#��<�
>�}����q΄h�@�GdP%x/J����{��b�[�9��~�b�FPr<���-��|#O�㓔<���y�`n�}�O-~3��NL�Q��Y�^�( W[#�t�A뾆t'�����kQ��Ne������w��#-� ;ˡ����l��������)Ub�KH=�a�-7�jѠ0���VP}��L�ʉ��7�0P7Zi��g�8���p�����E#��1������w��qC���Y�Lw�|d���B`+���t�X��vO�j���w�����EL�J*1�
�C�3\o�8�qX�V��*��(1��D�f����(�g4�B����I�����G��T(5��.A��/�yK1�l7��X�o��`F#1+�岺y2:zb�ͭ�iC
]�'�����8��솧��k^f�b�_���/��vm���7>>�:Lg@�L'����C�dkF������7���e�>�'�3�"
��X���A<5�&�����d�� ��?�=P���"��Ff�?jw�I1���ub���� ���n��Y��ҍ�H�4�x1O���]�Y�N���D��~�\�<|j�ܿH�ߓD 0���~��y-z�G�_���O��SW�R�^���m����'�>�ˈ^�9:�k����ubQ��w���۩f�)�R��p�[߀��t	�hNY��?�{��AXn�5��,��o��
QJM'�R.��Q�<a���}�X����7�s��>L�����~����[nO�0���w��m��U��E�//b�I7-S�HRˋ�-�-�p�'Ol,l���������7�j�?Z8.���*?+tb�O�?ƪ�(��UՉ*��z"kn�(�-X��z���J�b�����`9#�r�bW�H-O�{~�y���4��ZC����*Wdåu�z�LЅ�6068�J�g(�.�cz�k��Bxcrq�B�����^�}hP�N�K�����G�9J\��Xa׵�n��|}�!����W���!_s�Q��<���1�5e����&^�A2��J�� �K[�8�hl���1�0�W��	��F�j�p3�V� �k�0��n�D� ��8���<�Q�uG;�H���B�wm���P��w]��箿���kV�wkӊi���}�����mp�V����_/=�17���i���et��\�w2�{�XXίy�d���H���\[�R��wɼ��{+�<֖����\jj�{}�k�c�*6��=�Q���!>�@�Q�L%�`>�3�ݥb݋��d��y�ӟ��A���ug��P�wSʀ|��y�sN�	����i�0��Еc�u�(�j��k��|�\�ht����T{8(m�Ԕ�p���v�Z҂@��������G�h�s�Ӣ���Ǐss���3�������Y�܌sv�d���S�q.�a���TTjn'�V���)U*���a������4b�R�%5��;�up����w����z�"$kl��`o�-q�Z�Be�_k��m�<V*�ZW��0u7�����P@9�T<�Q��v��7�ǘ̕��7,G/}��gvWj�>Xޙ�5�3��7�{zp��t���罿77�||�|����ء�0��F#���E��5
ލ�2�ܣ��_1{_��qrQ���S_Ť,�_��ݟ�j2�(�o0���鬠�~w}�a<%Zo��s�qk���.��==������4�E�pr�|"]I������C��� �+��Y�j|9��
�L���^�}���O(*qP���Y}+suR�R���G��Ix���,t�o��C[�����0���W����Q������yY;n�9��h��� ��DG������}, З{���$Ew��8�R@��=$�
)�������IGO��I�߶:�\n{�{A���^��bt]R��$:9^��R�ҵd6��x�Ƌ�Ea����n6\�~m;a� �0����=q��)fp!�r�ӥ�_��q|�r>oa��MGl%��ٹ�@�j��J��!�}P~,[X�D��5�-e�dY��Yz�h��J$��n�o#.���A���DU��8Txy/ 5� ����n2�lZk�!���yC�}]G����N���͔�y�ڎō�T��/�c��3\�"
��V�=Y �:c�#x��������؎eoG�ݙ������_����zme��Ѵ�Ԩ����d�����@Gg@8�:N��ᶝ�0�w���E���}!r�%� ?�L`�`��_���v����:Y}w/c��@��tB�L<���	��)9۹�U�|�N�+s0���24b�:ܭ;tJn����=(��y��Eq��l6�N�yYyE}S5�l�c�LKO����{U#�ijU-*0q��&��L	�g���(�,� �	J����ӌ��,C��WM;��
��?�%�M���o��P���F$��-ぽ�վ5�����	ST�x���'x��J������c�݃�)���
�ϗ���)ɴ�u_9z��-�]�М\�+�E���Q0���nB3[�4����`�������f�����kv^q�T߲g��>���2�����j�=���Q���`~-�2�؄�=�n�11N��
7,k6?qn�/"��N�3�����p��`�K4�^qE�q�v2�68�9���t0�l`�����x�쓼�M�g�rF�4����� q2_2dPF��w�~�ʬ܏��/k1�=q�|����������8W�j�K�U�h��a`ŋA���y���S����x�r㶗���O[��8��}�_�ǿ��df�7M��qQ����
��&����"*���@u�H�(�O�XGu�����C=��p�}�V^ۭ �e.��4tI5�CXl]����f�/kq���{-n�*7��L{(i�J'�L7�	�����/u��C�y�#�ŭ>|l��n�Y�ڥ�w��2�'1WK�4Al79�i�Ѐv�zF���?�ɵVx���4x�y���)y?����y�X�.�c7�o���;9a�[Ub�~���Ep��Z0��K�D6cP�J�V� )eb7Kr���\�˾��_�?5K�&���3���#[���b'���#���&���y�&>���u`z�IJ�Z�����9Dc��v�(V���C�0�^�닌��%���TA�O����H(o�#��=��\��% &uW� �v�Ϳ�A��{()�|A�7��u2�ݾ���Q�9F<����jxȏ���_q��|�·�����΀:�l,�5�ޮ�.�_MZ:!#?�ċ\���Də���qC�d���d��bH�J�^�1������bO�#�h�:��I��G�sͺCC�4G7�=aHk��+'����c�p]�!�aM����.��-%�j��^9$5E�zY_��q�݅7kx�ᦫ�I�Ut�T�G����&����3��V�c9�O��U�*��.�/�ŷ:�?�w �ц�b˸�3�A�\2�/#N����Kf�u�<Y�1g�O��f���,HE�����+&_8��m7ڵ뫊k1�Pz����ĬKzl��MN�/qjI��{��6���s5C�(XfZ����~Ҭkra���['�iN�����ŏ�kza�&�; �E��Jς�?��V�!zX��o��)��|��k39G��lY���b�[�&N[[�^�ʈ�����x���[2������d;�.Ӑ�ӭ������i�����Q*%�жt��G���2
��}U�k��΍�T��r�k�]�by�ɞq�>f�H�~���W܉���O@�R蹨%2M>��41H�Ө=Fb>L��x$R��Bf*��V�������9�Wq��$�5����DDPF2��$�����P-�3�71e�P�^!�H�����ݣ����o�mmgdT�Ϲ�t�E`� �&m���H���@[$�л�K&���5����_�g�o����S��6����\1���8��⑲l8X��k����4J��8�h��@g�� �V���&M1�hqRPZ<Vv�)w7��+��ig��sҴ��'
��0�H����C����~���D�ϡW^�1W� 4�B��k$��,��U�q�3?9J�:�>��υs�|���?��HN�
5��f���B���*�!c�("����C;	aJ��zZ���l�3�(lCcgk��캛
�	��+Z�.�K��3���SUWě!��pQ���s	*婝�_@rЙ����OC�?vĄ S>�<���kx&b��P�ƥ���u�`}�?��Q�b���	K��Q����/)�_�� �.u��2x��뵲}�Q���,aq���y)��C@�fy_��o�?Y��1��ɄTq�q� L����(�\^}��������s�k����Y�;�\�ѻ�629�Y�3L�?�l;m���ͽ1�;pE��Q���E��-[������c��=���v0{ZU,#���rP���ҟzu�ֿxM�+�p�}��?�R�}�#6�l$H>��;��}�\;��O�&�[Ȭ�9̸I��DÅ��>v���=�		P6F�E�'	�7���A�yǵ�e�]�,]h8��c��լ=[�q������傳U7�'��-�>�h�=]�RۺLү�Qh���n��J �����������l�(sIT;����N�q�q>}��>��7H@���{�%���"s��$�{	�w0�+~�p۹�� �MT���y�)Z�Iۚ�z44�������%J�u��Q>�j�y�+4cN�P��L�I^3�,�ad���L��z:k'�Ή[;
ۧ/�aGf�eϡ�A�]�k��@�Z�!c"�o}<\��bI����+�b|p�Ch�ұ
��v��J��AZb����"���#(}mE�z��r�6���[[wM��`��@�2�)%������������]��S�bL�P�X�M	\���̅9z�q7���lܠ�d6�'������q��������2O."�]Iv�ÖJp�fc^�5,�`����������A�R�zE/j��S�X*�:82n�߰�����ĺ��¶�ǩbQMP
�QW>L-��W���o:�OD-`<e��i�}[Υ� �\vb�k��enk$Z+�y$��R�FJ�WW�ǻ�=�C����q6'v���������f$�䉯����iU���u�齫���O�W�������l"u�4�߈ �ڈg��$�I���;�+����(q/J1B9��,[Sk���*���/Z�T�	 "�@Cy��1��g܍S!@�˾M<�#��V�N�0���K珕��͝���Z?4�h�������=h�:����B�<��;gQ�HO#l8B�h���f��3��GVf��4P]~�m�4��a�o��[!�5,�;�ʐ�yS�Q�5��H�<�}�!RC@�4#Eԓ�l��jab�u�����a�+]�}QD��ڝ� N����u��3��:L>�����X��hH�7&��{�=	��{�z���k�r6�l{]eN��w'g�r� �����DlRLT����7ʫ�+�K� �����N�?��5�3]�{>��z>(��(�(����k(�_gf'`e�ei�	�V��I�N������ބ�@�����ce���eN�#��~^��k�P,��}���� �ǽ���K'�"Y��u&
Cd}�w�iP�ڕn�)졟�5D��tׁ�:��0��|lQ���\.Ɂ��q�WX�h��	�+~E�?�XR�.{�g-V+K��q�QL��`����ꛤ=�A)d$� qȡ��" 0=��?��������m0��xSGR�$z�����[�Lp�kw���ӗ:ݡ���n;�;G����K����N��%��~#����v���91��x�5+���7�^�s�e�<^�M���%�$Nx�g����<*��~�^EAtep���($>�Ȁ)��T)��\��a+��!��^/�W`j�1���g!?z�%����^Wn5�x�L�|L2�����G���n���ݒ�yY�Ha�R��q��u<��a̕�5#�~'�6�_u��t_ԯB'[�Jf���h4>6`�?�x-�g��w�Z��Ш6��
������f��vIsH�V�N�F#�ɺ#Ėk_jX��/0����z����f4���g|�!��g+�'-�a�vE��3�T��c�J�+F������RPpÎ�ǆzk�':���˿����GQ��-t=i�����.?�8����&R�a"�*�e�_�s{��w�(�]E�[_ߞ�g����5�v>l�-z�[�cޠ��o(��˧Y!������(�6=гX1�����x�0\"�Sg[k,����CRM���������I����(4`gË�n�����5]�1�V�����gJ2Q�=��#��]��K�^�`�  Ɵ�N�n������Dؖ��D�Z��;�,��kA�gY���iŘv��;Ǧ���s}�V���nw���Ѝx�y����Z�h�c��o�M� 1YrU8�/��E>9�(��s󝸹=n�hNh`�uT�K��e�Z�Ybc�˪�C�;��8��9&T3��+g���!<T�6�j���JN�	Hx=�#����o �n'	7Q̚ݱT���$-w��^����mg��K��OT��%k8��aJst�5ϑ�ԲZά@q����Y�2?U��[�8���4 ��z�3�p��Ah䡞�{
;4
ޯ��*C��k���4����c�]Z��X_E����;pE㵡������:�������?�#�ѯ�J��w:��#C������#E���42�(p`�����j5���^��B�vxw,!�|4.f��R�޿�o�&���O�&[��3ʢh˩S��@��m����a��~^��fD��գ��rݭ������/*���OR��+����2Pmb��"��"B~H{��bm$���h���fJش�Z�RL&���p��6�S�?)^n?9��Vz�n�hWdZz�- &�e��2s�-B�TDa�ReYA�x���B6�|%��������YE��jk��O�����$�`~\��4�b���`	�R�A��ڕV�}�77�,�k��`R�Ϯ�q�a��0�%(d_�w��s�1��`�$E����qnt��I���Kq��u�#Զд��Ud�����zK\�}�"�Y3V�hOE����.��̆�+4������=n�m�zr��$y�"�D�a�9w������;i~� t�����ΏM�u�_jEu���5��-��,�F���eSU�$���[	Eiׄ���-GkU�{`�v��B%Q5�Yu
d�(����B[[����w��I#T��b��C-,K�00;��&��:��R}��[���#�v$ �,���`ђ�E�n�jԲ�=lY�ٸ/vv�6
�a��cg��r�ֻ��O�FE�K�~]��,oWK/x����6�:�(���͈�m#]�2cj�^����.Zo�pAੌ�)2F�mÍ�-x�� �vi/�l縛l/����C�W@5��������R�!!*�J
#��H�(!��J���Q" �G�!���L��ϣ���9���x��]�~v��?�������\��Tj鈨�g���1�s�4!�$��Tɪ1z�.��NL2���N�*=o�`��N^����W��z�\����k��uꜩ�����[�nk����M�d�p��7��@��"6�PI����N{|�u��\��	NG!ӆ4�߇4���y:eb��q���r�8fڻ�%��|�x`@cK��n����KX�7M�T�AD�,��P��	�0�N��Lq�`
0�$�Δ�gԹ��y���Ip0&��b������y=麤�T�>ǙB�;��5wd�׺�b����)7�˶ۛ�m��	ƣ�����^t�m�`L� �v<ꭺ�s��}]���3�����bD:��[�S]�ܵO�)Hѵ������{B��H����B��}#]�fiB/�%'K��}��D���M�s�����ࣳ�L�l=��� �=���(�:7�Z�����>#}OPdx��.GO�&��"���W/@'\����4'` �b��Jms#S�
[i���4��HM׾�K�:�<%�YYƶ��K��ii��<iPa�a7W3(�@�ƴ��0�s�h��"��5ϜA��8͡=66Ei�w��Xq&<~,m��G4�9��cV`�)[��ޜ&�3��Ѡ��BQ�d͡�|n�b�B5,��[F���ш���eە�yh'-���}(�4f=l{��!�R�[m��a��ic��J-㽕�`��R�f^�31~d|�)��ו�"Phc��}�����Փԭ�JΕp�7v�8ڻخ�t��5Ui�=�i<<��ڹK3^��l��� �v �Zvf1��5��y��T��&h�?����FY�EͫVc�S��ce����M�݉jme�%�q��^o6�o�,0�B��M*��i����o�yzw�`�̊�����B�]�gV	��D�g;�w	NL�'�V>�_bj��xa�����jB%D��&�����V�@'`��F]WHtLӓD����{��/�=\I�]��_��X��i�Eii[*��m͍����o%r뱧�R�'W��|n��d�A���J��&�>��-e���hr�=�[g\=��!Ot�њ@���D.[+���

�=�A��|�������J��AQp5+]�{�l�����c)�h��(9|�tY�J	\fڍ��C�p;�.6�Ą�?�fK`���5�3���{FOG'�:�hm�K�,))t�k���u�s�=H���ۄ�#/|בn4��۶6����8��V�^����L%e��o�T���Kno1,�����6�uE�g6�w,3�\b麌�k3�&��{����m�Z��F�͑���ϥ����S�2�˚P>>��&f�8I���I���B�)��k��f}��Y>#*
��e��a�;�{4xyEƝ��}�C���zQ�y�4H����aa^�j��Z:#����U$���N��{��n�YFD9�W;_�v��ڟ8u�U�f\E-�?/&r�-�z�~B�[~����AW�VZ?,-v=@�õ����s����{0���Qf.�;��t�k��`h��v��<��Q���*�>�,��G$�U����f�>y
�m��H��S�z����<e����u�
�� ��5�C�tf0��z�IX����g?=�bX�39@��zl.�+f�x���$gp._i�iUrɀ�`�2u�'�1�	��H�A�>�>q k�xw��?\�^�΍�����D���i�5T:��#+���E��,�z��o�7�Э�47��+=�Y���N�.�ۧ#�U�^�U���VL�*�K>J�g.�%���Bġ�#���٭����A�ū��D��v{8�Ҹ��r;�zPjmP�7DL��rKtV�_#߂g#sl��C� T��n��d�����F�S�$�A�	�fܢ�-��p�uZe�]�{�k���Y����z@�X��鳣�%�)!?�3\�dBǩ�#��uX&*$L绰��fG^L��)>�|�i_�
�1���h��T���I���b�ݶ�
�
J,�	Qf���}mX6��U����6i���̢X#ޞ6�m"M��eI�?��%8�M��O>�s�?�����,䲴�(�����|�m���o�
+��#d�elg�+���O�ܥ�
R�_l�SŌ�J\=�BYgF�q���p��������:�/����m;E���([l���$se��� ���xN��)O�R�SO�"���2u�;7d= �>*/�N�5dKܽ7�٣ڗ�+"k�}F���9�c������T|_����E���[hH�iAd���YT�
���-�<�V��cޅ�aߚ��P���{g������Ω��y;Z������A;FtJ�����M��CQ@j��(A��ׇ�e��Z���]bhpX����>[@�ؠ�E**�6^g�lĵJ	��5B	�.�o�\�Y�n)y����a���\t߆&��pjx�ﾰ)�ҹ����<�:˙��J�ܨVu>u� a?T��kk\&1����
��姑g����]_�@H�SlGtun��h��9�5F[����c�@{V�g�%��r�����=�O�{ڲ�!���MǙ�u���E��5�3:�]Z�5H�$ҏtҟ�r5kO[6�tKuK�:\4Kj\�ԩ�.����C�.�:ń	ϧ2z�fAM���E^�.�(��O�}8�9�������S�L�2(�#ص���O��s���Z�AJ\3vI�)2��H�2�sPb�/dB`��9UX�s��O�n�N_����E����dw�w�N4��ҹ�4�R���:�H�����e.�3�k�vԇ��ڱ?L�Z�@jp�F�0�A94��U�V�"`S��5T�\D���:-�08���f�#S���~K���#���u��o�,硢�V1�o�4iL X�Ta��}u�r�a̡F�کZ�J��a�γ��I d�И��o\gLl�����9揎�t~�Gn�>Ѡ5�>��Jl����2���s�B�if�'�W�$��*s⧂B�P<�$HfWT|�u��%�Exٔ�|���C֑_/���5G����:	5� ��L���9�䤎#���?rV!4� ��v��GP�F�Y�H����mC'xl��W_4��o����X���X���F�
/Y�}���
8��7_��W��G%��}h��D7�^�\B�'�\A��W|ۯe������,�y���"�њ썝ȇ���[,r}�Ӷ�D/e(��A�U���c�;W/�[m�<�G9��(���6�t�OR�h����߆
�7ذM0IxΩ�Q줸]�z���X�.����(�c�Aw�iD��'�������V�%��s,��r��U�*&�3u���iZ���p��֋Mw/,��j�}��e�e%��C5=�c+N*;��&L�WU��]~�Y�R�ι���۞�귋Q�)C'��L��!j�N<��������nG��A���n/�����"ڢ�F-��ٻ���.U�k�;�4�'��p����ю9�N>�A�{���R)��v����TI�?�2$�i�)~��7�=4 �9�w���#I�-o�����j�ޙ1��hE[�xaUTm��i����T�Z.��.�*[�!�.�O��Дs��Sk;����{�
�?j;^܆�nj�=�&�ǉI������695����� z"&٨��
��0u��dB�t]I�khw8����G��Q�wMK\�l8&؂ �5V�47�3��.3#Bp&E�Y�Gӧm��v~��
A�	��D��� �!ߞ�W[�����B�,��4���'��v��o͊��5�i��4�
�PgS���vU/ �1��p�lf6Ux�W5�U�b�k��F`?����&rrȈ��-4f�u�&�	��V:��D�h�dKΊ?�V_|ڋ�;ŻA��C{)����^y
��=5w����M�o����b@����^��vt��(��qK:#���͉ 9�y���:�g�0h���$6�K�9�'�v[���r����Wr܃��Y(�-�IA��c���ah/��X~����K��k<�n�i,��ښuT�����IU~j']�e�����񎾓>�HV�]TG-yU�ߘI��;��+ٚ�i��v�5�[�=�t�"�DB/49痔j=Y�9H%I�]%l/��DN��t)8u��u
P�w�����*I&�#!)Qp<�$�vi����G����]����0Ѳ#�g&z[��\ȍ"�Y����+��X��d�1���A�s���o����ãrnޓ�R�%334�L6e!k�a��F�r�P� +��Oc��w��sn�W�J/f�"Њ���<a����.g7���*�=�=���6%#R]� wG;����O�[��8ҏq��}cP	�?;���(e16ψ�v�T/�<"j�vq����6=�ڤ�	W� 8�����w'��wdPׁ������M�{7_k���u<���>�ʲ&/I�s�aa=�
]��V���r�)`�a�/UR��z/Ȱ@�>	?`�0G#�Q�.�#��۾ul%��Z�^Y�e�0�[�(�Ro#���י?6#/�#����v���$���e��X?C�*ٌ�@#K���U��&��,g8��I�u_��LL��,~
ƏI}l��g3����K�g2��P�[�hj[y��x��x�K]_e��������T�x`�����k|b�!�~��D�2�tb��Nq<v��f��wq�����1��o-,��w�����^���t���I�@av����Z�e	^����vM�C;��A�-������}̤����$CP���ϩ~N�5���$E�9(�>�qе3��,js�9	?�Q��^�� ��'��nO'Ӏ��Z��m89�Sv���W���2�l-C��Oj�!W���^�י�|h���+��+��tpN��k�IG��F?�Y�d�����QV\�JJ2�Vl�5��)>�w�������##�������Ș�	����?�;�-����|ը�ZS6����'Э�ܱ�[�r�{�{<�-0D��i��i�oS �M�� 
�t���������o�A&�*��vĽ{}V�����M �S��:�$?�e�R �)��]8Ѩ��1�k�m���*/XA�H�b[�\��x~�Ap-�]�Qv�.��_�9�(�h�NV%0$�,�m@����R~�ըMY`�V@ƪں\��@�
�ƪ����s~):h1��w�-��W���r��זzuߠ��gJH�	9j�+��)�N1 3f2f�m�w���.�&�
q\-��.��S,�qaq�g
@B�ʾp*�|���kpj�Ҽ����8M���e��G���w{��;[Ok�;(��V��$���(*O�3�M��#q�_��P�C�p��7�MR��&2&�W�Pn���隈��o���'/�t	�|�hJw�yZ��4Sf���F�pQY��c��*$妰K��6_�9u�����"���L7�*�/i�M2����y�ĘTL��ܠkP8Zc��d��
c��C�DI���l���6H�ˡ/�jVSKb���x�R&iձsy�j\��B�����{�}X������K�@R���C��g����;�}G�fc�CU�/[W���I3�C�:'D��_D���B��������Bi�N�i��I�V)�{�G��D�v�(����RoSp����Τqp�rp�;>�SL!��3��)��b1��ͷ���bw%I{t+����;p��������'�������fb�6�{p�:r�0�ĺ��3I�k�{a �Dm�� ��6k��_"և
^a�u'
�l�(���3`s�P����_�U?yf9�]X>�e%�#c��Ú�2�'���"ۨ��j��i��;�;͞&�s�R��k:��v�[�9��h��kgI��VBNd!��Nw�Ω�	���Z���yr�BL�ȹ�4(ǵ�ݼx���__6ɿ����;�C�o���U��O}�4[�%�l�Ae�z���IžT��'t�>g'磷v��}MczL<��c�`��u!��a���=M���cQ�m]% ò�f˅EHe���?d��hX����Wڂ����y5]� Hd�,j�����\��j���՞�g���p.��Š�=��]�?����?:��^&4H���w�d�Q�5�D��E�l��7 ��`���@��x�<'{.����A�޾b̬C���q�N�G�_�X�a�݀0���]�G�V}���骦���J7�t�yul$JU���/������a�I�D�-�پ�,��R4�m%�Ɠ�d�
��K����Z�A/��J}����8���=�����H�~��p�C��}���q�n"���g��M����]���aҐBt^�k ��P�����P�޷4��sR�����%��y��B����"�=,��q���f֚5(L���\�FM�*��Y􃶫Hl|n�}�;�Ee�.���w����{LU�� *��E�CS� ����B����өH�5" �͉�]|����@�n"r=S�D��'9f��Ѯ���N��E ����,l8���5,T�0L�Ӻ������ǈ
�$j��VZv�)� bv����������Z�w������kc�;�oYK�o�l�Ԣ����#]�����{,���(ΌcMs,y��$��B;��+Kj�9=1k ��{�­��ݥݫ΀�+ۊ�����tO	����i�#;K��!�k��4�d�Rg�+���K���z;�*��9:���r��@������d)��;C�W���M�s�9b́�FL���t+@'@�Bɬ�)748X��-C��`�H)����x�麀a;;��ӂE��/l�J�Z�F
J���^�^2T\��O�op��7�s�LR�s����? �7��-�e����h�Z��ᩔ;��q>ϘxVZZ|\�}}M�a�j��r���FT��۷� +�g�_��^Eõ�ݡ���<c��?�=��q��R����NOȅo�ř��?������?��K�p�#n�C��WpAяO��Xw��>t?�ņ���1�	�ť�K+{A�En^غ}Q?�޽�E�=�R5t�P�oG��7���?a�l�+ќ�� ,9:�=���w��L"D���h+��h8!�s�t&�;Zc�7�^�����C�GMp�D���z=�2D�9�J�tw�(m~���57�5���㌭�^�wC��˗*nx�}J8)-E`B!�Y(^�ƙ�l��l��Eҭ�V��n�x?�q�"�'ZJ��1��FLk�fD�<C�@�D�����?�4��h�LT^�5�BD��fq�s������@+�c�����b� "j�[aB�=���?��p�d��T��@ڢ�[ozғߊQ�o9zk:�nl��H���їZ�����-c$�ҿ�N�����'A#������4l
A㾎(@�1�ԈA�P1�2A�_���>��(�|u�'m����4Hb�n���L�����k�g�&d��O�j���z���'i������=8��#.u���1�z#�	��c�ȣ�5�SӞ�H��k �h�S��G�p�Y,�U賹 L��=]~��պ�5����"���ޛ߁ic���lLy�ƱXT5ҞF�BT ���5%��ۄ�8
VxAO5�f��[�����~���"������&�����y��1~�	,���@Z�!-Qf_g@�|F �7�l��y�qt{�<g3H���_�R:��65��+���T��[�Z��]�I<��+�D��㢗�6ب6� ���Nt�,xOS �.������b
/I��S��l�M���&��r�#�/���9�Xߋ�e|+P@>�;�Dc+Ep��1J5$�m� ���H_���OK�Z,�/p��B�\h ��Vh���LpXϫ!p���Rpw�
1�e����5k�dp^�3�gn[��n3uB�M��O����<%�1d���G���;��K#D�;R�~�~�/�34U �׊q�iX!L�A� H()�L+�_
/���~��cď�
�ӓ �O��e5�Q���ɻ{��c�����A�E�_�>����U'(���oQ�:3,�1�o��|t6窻�`�y��_���Z�6ʂe��}�n˘�>�5Ď|!����ai�hs���W��O���g� �-�c�����S�㶑'���
(��`��M(����%I֍t�|���C��3��Yw��~������5�l���S�'���|+��{'���nc��$����ce�G'�S����5�����G'o���v�����/Z��� �|��7�v���~3�B���c|f|�Q(1qB�q':��P�5�>G_��[�67Y������x�`7鳹FX��5']���m�Iʁy�Y��t��HW��*��!��?F�������dn`��c�T܀� P��0�����4b�M	O��H����+�ֿT�>i�Ox���ocl��>���o9諟�o�P�Q���2��V�6�������4ʷ��gh�|���&%f��{3�k�qd�oP��6H^��r7s��*ʅJ��}��{�s��y�.���?Q�#.����/���*_l�Ecjh���#B����@y\y���{���ci�ǋC��PU0Ah�ԯQ
��'a)8؋;�;o "��ؐlͦO.� �
è�mi� 竫Љ7)�^R�S�$�P�J��3�2�Ej�?v�q�����P��N.f'��n）��x`�������	���~hj-�|G]�c�/�˰|��.�Ogk �uь����US���~m:��hY�ђ_��z�j��a�l���X5�Z!��yw(��V������U��NS�>0&� ���ٗ=
��QR��!�>��-)6��MVU �j��jdf�� +�U����Yȳ<r��1S���{�-���\5 "�,B�g�HA��N�P�0b�x!��.;}�`A� c��hqy�t�Ե�@&�s���Ė���y(@�*4����|v�����>�6����0�
��������ar
iw�.{��G1��l8w�O�yd+���F�P ޑ�Mr�'��:��Q ޝ��h,���  s�q՞{?�9R"o�.mI?�+�T�����9����S���8F͟�S��G�\��F~P��)^��DD_�
��0\��������Y�Z�n\�R(N*։�Ϧ���gO�N8б02	�3tt1,�E��09��>! |�����W���&c��Y0��A&�#����#�������������{)�%k�=[L
�c::��B�or�1U�7�#i�ב����*P�		N�n��d�Ld�@ܾ֢���+���>b5��Q��ؤ�.P�<�����/��jhe8���ѫ�?�&d����I��}ۯ���������YЫ�me�e�.�`����-k���ʨ�it[_��+��l4��c�xi�O&�$���!�G�ǐA�W]��k�Cq���Fm�\��PRK� ��@uȟI�/�����2ЋRL��g�uL�6�H5�ʵ$�+��B�0���g0�k���l��?��U����1�1T�Ւ��7���\����9ɠ&�v�,#|Ye�u�,9����$��9)��"����6+tX��~ΞLI])Lf��S�`�xw��67�D��8�'�����MZ��/��)������V�S;E
����_k�	� �o&����x�v<\%~�uP����)�v'� ���85 ؕY�� PU����Gǖ)v��Q��1�&'��V�Ś'qi|��c���"��_~BE�0��.��t?����|��k�M8�@�Q~�M�9�ec�B��ꏩo1�t/C(nQ��tYb<"�fMד��z�>Wa�|�0�����/�6�ܙ��q�X�S��B1ǩg8N�(���;+��@�͎�W�����|pAǦ�$��i�-��0=tb1����d4ڏdL�B�#�����2�����]��R�3LPʗ�8���6�}����[\�T����e#�<�f�|�>'����'V�Ɋa-kO��2�������������eS�;��٨�1&N�#��3�����O�j��-Z퀬<�ڶ,#~��i���iJ?��8�1B�gvB���WIjM�79EU�X"���ɔ��ɮ�B��v��\�
��E�����nv�x� �TVey�W� 	�w�dƁ���
�^,���1����p05�Jپ58=�O�nHJ(��{����j�7���|����f4��Z�y�Lʃc�h�T��#�V,�+�!3�qsÕ�@>�M0�����~ћ�D�M��o5�s<8k [}9���م��~��I�>��ŉ�9����h�b/�@(���ʫ�8�`����r�;a�L��}Y !J�Q4	ԙwd�c�[0L�A�F�j���H��ey��l���y	���扉�U N�m��g V���9W?�oNτG)1`�zr�[Y5q3Kw��1�P�8���U�;iz7���-��4p��n�D��OQ��ϓ�:��L��Yple^;�Jhb� H����,�K��n-�j�� ��g�@^Y$��ZǞb�_���W<�b��2� h}��r��q���e<��AU7�}�T��m�ݵ�^�)2ղ��RM6�I4���W}��cu�s�wv�F=�F9r&9�OG�Rr�J��j`���6@0��)$2����5@>~�Y�V®��g\d�O�Z�A�I�B�uT�A}p*�\Գ~,��m��������Eh^�zÿ[U@Ywq��'r�@P	
�U@�m��O-��KH)d��"��$3)6Wn�2��v��}!��E�V$�@Y����hKrL�܄��a��گ�Rf�M�I�TxK��kY��n �*���b���0<�G�� �*��ͥ�}���N�7W�J4�sh����
ǃ�A��`䯅>e��*����L������r@x��X
�D�d%����[�2XL�7hpB�m�ɰ0|�
���aIw �C2�&vVtc��l���pI��$��NN��~¬E�	���e$�h�qt#h�^���[� vM���e�ź�+�)(��j�������Ʃ���5���i$0�3#�@�wQ�`�Y{�ϯ_��N�\����%�v�-�d_�����R�&�Gj��Oo����,�7���r>1H�t�Y���g{��M�dF��N��Ԛ!ǡ�<Sx�j]�d^yK�ڧ�!�u>�� ��4|�zN����u��V�%�	��y,@��kp�r��=��Fe�H91������|�Ϲp���5Dԁ��=�&{Y�g����<9"��(
m 8,t�H&��Lދv�]��p�jl�x�\v��|2=YW�6��z��" D��:D��O��R�F���}�����&\��2T�a�8�r�҂�2X���r�.*,��}�6���4�Y]@������Z�xqw��j��G��)�-�n50���|g9�B��^7p��4ӏXk_F��MG�tU=��ߨ�S�FƠk`�.�&�߻�Q$�����YQ"�r}4:��Q`����X�DZkx�jc	 ��ό]���fɑ4�iRD���8����UZ��6�i[��w��0g��"4ݲ�D#�J-O�%�'��lϯ�̞�pUEp�ďb�-��YT�B�{
��n�㙛]d����e!p�����d�*Hn��S��?�b���G�ƛ��
�(��H��.U�����R�*>�9�I�jޅSD�WB|s.47dW����T��fUvrt��JFҙg8�g�c=����Q�Q��+B�Ŏb���tJF�}�-����ܻZӪE���o>ۛ��I1�
QU������S���6BWB@j�����`S�o�����L��Q��lx"��h2�Q�z� k�@���)OYf�o�T���M�*��jTB�B;���Do���IH�Y(�NK	�yl0�ƻ�f��w�mG�0�L?r�Գ���#�òБ���$h�E6�:f�q����4n^�ᚇ"i���i�X�Y�M����sX��fҽO�[��-D�߭���\�޴ԍN�jkʅ?��w&,+��<�fJ�U�Y�>'�7W�w+	M�Eﹺ��8kV�?"�6��շ��N�Yŧ�2�*�{��i\td���_�=Ox�&�|�A��NYZF�����`v�~�R)�-EA�Ɲ���P*�y�t�꽠^�<x7�ٌ]�{{|�)i��`���'s���+�[��ko/�y�U�7ܰ�s0�}��y�Q�����}�	��ȥ�p;��#�ר����dj��x��w���&����PxƤ���N�U�����j*e-��*�;h������p�he��i� `�����}��Ү����+�X����,�K~P�R��N��Jt�˪�[Aop�Sh��r�j� x��|l�Qߕ�+)f�S�]��-���A�߬h�je�Jfr�/��UK��$|�1��n�'��o�$7.�H�@@Ĉ�*�V�=y=���GK�w�������	��92&?��ͤ���Cp�#ٵ�Ρbk�j�:���@C܈}0�U�<큦�*G�������ҵF���\;y�D��l�>����r~�+U��lmh�B�y=/0v��S�~f)�u�ԍF�0DRY:��,#]UJ�x�?��k[�������7��xG�em9q1M�_Q!4xb�hG!`:��1�E�s	u�O ����69<������n�6�=^L���,�}7A��2! �G.��+�Ӿ�w��'L��<ü�c?�3��ՙ���&+�ˬ��&_�Ũ"#%�lXs�ۙ>X��dqhK���5�U�/i3$h���O�N�b�*�Gpl�;��z:�S�_��F-M+:�qE$����Uxu��}�8��7nwGh�������.����}��0��TE��%�	����}X����9e��Q��m���v<��3y��/<���y�?��#�gGӜ�lby�p`��z!��]h�C�_��"G����ȏ��4U=��ɰ�7E�)%����2����-;���4/�g�r�Ɇ5��va���5��
)�y��+!D/b�oMC��������@�OKI���<c����(��l�p<)�l�,�3Q�a^�=��{�f���!'fkK��n��,��X}6LӑgI:��.�@U��S��OdMHu����D�Q�Ǫ]^<^c�;jۣ�P&C��	5�k�m�u�I���a�ö��6o�|�����] m�	���:NP���7B�Uo�z�U��s}I��ۀr��O��4<4�}S{�'�]�Dw(m�g��Yl��i���$�S�87�R2�;-���H/�Zڼ%�J�e'��衒�^���͗n�|[B,t��]�
�=�?:s��>��ٕX����~ۢ�Za�՘�1H�=��J>Q�\��������S�;4W^�<�&�m������x	�C%�x*����"���d��K)׵P�<����[�3'qW��<M����RA٧������9�f|"��x}2[�1Uc�4�@O3���,7:ͮ�cӨj�f��@9�u,u�#/{�J��rtYEpA؍�y�v#�%`�i	���Nɪ�WΓ��뗝�味[��W�|���L뷖�p=C�V6f��7Ҵt�N*�s� ً���V,�;I����J��1v�2���W��`�H9IAvj1���(�w�����^�����o�1�.x��kʛ�>���t�~>��E�������΂|����n�*R��Zb0O5����K�g�z��ܤ\�ۃ�b���,��n��yw����PT}���T !���:�cc�x,OD?�H�茬��E��g����@vQ��K�2ń���{Fr���mo�YvN���xQ���E���^��� ����3��#�gsA����	X���ok������-���>zy0l�#l[l���|�CEa|�Qr��X���~��F��	�?H���x���=��z�i�$��ӎ��9�e��f�(W_�������@��G���B�\i5=���cf�tBNA�jl�:�~�cl� 1�a�o���E6��/��W�������n��{2�&>��sv�`��~t�&[*��8!2"���-�6����Vk����8�6��$���2��Fi�k�i�s|G�p�Z�	��jq��d%��}b\���iLv�pRƸ�}(]��ϻ �U��i�<I5�h��/�@ʩ�����fx�k���@�δ�F���w����x$��������(ԯ��o?t����V���[}����z����,��D�+Pkf�Ρ���f����C���%�|Hl%��	����N�m���SQ�!����(2b�<�}v����;XP6��aUs/|����7)�hw*ոDi��~G����������2@Z���B�^�m?C�a�N�G�Ntw�����Fa�����̔��Y��X�P�����g=w#u��sG���D�Moi��^�G��g/]�W6E��:h�RG��!{k-k�s�r����h�P�����Bl�*���I�q�M���M��v�â@��ǐ��@���z��F�`��!^,�u:b��ݨ�,鰕N���l��H� :u��G��	_KTZ��{�v��6�������Y���U�~�[�x�O߇��,,��J-���t7����QVtb�����K�6"?c��)j������=���F�Ϲ��ّ5�Ra���q����r?���Z:5��7�&?0��x��������|�	�:}���r��+�IQ��0.Ҟ�E�fdb`Ϟ�*k�Ў���$��89��^(�@�wծ�"+`��5-3�7��ɣ�e 7��,���Q;A�2^��b1��ۯMq��׌a��7��{��4�
otB_
�J�ğ7�3!Cvg�˃kʐ��4#�H#��%���=?�|�+����n��ҹ}����djڱ�5�}b��Yi�wlD̒�A���n��.c�iQ�}K�.n�"��ʳi������nX2����-v��f�'������Y�>k�RL�O����O��<��k�l$Gx�p�$�%I����Q�hWe�/�?��P!�9�:O6����ڟOc�O3_�W�.$JS����*��}��뤶gs�8�w���L��2�n�9oRvŠ���:�3*�Mykә��:m?���2����:��Kĉ�o�}���իz-�t����L�W!�Њ�`�"\��_?k?!v "J�����9���1qN��k<��]�ZYA�r�v҅�*�}��Ft2ts1���8X����[��F����w��D��E4�uG�,�~�I&�����ƺ� ��Q���-oO���Ԅ�
����&�r�@�2�ȶ�{ri���k��E��p���u�s����t�+QS�s�X�
tޒ����R��b���h<f��5�^�{+��RX-j�Z�su-�J�K0¦0���m>�yQ��?i;��!�����4�J��u[_��s�C�~_G�yM��
�%)��N���c̈`Yf�w�������֝��[�q�S�!1g�}�Ҽ�z��3��?;�B����iT�1-�$����D�y�f��F�F�����������Gw�W�H���i�x���Wj�9N���������S󐀭M�V��I�����ݢ�i�aQ�d12�]�M��K�D�@����^��`��csq�� -�6 �e��:-�z����� s�Z��-�X�Y=b�E-���5�++��?����Z+�)��	Wh >�y&��O�&�����J��t��T����>J��#�*� ��v��s�C�[Ֆ&t�o�;�%��vߕ�}�Č#<�(��8f��V-A��h3��_]>�wm��S1�:�+� �\��
�;�:��&fSq�b͗w�_/a���pBŌN���J���'h��˸�C�(�,�ƌܤ O�p ̽w�EO�J��K��0�}Ď/{z�%=T����}�t0Q��K�_Ͷ�� ��̤��#�k�!#o|���Q�In7v��/Ƭw�?�80�1oR�jR�q�h��,�u�}˸��7�������"s�z��� EUXOv�Q�K#�Ӟ�n� �&Q�����i�з)�yEҗ��sb��	��Fǈ!���N
���ya���6���P�8��{�Ǖ�Jx�o��3�(����[U	�`f�q��⠇��h���DpT �?m"~�9*ު/�-�ؗ�A��5��uI��%j�ݜbI|H���������6��6]`vw_e'm~���ۯ�~����l����yj�Z���aN���9}u��K({���{5C[_|�@��V�˨6�����H���:����l��P��D�z�L�?JǠ��r:�h��?�n�l�Ѝ�}'� ��F��8q� P�e�W/��%��I�'�]
�6��6�A��Ԡ-}���=�g������dԙ>KSP�G~5�s���OY��!��t8P�~m��ŧ�q#�lЀ��jڟ5oF�Ο����qq���z�u)a���To��y��)eo��N�xn���R��箖��mᆷ��x���Ta��=)׋�I���c�ӄ��O��DD��\CZn�XXi����6%�߲ap-m gZK)���5(�!�s���b_���Ъ�w�f���U$�3C/����k���(�հ{:	�7EZ���� ��<�_�S��9��&����<�!��}� ���}�X3D����d�K=Hy_C���c�_O���$3d����o�#�$5��Y5�	������5�O��`�&PS)���V�;#��ݧ���5u�K��~�=�7!�?I�m|y:�q�߭���_�����V������(�a��w�e���p��z[J�a�7Ǜ�5s�=�9�n�(�"W��J�h�?�;0�$x0Lu�R�Y��
T��� UE�i)�}��'������^:�L2�X �+�e�2�`ؘ��=u�/�i��N�ԂG��Hݬ��W������~{��҈��(*�׾���������1��T�������s��T��ޓp���2���^�?�h&hզG�7�2?y*���G��5����g�����8~��UĨ��"� 	9)���\�%��`7v��-N����(�f�؁���~S����q)����|�r{߇U��U�@:DPR�j��=H�P2C�J�H�����PC����C����<��?[��?��r��u�u�+���Z��I��x^a5d�R.R��%��m99[�.���a���a;�6p���	UUE��)�.<��`4��OS)@5�4��P�_o̩�ʥ4 �^����<���v�rX1�����53���zC��n����{sxn&��@�s
v��;Z^���j��ɺ2�K�����7�����E���F-����j$��u��	�6AY��t):����t�������RJN}��pq��?]7����|�vc>g�ťiN�O��_���Ͱ�a����RǓD���q39����y�pŔ����Q��j��d��H��K�ȏ�DSL�c���]�����C1������}?��-=^����wQ�q��ﬠ�G����2F�!*C��ZB�X$�Gײ�Mm�YfWr <k ��~亷d��any)@�U��evR��o���	�}�,,'9��R������tuK�R�w!�/�/(-����,34F���B.fW�$C�?�T�M8� 1.�
�I8{7�;��CI/ז���7-�u�ɗn��Km}�?h� BI�|��hcV5�Kqa��V=��?x2pR�Dr���=��0�иjL����Y������ň�T; ��6�ƿ��
\P��3
�++�cu}��x�7bQ1[@�-lU`��o��'�:����+��v-��	;���'m�Z��~S���16ߺW�*;,<�k�˱�$������~?s��M�Gw���R����rt�.�Ykv좪�9���t :�������4��^�&
�bt���|���b8����kH���K��Q�9��<�;�i�<t�#.���L�pT'��x�Ԯj�9J������!��#@=WjqsR�36ˡ�[��QߣU���4C�OK���ҷ�_0����DØ
bX�0�͗���S�}9��6m8%}rm��(�<���dm�WX���Ƒ1A�Z^�4��}�̤�� &���UI��E�D~����n�;ڴ���)�0��m3�`�ۜ��D��R�(��uuX�^�4Ɲ�����Z~��I�m��z[e��ӽCt*N��-S]�Ṣw�ؕ=B��f�����*�c���e��7bv�\���>�ڌ�2��
za:���o^�����;U1�8o�bnCJ��j�0���������3��W��*D(z�c��h����n�d+"���1�y���M�'��]��ge�9�9�8���>3�q���B��6o^�y��^in)�����r�>M�bb�� D�KNK��;j�6��������^�h��Tl3ˋ��9��� x��`��f����*5pQi5��ќ�������>��S}nG[���$�:���k z? �?�L�tP%\��jY=���],�t�c~ߢ��sQħM}C�Uj��U��@c9(�4�5�9��ҳ�t���`�^ˌ^r��ǟ%��_|�6��+��{/���p栱��̐���SCaA�F܌��>�Y�L��?.��ќY?��Y4iq�b-�'m�򭬱���^���s��n����Z�r�\V�XF9�<jh�C� *ol���]�WR�u��(Jw77���G����~0ǓLe��v��(s,����-��ƘYi�D�ѡ�B��jox��? ���y����4d��{��(��i��Ծ��$�r��1�'�?}���p�JF,�����r�d8���[$�~W�̑gI�3�|{�̗0��~�������G����{����F{U*#��0U�)��up�*M�@�Z�F��!3>�0-+��:j�0����ƙc�z������+�n���ueRq�}�
=yt� ��j���7#�B��I��(�J�;
'�٣I��N	E��:3U�x���<>ʼ�#�S��C�c�R2�Kp}��Z��b��E㴇@.�S�S�q�����M(L�e��F`��Z��8Z�㗥d@��F��M�	g�CXsl>�_���j>������is��'�(��Z����H����̙��ɪ@ã��&�-�n��H���b!�]91g�[�}����$�Y�xA����Wv(.;�:��J?n	:���ز��BEF�� ~����I%���`�m�6��w"�d�6��8�d��o�NohY����oTXgϞ��:P>�P%X������ՙ�-3!�A��3vv!}���BTqXpv�kkcc�U"����5�5����Óڍ��r���=��5�=\K����Q��ꁊ���ml^�ЯS�>��L�E��&J������Z$�mW�,�����5�������FTg�2��rg��㩽��ӮH� ��*6(.���)�u�p~���R|X�{P��KC�h�B�ڌ?Yd]N��5�Rs���1�:t�����2z��t����0.���eaJk������h���k�CP~�P���;���_im�%��&`��?�J*�_$m�+������J�k��������Ҹ��w��}�������ؐ�D��ٳy�Cq�@Ъ}A�3�C�+m��ƅҬ�HPX[�"~�F�m���e�Jf&�\��PGyee6���r��ܲ���Q��%�*�O�ٟ'�t����a}jo��L�^��nS���5�Y�-�㼭~Hv�O���[ǅ��H�o��L���jr�ϖ�n|<Iw����}�6y@p;�:;�˟��d	�>�I��V��������9bA�Ж�]�㤫l���\@˨��m�C�.��Z�����|p��eiOܤ���� 
���w�q� �y��I,���J�ge���s��@v��ٛQ����-�oE΍�J�̻�~������f����AB�3��6v�V�#
��їt�1�i�Bx7{��s�{��j��A P�	5�	��{��ך�����7��\�'�����囗;���X��"�Wm�~E_#��>I���<P��xM������@R��oM��'%ȋ�į�� M��/}IQ�m%{�ѯ"����`��t����2����d���i�q_�Β@�p�V��݃����.��b̷qtmz�> YOEb�
Z�!ӭ���J[����C����@o�I�����d�9_�l����I��G������7�82
�#�f������S��ɀ��9 3@�h��o�r03?{�|���'
��r #{�>�$ܱ�A��tT�W��U�	3'�C!VB�d�>�����w�ߚ��F.�7R�[`��l�|m�?����<{m��<�o�
���N	�Γ���~�q6���eitߦ�ƏcF=�p���7?����n�O�a���|�g��`Yj�բ1���7ۏ<����;WP�+K�������v�Z�#�UBr	(ҟ����xӍf��틓E.N��aޥD�s�1�t@��������i4i�'&�?��ڿ�vT���9Zn5pp��^&�)-�h�����[�v/X���W2�??�Os=2?��d�m��c�,s��Jp����rxYFs�CKk�,��^�..v�sΟ���S"eP�V�c�a�^ �A� ը�'�fɉ#;J��{�_�\9��-VZF>��Nc��H���&�ƳQy!�i�BB���qc��J՚u���XZ�l]�m_�wH�|�jG
��I�g���	I8��:�8����e������#x��Z�8Y�z�Q�8����l)�a��]Dq�{�x��~Lub38�U����~EV���!�8*��R4i�hk���֛_��}��9�8�b/�� X3�%�sDO��������.�j�&��]����u�ܣ��O����a�~$F�`RKdl�����sn':�"uZ�|'�̩�;��}��5�j�-��f7�
^i�������hXc���h�h&���J���t��-d�u�'�R{m#D���r8�s����%��2vG�%;B�t���r+�ۨju;�
فW���u`jF�N&��gC��T
��>�`��;��SOl�j�k�6������0����0J������H�+b�Ϡo_��c��9�U��Uo��L�Ԯ�U<S7>�o�O]K������Uà�
�Z�StN�m~;$�N���>2w5��`��2�S�;��V��kO��������&Ǻ;So�����w�Jɹ#��i5�a��}���,JQ�2����H*n�#v�),Y�&��+�>�������	v�Ǐ[�mY�"�I9|�WD���B#s��]+���>j��#��f}R8@T�W?�,,H%�#z��N���_~/�]��z���.��\��D�G�a:�g�tp\��	UU��%2�O�+�]�LJ'��t����M+�W��tU��Z�� ���4��'��
.9,�fcXS)������Υ�G�+��hKQڞ�GU���������_鹧ߏb���4A�t��5J=+��T�hO�ɼ�_�)�����U�;#�ú��E��'�A����q3=����{�0#L}�a�Ѻ�X�Pp��$]�j�y@{���ll��M(�&s�]Q��޼"_4�=�1Ax�`�im��6<�+Hnv���,�G��2�[?���~���Jo� �i�twU�F�]�_I�A�KջY8��W��NU�5M�<���Z���|f��43�7���<�b�~F����&�-LѪ~N��>8�s���X����K_JxIߨ͸��'�&g���퐑#;vy�����.�J�Ne��#glW�{yWww��b��v���`�{В�����eS�m)h�v���r�{�b�΋r˩�d�a��������N��zf�rW<N�{����k)�J���������n�^�t ����ś;�E���+S�N}�c}������WL�ο�y���:EqmH�=�	�(���iv��A��ۉ������\ҎC�(�ra�N�� ����;����?/�9�qb���pW�Q��ж��3=9��6�\����^̳��(���ƣ���|�;���
���=J]�W;��~B��_�����S������u��Q���f�y}��hy~u��m�vQ�ڱ�=<L��C���Z��	���䉄�h�p+�k�O@�t��|�J%�0�jC�h-f�����B3������'�1y�e��/:JXfe��Iڥ�b�i�;�l��&jT��D|�S����ou�z�/����3V�n��@`�Wwk���:"�j�3M��5�^�j��ٙ��ێ�A/�#�l�ޑD`��*aJ;���7q�9�T�n�a�ݙ������6��)��d���2��v�d��iG��S�;�H4�ov~T�KV�禝�G�����;Ny4r��:��eW�!\?,\�VQ��<q�
L.3im��[�����G9ĥ��\���Ҡ�ɡ%	�I�%�Rt�@���$4Q���ᰮ�������h�0���xs��p"14/ ��(8}2���/�R�����C� ��t�S��X==�(��ld����ʺ�6�Z�A�s�_J��I]�Jz�(K����;�����
�S��'Q9��0ԓ2E{�z����/��㦜<��	Ykw<C��f�ײ��%A�q;�J.�g1�I��>��rQ肸�r� 4��,;j�ś=f�3꣊��1���tϦ#S�.ˍ�P��DC���e��<a°��d~����1�Ҽ��]	+b��Yut�U�cB�V�O�v�/n�{e��<{[P��������N}t��U���b��/%c��x�A�ÐddL}��pF�L[#6&�e8��5��a�9�5��T;�/X���.>rs�j��Z���Sk%�%���p�Þ�{�s��#�u�Jww��2��?�	�q�d�ƺϕ�������>���U�ب_,�m���6+�P-�v�'Hr������&h��5�%��ٺq�1:@�p_P��Z�D{l��� �VK�{~Z]�=�.hZ�U-�29����Zp;:�۶�]�>ԙ��8�`h�����Wj^96�9����#uB�E��,Ѭrf�FH�3r���5=�� 2֚�N��e�f�����(�i��pֵ�Z��{/P%���K�v�����W7YmY�6����c3s�<��׿�.:�+�>�u��l$�W�i�Mz�1U�E�є#���gd�Jj�^hUo���Ml�W�<�P�����C���Q�8��ķ��tbr,uU����D>ډg��2$p�Z���Ƣ�� ���sV)8:�����GN��E��:,���0ܺ3�L������C��W��@>���6zrX����*���t���Gk�U`���c�W��X�"�qku9y[&U�]���1�7���A%JY���F��=u����у�g�YV졣`�c��Ȅ}��t4�Z��r >��A��bz�D��
N�`�� ����F�cjq��J,��U�e���u��n���5������^*	�������8Qch�����8���y���~Ƚ�+��ߪ���<��2м�L(
�z�H�S���<&A\���^ܒ'"�e���rx����˯�q���S������0}�46��|��r	�mP8�gc�^㮘nT�DV�+ɕ/Jh:�N�I�9(��{�H������,n0�<�Qv�Sv���^�_�� ��=�ɉ�B��U*ģz�@a��`?����o�82��_���wX�g�I�E~Ɉ@v�A6
�+ lD�_�p�]Y�VY��"��jb^���tKk͝�\1��"t�3^�Ɯ}�����-�yA��}/k��U�
�jy���'zb�z��}Q���p��{�ޮ��a���yi��$�O�mY�%}�@�Bz�PQ��������
��Z�|��)|��t�����GAj�Y�䏰]�W�S�B���l9V~�O�&�w_��k ��Q	/�uc+L^�|m�ž-ܚ��@�����뤖�urs��;l�!w�b.�	��?C��e����1֩h���k�hG7ӂ7��^�g�Ld�=͗k�#l���8c�(��
C�m7�@v��&ʀ����ڻU��n 
$������kn�a�DOH��J��޳1��"�U��L��j�s���m����Y,��Ve|g �>,�bN�K�8�K�G?�x���q5���r��-+&��J�=�-�v)ﯨ��m����[�z҈�JأlP���,��j��X�"vKZ����6�t����V�����V�C^�X�}`�����Dll�ܤ�X��2Dv����02|!ۑ+B�Gv��r���\��v��u�v��S9�K��oS�)g޽|��o?S7�ܔ� �[�5�ؐ� 2�lm���#ųGz͊"�`����[@QZg���q��3�"��C�
(�K��/y{a+v����XGܞ ������s�6-��1�/�̴��#<��6�l��*}������`�?������~���q�Hz?��0�m�˸'��Y�I�'u����ܑ�{Q�X���n�<h�d��6������Q}	*����wgC��4NP��9s��S�n΄`�9 v�Oa'��������\:�������U7q���-O��^+� �^�U��1hg��)}��9��~��=6��'T�/��~�-�(�RX���m{?r��\e���콻e����ޙh�Lg����j����vkc�=���g�5֊�*`ĕΛ�)��8WL������r���_r>��n����)ޫ	1��w;?�����;ͳ���H�R��ކz�"Q��Ѿ��C�,d_sC�D�+0O}O��U:�<�]���u?�ȝzXEۦx��K�x3��������!?ii˨�<�	��=�F;�����2.���T�c�$�JoH|T�sT�*��=ڗlx�ͬ�H�u5[���S�kӬ��>�Ud������ّf�q a3T�U0�:�Qa��-AL0���O�	���u�<��98�UȎR�a/�ۇ���ȷJ,���3U:d���RyE �� V�%�Z���]�y�Y�w�JtP�6�̊�D8�=�>��L�s�$�Q߂*F&�v�1��k�0-�X�x�7r$���+g"��F��R��������7_��Lq9IO/�?��Uɾ�=X��ZȒX�oZ��l���U��1����&]Gs�&�4� �GOI�/oAHE�Z��U��E�.����a��UU��9 Bx�,oi���b�X���aB���K(����9�óR���Z�uX�q��,-�C�e���o�R�M�sT��W�W��al����`G1/�x�@��� �3��7�S�(0=��[So,N~p�Ʊ$���Uu�au���^�# �c��r#� ���g���z|b	3���j���J:(0�R	7�,Y����gu7��Cg@��CE�K=6%�����V�޸2���S�q\>r�	�;���l5�UspZ��Ϫ�ᴤ�?�i��B��h�m"����!�Қ����	���ڍ���H�o�3E�����k ��y%�_��P�@lV�@e��]/��#�pX��rQ}���	��0t.n��!H/�k�$�}��)�1G��sD���9�C'j��B ��g�C؆���[�	*^N��?��Mw`K�U)P��A)( 1y����0Snk�{{��#�"�7,�%��}Pŭ~�#hm�ޞt�f%h�,�/������c<>suIC}����%�����A�4��>�c���e�+C��<7��/��)���aH�{A#G�%)Z���?�q1�U��G�Ǡt�*��ꘕT����댏��lT� ���<'�a��K�*�U���� ����"[�P���`�٥+iA����g��zť���G��%9�e��T�N�e=@9�]01�?��N�)����9�$8����"��-k�����������)?5�}�li����D���7M@�������ω��\g�-��+���V��.aH����N�Ɉ'a����R�m�����Ge-b)�̔�jM-�ǹ~+�"_�ja��C �;=��-���a�g�l��^����S��*�dJ�=z�H�����X�b��^��+�N���F��'�p���=Ʃ�&�%�b���͹���-E��]<��5�ҙ��>I��ӯZu���M�^6~6�2i��%�p��B�$p����Se�|�	��4�������� �T�;�H�ة~����W���U
�z3�P��#���IB	�7��
5ֶ�Vmv�Toa���c�#��55ϖ;7��v� f�'��9!�Fb�G]�@�)��d�3;�֡���e�N$	5=��m�Wܝ3S����65��44y9Ǜ4m�9f�=b#W�&��[�DUo
c�7�+SP�h��k[���y�>�H�΄��K�Y-
���n[�?���e -�-�^I�Gҷ�i�ѦǣPq�u�}r��=��D����n�?�uKW�8ӻ�ɚ����� �֠���6���J"P���Ƌ�M�-Q���W��9crΧi� =�:��=���� �('�_��C7�� ���@'���E�ͱ n��h�{p�/�r=��ΏO�x��; �] �v��u�8U!��kՎ�l8a$1���L~A�C��q=6�~F�z����;��b��񦣮��Фw �Uֲ��q#o�Z�ڿ�  	�죊m�vP	7���)6S���sG�V�����T��=�WV� ������1D�;�h�>���Y@�%��S B�>/,�HE��!�{w}uGΠ�A1�L�%��P;���E�4vTB���g�-1��/ø���%�gQ���&c&�M�}6�5/���|tF�O���M@�p�T�0��#�=�&�(�W菔�r�KOL���23b�!l�%���k!����pkk�]�f�#�]������x�v��A<^?%�o#����D�j������U81g�>�Һ��ӧ�����Kz���Y ��zڲɭ�9�$'�u�ՌU/Ů�{�� BTug�A�cEI���x�"����Ȩ��p�����U���0�|��̱��N��y�����nІ��X`'����^`츷�P�I���v�������(�?��܌Ֆ���zl�>֫�t�1۴.l@���t����Ð�/��f�ӆ�u�����8׎W}�>z����|�n��7�osR�+w��u�}���k���n�BZ��qmp�*!�H[���еfb<�<������1��s�]�{i�K>��EG��G��;s�5Osy ��k)��q|�񹀢 ]�P���0��Y��G}ڐc?@������H��H����� ��|�z�m2m`�]w����
���Nl�Cm>����7��,���/.,��Q�it��3��Ν���b~���U��pk�5��D-3O�ak_O�-�gQ ��$,��a�/f M����� NV8���GPIwTMʡ��Z_U��.7���R�1 Y]�[e�Ic�1�04��5}����K�:��Le�gl%�}��[<�i����?\��? �R�Պ�j�{B���@g7�y֯������/�˫�)�;t�Bވ���l�zCG�[T �R��m��7�`X�%'���B虫��;�)�����>��K��f7v��Z��ǘp��y����������j������7�����e�%�^e�	ꣿ�}^UR��� ��ky�<�_	��i5e�H��ȗ9密���S2 ����qmq�˹lPx�L�顊 �._hlx7���Ўn]�2+v��[,�Kj۾�������>u��A Q�_|���NFp�V|�t�E����+�_®�� dC��8��� ����ƍ�u-<Ѩ�y��qyme�ǉй�?��no:	����8�!�u=��Е�&5{H,`��c������O���j��T�=<�H��Irlٓ	�#����I��FS�%�aP��5��4솩q�:��B�7���D�L�_X �xT�S�Wz�o���Hۜ�$��~�#�Cn�*�Y���`ϯѠSfs-�2.���"L��E������d!�C�v�fs�t�Y1�e�v���G��T��J�'�d����+�;P�ML�>�ո8��q�t)�ؙ�X'H����F�5ޣ��ӭ�� :�,y��u�@���x�@�!O�y�� �f�Ʀ⌕0�{�#[����6XA
q���yg�>o�CO����x�`������
�?�|�"�Qv���-n 6�9��_9�+�2��V͈� ,&%L<f,��Ɩ���#�&\;ʅ6��*��	ӟS�O,��1���V����L{Be�����7������E@lx�a%��>V#+�G�ih[�)���g����
���7�3V���ҟf���}�L�ͭ
s"���mM�D���@��K���s/�a�|�9�����I����J0޼e���w�r��p�?��h�u��Tfp_é��+��>4v��_��]�6�q,�6˲/��s��##G��ja�E�5_���_�,�%5���~����Ā� �Ta��\8�i#�n���&�a�@�}��^qN�8��K-!���+�����i��fwD�A�*O�4>a>x�f!s�Q���9P"B�`��޿e�-a����$�i:���=-J���ڡÐ�7_M���D�6&Ѕz��(L��7�Պ�@F�u�\M=���ގz��(GH��M�D����uϽx�ޤ�*r�)�ԇa�S�Mf~F�������+SyqQ��)Yh�5Өw�6�����bS;���R�b�8N!0���t}��+�:H�;���n�V�II�=%gwٍ�qߺ��xI"�F����s�O�E�Mp1mj�*��^�O��l���q[ Ȅ�Y-�pT�+/\C5R4��2YV��7��*Ӵ����ޜK�&$%k'�l��Y��{_��[}��\܌_�* ������7ƤL��`��@�{z:��@0�߷��R����b��Dך�՝�O�h~���,qmZ����譩�)�r�֦A�a��9(�@ͣ�Wl!��y��s< �#e[�N_fLP��Ֆ�Y-�wb�uE��i���O�kH"�z�S��|�<��@��f�)�w�a�-�A@�u�0��t�sC&�6�+���l6��g��%��쒌�,
��>(�!����SS!��q���YtSq2p?���z�_�G�+�^O}hП�|#eЙ��؃*�M>��JB��S>�}�_6n^�˨�|Gߝe<�7� ���Ạ[��'�r��C�f�J�i¬c� ��,z�ƐY%���X�3�?�ޤ@ߞ.�z$P1%�?��	��bH���E93�P_ a����v#����H|��1'�j���RJ'4Ԙ=W�r5�u�
6��.�K���K���Sl�y�c>���5���{�>�Uy�5�Z�x������܈�OjGz�0���G}����*i�Ɲ^t�� ��L�og���+~P��h�>{���m״{'�����L�œ;�V��������Oj���A����jW�D�[��\s����,|� �����iw��V�`D���z�Y��2Ґ�6�aa3��6��Fǅ\W���zTt-�t�`�\f��0�J����{DY�p�)��|�H��{2�,5���*�6��\�m���nCe慨�0������!�]��h�S�d*i����8�O��T�]�>,̨-l�͊O�z6�����++��;�N�V�-%q��'���|�:��b߿5�14��'݈+�t�I��#m�u'�Z6��vã�	���,�ukE�N�d&�����Mq�A;�*�i�|T�2r��ϝ�5�h�����m<?�T-�Ƀ��.�N1�"�S�C>���h��L�Xǲ����(��b$�z�s �U�y,�1�7>C���w�R���Љq�u'B/�,~��ɌC���`����YF�����<�
������m��Of��͙wY&�i,�.RW�0EC3!����_��sZR�
�j .� �z�L�{ڟ�1����_X��öh�\�L�a4���,#�*ؽ�>{K�G�Dy{�rj���Y	 `/�pA�������aP>u�ʞ���_�:���0��ֿ�&}Ҵ]#'mk�92��/��ND�isg��b��\'�$�y��w�-͉�M�u��	��r���Wi�5>�~l�}������ =�����=�?M�AB���.�hq(�n7Ɂ�l�Lnم����l�	��%$g&d�@>B�����̛�C�����#��ߗkM3��c�>f�	s�5�<o�Z�oi�����:Ǯ#������.C�Cέ2��@������u�+���*��f:uȕ�J�35#R�"3f���]�{� �o$��N;��Ƶsȃ.�+_̿aDB�X�%���Tx�݌C_���2����|[�X�����K5�NX��x�M���V�W%������{�_e}z	���JJ�o��P���S�XȔ� Lru*=��f�����E��\��<�.BPAOd6ĩ>ͫUGS9����m�윟�X�[(�"�Wf�F~K�p'1Į�����c�M$�����M���+&má-nB%���c�_BGx��m���xk�8����A�$���{���e����J�����lw�/8��w*Vn�{A��'��o�M���T"~R�:%u�Q�M�V�+SM:��<sR,s�w����p;�+2+e��3藏���@�-� '�9de]�C2���J^Ss��� PM<Tp�U-50};(���霒+wR4��G:� �lbd���Ξ�}p��������ʤ1�h�Z���EAR�>��n�=�C�����@0�� _ă�'�����Pԃ�M��_�6�
�olU�ݏlN�3"�$Q��YW�@�����&����2~Q4��!L��QO��(�c�ȧk&�c�r8-��c>3�%u��>�X6+�8����%��D[��W�E��pR�"Eb��2�)�@�MG�wˊ��6C�4�7C�� �����u�)X���(� �l��C�����dY���zR��r9(��(ě͊�v�w�Ǧ=�	E�'�yC/�� (��+(�-F|B����F�-����j$�|j��y
U�[0����T��PZ�H�P>z�q�t�T�:�m��q6'�bˑ�o/>jT�P��3mT�P�W��_YLS��m-�}�-1J:߁�}͝M��A�.�x���^d��z�ⓝ�f5�H��Wyo���.._˥
2Ɂgr��Hp�e���4���~�~"��7ϗ1���$���6�H@��SD��3��{�I�Y�R�^� Y����'�@W��"&vڅ}�u�`�P��l�%�=1A�#�_���+J���;7Q�]�ꉤnV������Y��E魊h�.�*��*�1���xmg�ك�w�a)n����u�Jr�+����k:TIOm�-"����x�qs���x��|�B��퀊�J���JA���a���r�>/h�b�ӕLd�HPQʅ�Y�^!E.��lc׎椴X��D�,dG(y��s�A	�PSU��o&A5�.c����|��T�MZ��� ���@�|�v̎�ޞ�5c�ʙ����?U��nc�$Lʒj,��(�z�N+'�t�+n����H,�<��A��#Z^�}�YG	O��]٤U,bpoN��D$�6�X��**ߑQk1��֚o�\\��p�n���+��.k�h�ݺ���Jmʷ�gֿ�Eɧ�����I�=�� @�C	�����q��<���87\���.��6�iP�=�	%��Uk��Z��^��=��*�c�H����1g��nZ��b�ܞ��T�֔%���3�h���<��	�44ΐ��J���wD=��/��U�~���FjqF���б恲��=�h��=��'��Dw���g�O�E�K�u��V�]�*�:��UUq!��~P���Ae���fH?V��.�R�o�k���nPO4e��F��3��Ҍ��²��/��iy���U�������8�;���-�#́ܵ�g�b�cE�ɦu�����A�
H�=@bS~�_Þ��P�w��;|kS��n|L�%TZ�M,s5]4��Dg�n_�d	cG�i{�Dﺭ�śv�K+1l-�H���&�86'�'���l�U�w�>(5W�2�:팷�19�h����#��A�S���~��NxR������+����D�x�V�K�%�NnǶ1��&��a�ea{b��!L�|�G��יp���V�v�ϵYo<z��~��e`��Y3��4V:��1�*�N��zـ��)[6Q�}�\dS�V�wK�~ӎ�x2�MWeA�c����M�x	1J���`��jqr�Γ���xL�xD$!4��{̧�Q�I䞆���|����F~$L��1h�z������帏�^��s����ٹ��޾��Cњ}�1/��*���Z��� #���5z�����5cw��ʴ;��4ua�5ջO�Ƅ���L%�I��bvT���$�v�]����^-���.�AfY����g�Y�4���=�7'%�L�E���ZDD�M6�R�*�2� 5���$Oa��a������ʫM�F���SDC}"����B�݁��ƞ�����s�<��~���8�7;;���W��_'�F/�З�F};C�L*��DB��_r������9���c1o�4-���
n'kk{�ˈ�փYN�Y�"��f�?B5os7�w�z�2��9��Y5 �4���B�<�� ��K���MZ�*)��<��D�|�<r�]$<hR��w�jړ�\��t�T"�ʛW�y˧�:��/��W@	��{��PLa�������F��6��1۔���J/+~/e%;�������j��1����A��0�Kƅۘ�k�W�&4Ǉ�ǳ�k�v��]b���@
R_��a�=Wfq`T�a3�����ڣ�* ��]O���������>����M�Z{�N8�"=e.��}"y�����U7��i�N����l�.�C�Y׽����j�����vQ��#/���:<���(P5Ӊ>�u�|��C�ﶪ����hi>�	�^�\�� ����Y�}��9�Z1f�_��-�h�a^�^q�%�,� ����٭���ۯQ�13�86W�E7�����@�#(�1�B�*�L�o��p�)�]��4���Xt\��������,�0�p8�C]>v'_��]������	�*9�ɛ'H��&������rݐ���Oi1�8ݗ]��#Z7��7Q�]��_����*�=Һ��.�2�^�=7w�@6˗K�s�ZF_�2x�֓P��c�Ly��ٷ1��{���S���a`����oh�+#������Xޒ<��)f�����[�`-�q���*�j*�1<C�jFNU` ��e�ݔ�C%J������̎Kz�������ߤ>o0FE=�Ѕ�M̓=��������k�S�@�ny
�F�(� Y.=/�{���o�i`�
�q�$�
+�%w���K��V�#@�Чګ���2o�F��{��M��c���'��O��*�=]$ʭ�wd�i�F6]����[�eWo�f��p�䤮�~!��O�|=��$k�U˗�^˝6��TP���w$F�v\����`z��B��Qߞ��Z���L�3]U�i@��ϗB|��N46�z��x7R�>��k_޶�r`������4�1�G����)���Iqu�N3����)Q�	���g�)�|�tSO��۷�_K&V�3�I�������U͡��XQC�
���~��S�z���q(��_�
�g�5����5��O|���R�!�ĕ��!���]���d`��ӫ�(����B˖�����qÄ�
��L�g3���y�~*��*��=a�K�9[�Yr���gu��K�=7EO<����V��6`|���PN�J�g�"�%��OA�N��1��Ҡ7���t���!��:d�+��->T�R�ĭn���L��~׭�jY���D�6w�}���!����$Wh�1���h���VJ�W�5A*򜫑�>��w(�=ne�rw;����-���)�rC���׾���ۊ�([��0}�F�ޛ� �֢���>,���i�f[���"������Q�-
DY�ɍ��� �w�YW��~������&�$�4��Ic}N���x�u��,�ՇF��Z���Tp'�m�1�<��{:�v���6��-�����ʢd6L�G2(��b'��xl������8ϟ�W��:[���g��pn���*�P(��=i�f�n�W<����iC���|���)�nf�o˦� ���zR�s�~bc�G�m����<���@�c'����PQ����(~U�ŠCI��i����!�r]���D��A���n$fFrh��g�����=z���{�{�s�[�w�B�SQ��ϯT�;�C #����	�u�`1L���w���T��u�n��s����JH���VM�
�P��HA��>��7L��\_�6u�A�k����]��R�E��p��P�����̕Ŀ~,ps�[j���̷be�~p��^�]w��sTׁ���{ޠ��D#ؖ�[�M��U[�D�þ�oe�~<�M��c��!F��p�e��'���lTǭ��8�����9-qr!Ի�ί�`T7�\`�sw6�>dT�g��}1){��f!-��!G�d����-��	�yFj���\�����d��Φ}�OU4�aS�5�VF�dl�"���F���͎ٗ
7 �~�B���~R�_�\�q�?����!�q��������R��NZ�����nv�v��u�6��||�F�;<�_�}��J���Kum�#s�P����o��Ώ������EҖ��m��F��5�0^�Z��;?�����C�4ee���^ca)a�-(����
�>��x:j�"���:�(�$�In+���2�������?����J<�5��~�_d�c���0��m�����c˹�2*U������U,AXZ�/3j�PݵIV�V������˿��z�B�=��?R�o��'�1���x��V������R�ƈ @�l �\ 9���)�ǲ����ߧ�\!�6K�Mil�<���a�d���������_�b,t����݊�����,�qqi�AN��T�:��4RWj�e[�{-c��U#Su�l
�3�߷:���@�]L:u�����_j{|�r��{IIK��K����)�А���4A2zz	e����J|��J+(PJ���w���VΊ�3�ݾ1�*���U=ˋ����~(�S��q�}���E��*��<1Da.f����M��*9e�>}J�ҕ�ș����ޝ�����c��@����ǻd�;�j�?߿NN�*].���Ƚ�%�A�\���m��d�\�k��^�O��&�G+��ׂ������F\��+������<,ƴF�]m9mL��ϝ찺�BW]7^�R�z���L�?��=&~�^�8/-+'׸�j="X���k222ߗ/_R��s�7�d�j=X���0���
����`ؚ��1W�n���nN?!�O�dl�����:�����CV�{R�׊:&\�&͝0]���Ls_�c��ܿ�3��S~5_=;5f}��Q�`����f�\�e��X�v��~���̌a,܅�]�"A���h���Ԕ\Z:��ܥ�h�S��&:۸��\{�noc�7�zC�����e�b_׏����]�#�<�L��]~XO=�a^�W��,�:��>Y	L�՘k�O�����U]j��
V#����n멌$���F�9:�|@���f��`0��������)�C���������~��e���_pkO ���,Q�>��FY>�>e������PI�h�v�u��2o�i����aVG]�a;.�CH��C�cݪ�w������*"	A@5L7�p����b�b˨��F-t3M�f�!�* ��^�	gh���pQ(��&�E5w?�����߯��K<^�4��!0�y�nO@��������x�y��yP�,�>�:�H���L
��Zia�Q��EX]���U]Jѭ�����?��ttt6v�kk��/��Od�ſt�W�B���մIϱ쵱�uO��]5��6¥�������*m�P�g�Դ>��ܧ����r���l�
�J_D��.$�ē]�=�f}W�>��연3o�QTTRRRv��2;�o�),���j��!I�����*��K���lT�^E�Ѻ䫠8�jU��um�|�,�\o��6��O�G�D �e�N旦���o���3=��(*���v�µL�j�x�_�Eʈ�en\"��G��q�������;�T��ml��zǫ׆is�B&��w��s��\f��O6K�����a�i��5UYM�(��sZa/�no�K��<�L��8Jb��l����sE�4��r�Z��#?�,�������4�5z�mvҷD�|�v��S��2���hwӊ~_����LKL��[�3�.����+]���55��>ZL[���}��R�m�5L=�ȳӎ�4�^*D�~Jl�yP`2L���W�����S����D��'3��6Q�2��\��7e��|4����J:#��E�|�^�3��6�����M"�0��6\fc���+V�YZ��c-6�V
n$Y�m����ũ�����2�����)\��l�<�1p��Xu���y*akE a'�;��l�*g�	�8I����o�.�`2�`</g:u^��M���є��+P�C+I�����7��L�:[��A\�;�%u�p3a��O)-�G�5���ا��C�0�V�$������ɏ�l�'�+� �4
�QD�m.���	A�l��e���K�ʺ���2�&��,���`��5l[q���a�\�������/#T�nb��f���kl�&Uܘ����,�f��;""gB_D޽������r�H�F��g���GH��Uk<�!��b����9�4v��-deq�e~sJ�RΚ/+��/�f��?|Χ	�����9-�^|u��5=#���Mu�\p�g���'Z+Q���R�L�?a1>�J�~/�g�^y���?"X�ҝ�.��G7,�5�d��w@.�`�E��-C��)�io�ʜ6"I⇊�b��<�Fr���b:j�O@��m����J%���y||������3�L�F��^�|���i��&����=�Ϳ���J\GM�S�0+g��V?pQ�ig�_���h���;��q80x�h�oX�|kk�q�����Enddd����fz��=��FicxZ����d�>ܲ�kέe�lC�b����� ��'��)���`�	�")����=>N9x�;z�z�]������W�T� �_�i�����������.��yg��^ݟ�'��͉k6 ��C���.,�����J�;7��闓�S��I�,�Nwc�4�4!�>m�Ld�u[�K�J�F,O]�$�
I��3�fQ#W�t���h��N�Rf�e��$I�)�����n|����:�����j�Ը:
g��8ب*p�J�a|+Ek� 34��t����6�ׯ�?]�[=%00���(�_0�����,;/ݳN~�r�H�n+���PI��1�}l��tԇ�������{
��������`��d���ה�����/�`�" _�2666�y��t��N�QBoE������W�Zw
�:�P�?�N*����0�T��Mc�uF:��Jί|h_�9�C����,�D���@�Sҁf?�Ƅ��F�7�Ya>ow�ͼ���y"ui�nt�oal쟭H��~G.���v~��h�����C�N��/	M��7ސy�п�eY�3=&������|�ĳJ,~�"�P�sz�ڇk��6���J��c�N�����:
}VM9���4�r*H�'y��}��_1��b��M�&�Y����~˰��"n}-M��3��T(�3���6���H�٢5�@�C�+*��8o�u���3ɯ>-/�Fi�_^^^t�o�GY�������z�h�^31q�,W�l�e�'b�g٪)�Y�%$Ҕܦ�����+*(¥�_�Nw�Ǿ~���jVp�+�Ib�8}���*�QR�����GE�ŏ��� ���dK4����o�7����3E��WUQ����\ooo�3���{G�����\/v5:&�|Y�]�^*Y���|u����åɠ�ak�����h����������M33��|�N�m�N7=�0�FOfl닳�V}D|��\�%+pqrz�kV�!1��n��=1A�B����¥�܁�~���$Y3;]��Y��C���As�����6�VXb㗜�����ގ��
����X����E����W�u�jY�� ",,,�ڲ������klۄr�%%�k��O�>yF;"@~���_=�� ����q�%\:��_*��o��K��/���ƴ�߿��=�ؙ�z����o�(e�::r��ӟ����)���)))t�Ԉ��Ŕ�\�����35.�>�� �~��t,�u4�ecckL��L,��>ܫE��ױ�H>U5���"� ���[�H���#�]S�@z9���9�p�bM���M�{N���S�\�9������6��ϕ���xs;;�۬����?�����-���-�U���]�g�-�H�#^����>M��C�G3�;�B��៕��E~�ڧl��D�?�����b%�5����<v�k<��5����&&&~��ʞ��vҖr�|�ׯ ӣ4����)��:\�>������ً�9	�~��C��/&&:�}kkk�����ƺ:1�o���OY��7n8�ϗ��~��̈+1v�p��&��S�K���p1��j255��@b��F?�"����#���]> �x��'�Addd8yyo�r��CFԻ���}����Qd�K�����;E���8�H��ޑё���;&�(�s�hA*���я��Ԕ��B�ٱ\[VV6��]��M�%I���+S���9ʁ|���C*aa����z�랞�� r�1:L}�=ql�����v����576h�5\z�9�E*�'
���[���ja`�����gv7�o	A�p9�X���<�h�*m�Y�0�׃�A�h��'g�M`RRd}���"��{;�%Ξ���^��j������JS"������A��bG����RQ!M��6p�cY�i9��^jlL��͛�R!E/� ��2�x��U�F���N��'�[�e����\\��[�{:.1��9Lս���Th�i��XAy�����`u$%�M�7(�[qqq?��>G�m��*pH���'�>U�Rʒ����i�sO!���63��A�ӝ:QB���U�V&,BFA�~mm�Ŵ0���h	�D�ѐ˸�(���M���W�pk�w@����NT��7~��#pp��o��3���	�gY��>zm��	�@���+Y��sq
	Q �;�m.}����n<���o��5��� s4B�>���HB�	��c��Y�VZzp
�O	���a��S_�63A]�q�B��`# �l_�r��C�o�����z�JK��ㅑɕ��Kf⅄׮A�,V�S�2ګ&���[W��t*����)}`8�{�" �����F�aF�˗/<[g�o6���!��	�6z�KN��$�Ȳ�&���Q�D�1g������� $ i���d���襢��ρd��$����N�kjZ��	>��~��G�bv�0�lP���]���0鴲�7� �*�\���oje�qg8���"\XS�'�F����kf�<�i@����._�,@Np0��`�w��U��g+m=5Fȝw+E9:��d�tw���4G���n�z��W�D;�����v<�]z��)�a ��eqL�Es��+�djY���� �Q��>a_lQς�ר���r@s���@�L���B�/u�f��)���M���EIE�"��ׁ+�|�>����%jv��0jp�_c�QUtl�(���ɍ�>�-��(R����j�����$\���A�433�p�kY�)޹Aҋ>#7.X���J����^BT��׃hd���\���ƩF��å �%��X���0���Մ�T�ٶj��'�;����s�oN�H^�oוl0��h8f�@�=::����m����ίi2jj����I���砓��Q�},&H��*��Tȷ�J�SCh��oI����] R�ӽ�u��WA�.G������9�f3v%��{Q��q�	b|�����>��n�K~-�U�r6H�)�L<�� �
���w�@�iθ�y���[�g�^�'>���`��[+(�{੕v-��@&9���� �·J��bnc��5�.7�~$���4��sb'GO�*k� ��_~����5BAP�7q�s�'��#��{�>������mB���*�4.*���Ċ�_��7[
H�<v��k�_��B>~������`;$�M����u��R���UmYY���`����Q@ �;�3Ȕ1W$�����N�����޴&���~�@�99��; ��uƿ����E|��i�<���׿����z�Z0��� �Č�t����͙
���^t
?��p|�X>i��x��ѕ��0(�l���i�TV|�5���c��>C�]��dR!<�
�A꺺�gI��v�4;tk>"YFs�҂�~���wڹ�����1�a<�D�	��\�̪*����_K1㕃e��}It������r�>��w:4�����Q�K� ��]�FVnW`Yly���f����;��\�?�J������.��7���OЀ?�~�O����G��N*Y٢T֠���W��B��P�[���OБz�����M�� Xp{ХN[�꪿��k�x�Ĝ<<7+]0�?��s57�ΟP�y����*i���GS���D<��:`%	��QRZ�$�qL��!�p��;���u���]�(d�F����:g��ěPut�!2�&��3�n@�N�=�{��.�������l�b�I&)���m�sr���P8�$ZYY$����!O
�H�(@y M��g�V��F%�G�a��,;I#�C�bN7SeDó�vbp�U/������I��w��V��"Em-��K� �G����L�ݴ��b�?������\Q<�7��-���m]8.	�⯧�|�p��K{_����\Z\���R��V�Ύ+�G�j�cS	�����)8�<��9��6{6ZB�+"_F���m[��ek�n+e����'�����һ�J��X�c�j�� b�Eƿ��V�� ��0�}q@�$ص)G��3pu��ǧx�!q���A^>)j���pv����O���l3֣�� �JtE�4�y!7ܹH�~-��?�B��yu@LN�!yz�Z��;�cV�����:F���P�t�u�IO�r�{�����B��g٪�^����*}�Vc.�_S�-󎄢+___��!(~�Z���;�94S��'>�K��O@(�C�����'�/@N6ttȾ�`]T$>>:��j� �j
@��KU���=��p����`�g�p,h]6H�t6����6:@W���$~����^\�8���+\X\���S؊F
a����T��]��4Ֆ��gA��LZ����ozz��8zcdX)��/ � `[�E���P�qP]�իW���ssr����M���~�4m6a�4���Q�~i'�t�uB �Y z���]� l�Yk�X�ѣ��s5�����ٙf����3`v#�?8�j�z{{����.��
e�  @�y�f�=�3��N�e���A �y���y(��.���?o���0d����M󽏏�6:� ��nYL�W ���`� ���XX�0��pV(�>;f��"�pI��{�w�#(����t������HB�Q�e����?H������p����l@�qm�0���<y23V�BN�T3�	� f��H�7��р��0]9"I��(�Z���������\iU�A�3S�| 6��!�%�0Hb@$LVʔ(����xzoYm��B��A����# ������v�*{��#�Ė���+�K��JV?�<T��4p��]'��!d������ jM	�3 �E�>��#�Q�5?=���}���uǳ3_$�1�Ùå9��9����o8���rx��$-��05�mK#�0"2��As�݊�5��e �L�q�~= v�N�=����e*}IYY� #=0W vH	�����oZ�Z��	�g�UB�-WX� 2s++8�T4H�oD���O\�1�vzR� �1�/������-.)�P��Tw�"6P�\X�}֕3�+כ)))������h`~'~�شB�"�j<HuE�>	���5����@|�m���������/��_�����D���x�� 9Ъ�??�=e�zNNNh�Pu���/㢑}8�&?d�)8FN�qW����x�"��&?<<<F}���LI�G����� �Ƚ	N�X{��1
�|#�T�=AN.u���q8���(e���� �I����ߎ��
���'�Gh��l4�8�;u����Up�'�H��9D��?��@���O��!�����;�2��P���A��Q>��5�s]*R!�����@ �{�2,B6���V������d ] ?��}>���j�nR�9��ܓ4��|�'Tq7�UB2�m!���v�D5b���^���w�lq�����~U7�G1E����jMa��S��wf��JU�k�M����
T�:Ju��V�e.���?g�\<�D��E���,RhXNL��H�@5��������dX��o�?�|>;��oƚe���>Ig�Y-����$%L����oG�kC�4����h�o)�]J�kw�.�P������Z�D��BK��"�IgC�bN���Q5�4R�(,�֊z-�b޹x�W;x-(�XĘN֩,FV��=�#�`h�^n���1׺K���6�m�=�[�LpU��ƷE����o [_���%#��}Z����x&��֯O[����]�/f���tI�Gc�3q��ލ�؉��M��Q;ݤ�|5������~|�cG�:�k+zǯ��5ۗ;-j�R��-��i�_��NArzeu��s0��{hҪ}~��s�����#�eI/���L����+�)W{C�x�D�&����VOG��z�h�����	m��ե �%b�����z��$�3�u�1��0�DC�}@-z{0��m�[��O�تt��>��������]�x�P=�����Q�i �z7rT���9�7�%��w���R����yRk������u1����~��T�x�`����� 1��ÆB HVaI;��c�e�붱1�t(��Ӧ���������\���%/�7��[�������b����=�[Y^~���P�8��QBO���ڃn��XĊ�~.��tŸ+�oY����6s�moo��=��=v��8 ��� d���\U饔�[��������$6�ik�gf/�v���
�Z����������˱\{s�6ۅ6d	-`�gf�������+Ǔ�u�\�O�F5�v]�ܪ�r@��������y��t"Da�\��=]j�p�@��5nr�*l��@bt�p�(��?��C=�ֽ���{[�E����N���G����j�)S�>�^��K&�d�W�"Iff]�_��`kЗ�+�_4�f(e7ez�9:کm���T�������{�e!%����}s �o���\���Sz���B�f&=�bf�kw�@��?vЪ���%��M��A�Ӏ����*���At�q����j;�g��E=o����E۟F��kׂ]��h����An(I�����@����o؇����%�klH;;�&�Fڣ����tnlH@|��2UΒD"�z��C;����'ڟ�%B�vk��r�����q_֬�Ȏ� U�h_�ՌY6�n���@n��hv��7��M�p/���H͐*������$�0�C{�JM�j�M�����_��m�+�Θ6K�����5�ބj��HR�>ĞaՁ����5�a��h�0W#�F�v�FG)��9���`rz�U�m�&D$��s(���[�q�$f�|y�(.)�e�+l�*����c����ît�ÞKGHL��z4f�~ѻ!������srv~�#'��%dk9���j�!{�~�����u�[n�?:W��r��� o�	�n��c�'����ǈ��
w�l����|����	@�ѐ!��KU=�}����uϯ]Ci�ny#7��h$X3����hVcv搳�	RᡠjL���L���L)�ܞ���� ����8���>d�Y_����C]x>{���h�6�Z�`7�M1G�6�L�y���S	G{�h,t�)4u���!�TSS����ǂ "0�2+,��i�T�7�5���7�)�+���*�L��F����l�ˁ����6�'f�V�8�)���$4L];�e�n��-� 0>8�9���K�z!�eu�}���H����q͹�A�R��Eg�)��Uq~��7�}'S����OL,q�1.����i��qV��#��/jl��3�J8~��=͸�����J��ᗤ[[��X�u@��5�o����m���}W��H/�1�/�5�ޫ�ܴ��.q4���:T�u����,�xQ����}����d�O ޥ���.k�w$�z���<G@G�L4Z�%���� 
'�>O���%
�GYK�˚��_?Oo��1��I��V�"��Pf��~�^�ڞ�^���є�7�Y_�'�c����\j��&��җ�E��e}~̿�=��{��%���D)�������&T��C8)�P�n�<�HL��X[�=�k�K"r @߀iJl�v�mq���<Q��e����?�A
���j��s�[Y*Y˲�A"��g�IR?Ǒ�>��8��8l8�)a�i��,fx�@PtR �Low�����M��Cl���+��I������Y�!� �JZ�|E.�c�/���N�1j���va3�J|+57�2ߞc3���ز�q�%�}pv���7��j��Z|k�fM�������c+�c�;;[���RO��b�,� <[���	�L��Ų�����mD*<�p�c����+�ȑT�s�H�R� z��s��������𮂊�����B�͊-w�G[�Q���B�#~����IVSI{����͓h�A
|/[�������s�'o�&��vm�{��E��F)�7~֠[;���+�:�-���&���t4?�lk��p��`M�L��~~2�&���̖k� ��qC4�<�Ѭ�n����V��p;!�f�6���_���=k�	IIIHR�~'%�<��5F*?^����b�����ir�{d���q	ѱ�%�)�B�^f��W�`w71v0
\M�c�s� �1Ķ���-Q��0�hrrSX���'�E����qU��SF�D�+Y�_���'�b���{�h��$�jƊ����&��1;7�	�#�@�-Dc��oK&zG��
��PS� C2�����4�ʍ��D�K�VG��OCR��=F�N^��`�B-���B��������8�X+0,333 j��������S֌��?�����
O��4:n�M�Zl)!q��3��N�&�<���]�f��4iM:z�v�׏�h-]���^��z��Q�N(f'��t�h���NK�D���XS��}m��T����.�|�nm���j}*�II�1��Z=+�1��5�_/�����"��-�b��v������M��$������jX��.
���o}���m�CLc�<�V=�u`:�ںjs*0n��GO=��Gg;Zo�L(/mD��q�k�ۥo��	Ōn��(�r���ʽ����7�{��碳��?�9�ϥ�Pz�6�8��������#�:d�'���T-�)�*DU�P�̱�<GAO�f�.=콟9����s��լvwA�H���6�Xu]��6�F�J� :�(r3�rk�y�w|����I/��me��f��s����C��9���#Z�IL���I�;��r1Mj�� ����8X^�N�ޱ(Km����}��P�n)��mz�sV��w���U��y�Sa��Ϣ?׮���,9���-�/���t��S�VYe[�Ń�:g�{�cQH��R�����C�m�3�ۥe���KL&{>��(��q�픪s�;��U��n�Ţ8	�tk	6��of��{?����h-��؊���j��QMp��g@W�K����	�p�e�E�
ͽ1zz)G�v�$5�'��� ��-��d�,%��?�m�D�D^&�s�e n�iZ�˂��x���I�(��;QsD2)�Yq��ͭ���'�
�D��|�~�h[���kL.`�`��uf��}���}?k=�2�ܦ׍�'mєG2G��
s�Ǜ�R�=���<Q&=/�۹7WE���^���&
��ri�ݯ$Bq(^�����F������*���l2�[j��Iy�|	�bU|��q�E%ܢ�9IS�
k� ��$�r��<w��������8"Mm<~c�b����Xg{m�Y�����z�H�I�Q��G���f���	��³w3���iIH�xm��y���伂
�W�?(i���G^Q�d���+�}��P��>�*G�O���[\��~)J@#­�������(}$Ad���U���&W�tQ�]��G3���}�������z@TB����",���6�`��Tj�L���笄I99�.E���y6z<�8���^�q�#>��[�9"4���0'�óck��l����b)rB/%�}�L]wF7�F�9�QL=�����_p�tn:�ˬ��S��`L������]y����>����YWA�q��lS	)�u�o%YFqy��Lz5+�I��_�	��9��&7l��!V��6#��7.�b<W$�U�����M�o߿��`�<U+���/����h���H�QeV�h�[��������!�A�s)�>Z�
?��j��t�d�XzC^|��[]Ʒ��Z��3~j�lx�s�\��۝֠m���Pf�E�c���\�c�QP��`���.����K#�x�5���%� j\)�z��U����a��:��i��H9݄���g�sH����:q	�5�7���3�����{��*#�gG4`�� N�XS��
dZ�gy��Mu�U����VH�i�2��̍����"�m�dnv�����
�qp�<�D#��g聈Kb��:�	8��?=Ikilt���ȹ���6������Ԡ9�	Jm���HDy�W�R,HB���0~��r���,UAe͡O,n=���#��*wv��ԏ'{��t�b���z���3E{c8H�@��N<ჸ��=���x;nPZ���u�����J5�TI�I��p�aT6�i��¹��Y����O��֣"�{}[�}�>I ���A >�j0��2ģʢHE����bn�h��0���3Z���]�y{n`�[[�X3J���������ZK�[yp�S8��W���c�!�d���ݶSO<��*N X�Y^���i݅���
q�B݇�d9#�"�I�d��Q�u�d�j����Z�v�#�nQ�b�Ŭ�U���	��_�	��/����4������`�}��/v�,�]T�ik�nJ�#��+�ƋJ��H�>��Ӕo�Sέ���=~��O�p�H0��ll�8���u���G�W�2��&���u&k�Jh6�C��v/��������y��:j�?~�ϵ70�qw�j��_̎� s�Z�a!����c{�6��h��\�'i"^�5��˜�
�^�do��"m�1�^z�ax���a:4A���7G�O{o��|0��G"X�����X� ��+$:2-?d�[j�+4���n�Dy`��_1z�-ҺTx��c[ݔ�C�y^}��#��r��9��9��l�[���o\:�����v+�y��KE ������]LQ��Bּx ]Z�l��9�; �1E���&P��H�;`E����o�&�#�ݜ,�������c�l�W��|��}�I�e�6B{=����Hf�$��&��휘w���#�Hi{Eun���ư�^t�(��԰���KK�k�԰��C��^c�5h�ݛ^G/?�(�#洿�蔡��*��5P��`$c�[-m�۶!�y�\"�����X��>p��%h�#譞L,f�]���`���^u����������j���]�%U��!����sƔZ#��^��7UZJ�u��L4�p��T�b�]�SO�pcU�[���L!`�@����QZ����Z9*���uX2��]���o/��E�Cw��L�����>�{�:��R�@:��E�`i>GXIʆ�Ҙ��`�o��+�4:Ô�_3�5g���?u��������й��E~�s,���hN��+��8�j�7b�y\}����r�5+�%�T�O;���RA.�#�����B*l���S,�w ����X�wy+0c�#5T�C�m��ƾc���Aa伄�|�������g�º���Rp@$��������/�Dϭ2`u�3Q�a�+�<l�.�x����������=�IÈ�J]?åG믧g�}7���]+�=l��_�x�>��{zd|�����+��+��g=��F\V2q�Λ��@�6v*��+���Q����z~0�i��)잁��m=�&)��)�X�������^C�g���n|@��\OvϯG�]�r��Xh��a�D9������=��hhj'�E��^�3��pMІuRr�@�UxB�æ(�COɘ=c�A�s����"�"��k��y&��wv�6�8_+�?���ߡa�	�Ez�� q%}�&)�ӧ_���!*�(~�xh݊��47�<闁�ϟS����p����*����	ˆW���S���ёm�}0�w�\X��V�|�gM�+)6T'\�p��)���������a�O!�d����tS7� mT|~��#z0B�@|�+��<{����O>��Ͻ
7u�
�}k��#�U�n�v�/�7Of��:̕Zo��f�b�}�������P��Z�䝒�]{k4���`IA�� ��z>R���};��[B�7�aN�IA\�j~j:�(Ց�jJ�n:��v�CC�	+�Q��76�Z8��&$]Q8���z ݑ~mˤg?$��{z(�'j�o��Nmd�5>y8�B���-��"-ک�'�m�2v�����ؼGh��/�_�W�"Q0܉�=����@c�P�?�9�74=��SO��f�����]�L�ޣ����@"�V���1�J:���+?0/��8�/�[�ܧ�O{o�{5�^����O���$(���8��\2cxu������yQ��$��2��
-!�#A�^�)�S�������sǭU�4���xd����G[R�RUp��O���+/��6��;���u��|q(�MYE�GpC�qP�Q��9J�U�;<�02��J�TU��#�ǘ\�L�}�dqȿ��	�Ȋ)�V�y*)t�A>#�F#O�4��a۱5[e�[:moǽ���|){�@�w��i.fgZ�;/�^w|K*���.�:���8γ�RI�]�����w������.��{��Y_H�:��[�*�%~�(vy�=��2�u��j�e���-^!��Z��%��6���{�����u'e2�F�F���Ā� K�sݮmIk�ˊ[sa���k�p��*�6�m�t	����8؉���h����T3��mc��|�g԰u�$p7�9�n���)���S_n��ʱȅ*�����'4t��:����ò5�#K �����
�JPԴe�x�Y�����؀��r
�*Ļ>���˹�--�����5�\{�f��Q1յ�\�I��Z���}v�5����D����K�&V���+]B'����m�Q��1�B�\�;�A���_���,P�7�'�!�q�`L^��`��a�ZE��U;BNU�`��ff'���S�{�FC��{3�tWbl��Vx�Y��^����x�'-d����@���R]���5%5,�a�Q�}�la=��ۓ��w��Ze�<B	4��7��L����'�ٱ�%��퇵�|��Y�c`����uq��~:R9?܂{7�:[7�;b�{�9Ɵ�L���\1Tx
"m��v�u"'��zޫ� �.4�����z@p�s��;uA�;���
4�>����N��������׺��qs���7��BNb�n��j�sI�����?�e�xX0dL��5�ͻB"6͵�m၊M_m�jU��^��&
zж3*C���j�k�u���_N�M<{>Xf����ͱ@�*$�������ɬ�Z�X�k_�z�]�����5]y�+IUi�:D�K�=
R�'���h�O7>��+����/���sU��
����1�W�^�U�7hg���_�J,YBo�Dd������!��mX17��MuDW�.�O�S�/�����?{Cv����*�s��m��4��?���fZ"���N3�2�:G����+!����2v7�8��J���>	��%�g��B�^i�\�~��fŸqo�o����gW�ɽ��j�ωt.�-\~��V�[FyѶ��ho��N�k�[�o���I�<7V�B=��v�	G�v����_�o����S�!�_y��U��� ����S2r�b;���W�M;�_ˌLn��C&�IW��mw&Z��ϵ��4�C=�!��J�\��E���C���Mo����p>�}p����'���7��BD�:��Z�������2����{3��hܩ�GM�fX?�s�R�%]Be��߷��kr��"�Ll��GNVz��Xk��N=.�4���'�rh]�\)V#�Y��k�����\��[/�l����$�7��>]	%/�ڊ�e�jg7����N�4��\3<���]C� GM��<�ͯUe�D:��Z�����&I8��%[nUm�ƿ߫��f*H2K�{�8$SK�ߪ������?:i���^�W��b�j�e�qd%�鞵�H���~	�C׷c����M��v���x�A"[K�Z������ɽ��R��u�T�Ӟb��J��*�μf��k!a�}�M˻��S������p���vF�n��J�[�5�����>����!�VOO�D�֮���Qm��6]�����Zd�.QpJw�����$v-���F��ˎ�\r��t�7{�zZ��z^*�R|�ט2:��5��9vd�N�z�>�Sm�3תt�	W�Aٿ�7��Y�6�0F8����Vk	�����O�DH���]���7��1�������.�A������+2���*�7�P��ގO�ꜚ�h�Y�ֵS���F���<Q`sO�`n�-�I����/��V˨�?���z��?��s�X��A':�/�Zk@�U�Zߣ`YZ֝��e�7��[�U��,��JI1�{�9�Q��)�^����Sn�펍���$��/A	��L�w6	ɬ��Xx`+Z�Ǯ�ޘ��`_�͐>�q�?��^��P���S��!��C�K���&�$�薊��=���WH�4��8O-QZ�H��,��z���^c}�C;T���󊫈?ܷ�f��V���#*B)U�52�c���1�g�-��g5>�7?����{�tt�^(�;�1�%�1���鐷�Zҍ�~��H����:#H���GGu�Ũ�����E�~�MU��{`���63�Ar{���n���n�z>^��v�^���)����	<�a���ݑ�q����ž���~�L�;�Ą�`r'�hHw`�v�C��]�yiXtxi�����s4$o���V�������Ki���V�VǶ�.S�w��Z�e��.��`j��g�I0�$a�o�NV}w<\g�-my#<R���r��~̀�����j�4�w��UlS�oWL�J��&?���\`x8�g^���t��r�⤜!������j%��h�@w2(�F�J�9��MSV[/5���5Q����A���9��������[��UH��zZ��1���Ⱥ�&����DiOi�ҥ�bA��ҋ��� `�J�EiB��@��ޤFB�bH�	%����S?��x8�ν3w�73ww��u �zǱ�1D�Y�N�Us)��`�m��=v�����[n���"���&?-j��Vh��	�*�<W~�<��?\�4�@��X�W}��r*���F�S�������%LYr� �f�ȸ�3L������.��2��	1揍�������e��Q�.�����)�m���qhӾ��y��fV���*cm?�����$p���8ʩ��n�i�o(�5M#{'�0I�T���#Jo����U�������(�z^nPY�L����Du��[�a|�?�:ĳ�,��r�$=X˝�6֖�p�mT�ɟ�S$J5J�P���ޜ��ѩ��4��cL2�P���q�[�s����h�>c��r	����������#��������UW�+V��;�"�M(�7�<�1���X�|p&O�c꽼��a��������/����,�Nmۉc���R����F��	�_#'�m�Q��yѺ����;KM�����W^vtɎ�H�9���"����Џ���{A3P7�}�W�R=���H�/�c�ޏ��vp�1N�G��yW��ۚ� #�E�Հ.�kS��'<�#ɋ��L%�~��t u�)��>4[��賿&��$e��#�v��`���&1]X_�e�;ѫ� �S���.=�>�ZɳLV)���z�!��<+l���t��|)d�)]mՐ�
s����m�`�u&\�j�q��3�R}��;��ѧ#�D�#�2���j�cA&�}���i	j�14h�}{�|�Y�0d�	?,���G5Mnƒǒ�M���\3|�Q��X������ܙ�?.����MY�|; �� �o?�;E���$��ќ$�}�0$WS������'��H����e�޲2������5���q���)�ma�x����8x�E,�A�/�a�"�����V�"l��B��L�'�P��p]�U:�GI/���N�U�`���x�-'�Ӻh���GGz~�=X�a}�J���� ��аo0�O/@�*P\1=��pu����}�i�: eӺY�{;�����@��V�H��&oK�MY�9巂󬒻�O���A���骉,k��x/I^R�������i�L��m,�g�;���&��B*!�
	-ͦF���ը�x+I���	 2��-b����4�U�ᄹY8�l��&��Ĭ��?ulw�p�f�Z`-�(	��|���Sq��!+y. ��rt`$i���$��JG,'���p�1\�~��cIY�����&��G�^~5!z(������7��8�&�88؝��,p>�p���CV����ek��Ks��$�mH�m�@���!� ��:px�MBl�{�Ա)[���׶T�=�񟉝/Y'K?��� #����U�f^,�d>���+���f��V�1�����U��B�����4����)���z+|��x��crN�����"�'�������i�T��_�7��������!���W���������ݞv�5�r�Oώ&k�g�Mp��Լ��)$�-��f�d�=����{_��$t��5�̬�w�e(�k)������I#�����]w�,����.]1� }8Pn�B���#�;��
4BpM���=��C( A��A�>���� �)#Q6w�Ք��O�H��,����Z�Her�ʈM��GS��� ��&��y�8K�>�����glu]�Nc�1�י�TGk��V�DD��wPIL�%�G���p3;/IRj�cIxu�*��iu}���k@����8��B�����K	K������dZ�"]ԕF�L�>ߥP�����gc��@Ѷuha��?8O~�_W�<��,k���J
�o��������̊n��T�ɛQu�̸Ք�����6��Jd��=D����R1���~��H�����C9$-W-P�J��B�D���V�B��4_�I�Y,�e����_I�`�I�}�|K�7?3�藄0g�����KQZ��Ő�~���� ��z�E�%\-���_60S�4A\����zwf�\�wA.]�-��:Ghnڎ�36��#	�=��{�w���� Y��:O��;��sjӓ�чr�B��=đ��K��7�AU��Eoi�,��{,:�4�_��
O��.��i�s����	b��Ey��M�?),ˏ�h}�^M�v|�s�;y$G���,���-����1��c6@"�6r3���f"_p�=�n����C~3�v����?��m�_O֮jrsS.Tm���Av�j{�< ����M�^�3[�9hi���Kn�Є����#��"�L#��I�nmE��};wϻu7�v1'ϵ|B}�L�e���m����ȯRg�2,��&�Wƺ��͟����[d�A��	�9 Td�F=4����j�:��ma��߳%1����ܐ`յ���
�,���9`��pm��>�DW�I�Dо�V� X:��O�GɁ����������e*�:�&�A,Ca>f�\fKJ}�w�~%��8��\@�W��U��$�U]c���_Yۀ�N�̅X��x6eU d��*��A�T��ٟ�W��Y�\5x�Gn&j�S��p̶p�1I�O.�]y��L��]� O�z�<�X���<�|�� _�*�� �F?�y���5��F�6�LM ��=�����~�Ќb�!�_g3���n,>�D~���(�J7)�zz��q*��q�fTkV/�z��k	��q�TfY�k�j�]!>������3���;��_�("�4 ��{|�j�x\�eQF0"l�z��Q�M9oJt�����RM���F�j�\��]�Pf{q�rS�e�ͥ�:�w�\ߪ��u�Ў#*��
��iċ�:�й�k��'h*�� m3�E�~k����
��W35�v&��ՠ��tS��5xuY
��LB��s;W��~r�bsn�*��	��)�u򚒪]����Ɵ40<={��2w���D�Dи�r�a j� �b����9Bl�
B�N� ��Vz0���D�O���J�-d�-nz���z�C�/3�b}��},F�{](�m�ȍr�͠��&$=��]���1o"�C(��μ.��	c�/r�ǚg����yVY-�9�Ǝ���5]6�|.��	�]���^�LqAq_��LW�ӹ?�=�V׶�q�o[��MUE�SV(ࡩ梪ôcxwqKȒ��D!r�7��n΢�Xݛn\ǖx�b Lo� �ޒ��]^���t��������Q��T%����߂LU-q_��2�����z�<�V���R8k]�J7 ��8i����ΡN㱚Bgc�ܻq��߿��癟�x0P��p*������5rn��c���J�����5Q. @ ���f�6����3^��<�hBR��d0�Z�#���et������]���G���DA���qn�6����{�!��ަ�(��n6��q�^D��B,KꂡC���ԬQWv��`1��a��'�!�ِZÎ׿���aj�3��]���r 3�7�>xo��k�U��#���s[���D�\�	�QK���~��t�P^i����d����:a��.Y�]đ�6�h'T�����߂�#������$�I6���xs/��O��7��@W�WR�{=�@�2��lz�� !��}Z��q��Q�#V-)���D倨��!���$�sȹl){�$fw?����� ^} O��䫁���ī(ҕ�0˙��ܧq�I1�Ǵ!���2lLU�h�qI�v���v�T/�=�]V�I*�,�X m�k��'����F�tƠ˝ӣ�B�Y�8�)�^����l��Lm����U���� �ء��B�dZ`L��*�g֘�Y�BK����e�C�:�+�e2W��
��-R�&<.)Y�	��Ȫ��A���DP՟H�:�52<Z�0xm$n��W�\���������G��l	�UVN|l�E(��9`�����Cg�H�d��.'7�<J7R|o����+g�~�*���ׂ�-��e9ЬJH�b��R�!��Ǔ�I2�^�C��RK�o��b�蜚��=��gј~@��y�_qg�
d���|Yl�9����z���n�՝qݧ� ��ӷ�1̜�v滝А�YJ�P_�	'ip��G�o�qo�P��蚶:��{#M1Կd/�uG6�}��fQ�����J&�_����rD��%��"d�f�ӣo^,���7�i!}��h���_��F�Rԃ&�V��[�M���nt#���yLfе�d1㖃/�[;�(/0(e
D��|�Fv��V�o�����l���U_൴kq��zF�Z���� ׎C�	ږ����Y��ü�]:�a���[� =��|\���.���'8�mm�h�U���y��`P�Z�{^������6�����;�:H����濪/$J)�+��Hsđ��+��=��3�|^]>:ﵪs�A��7Ϩ~�����N��a�H\U�A;���8�͕��������щ�/X_�j����ٔ:���oNi��A�@��gmt7��"P4���.�jtU�/I��~��+�{_/��K��4]�}e��~��X`���2�o�Q}'$���48��ax��Q8��^ƞt�Vn�50�[@����]U�џz�/���͂{��TB�͹Ǡ��.W�]AZ�8��p�ąLJU���9r�.�r�ii(j��7@'�(��T ��]�2���ǿ'AG�ٺ��Tp�H-Б+̵��呕լ/ͫ9��$��rĆʒjPx��q���Q-���ݹ����]�#�����JK-���x��:���~�OW�e����E�!��NFN��A>�Gm�)I�S����.�zhK}.�ud�j}��گ�����s���1O�1-M�٨#��_f�)c&~���,�ϧ���A�*4b�V�@H�ĩ��@(.katW2q/B��˯�M\�I4z�T�4j6�6.�=��a��!e#X�3����0-�N�~�P�_�D���i��7�^aS���>�R��I��o��JZա��~1K'�o��.}Q���n0W�ee����z�yw��U�<l����SC��#0���j{��ݼ�Z���q�~O��^7����5���t�}5�b��c�@%��uy�4�}�h�o�1���90j��!hc���J8�2���ї��W�Es��G��s�P�xG�[J�U9�Ү�H�'
V^�2�q[�U�l��h4{����$pp2��D;WK�4�J��m>9�~��/�V��XE��7C�hk,S*�M�z�]A%�4�����^�f�1[�}F7���ȇ��}����}�?�}d�s��~���{p�Q�q�-�}�z�AveВ�4�#| ��ӽ�}�o.�ұN�s��Śf�
�O��Vi���Tl�����:q��tS�;�ٔAsa��o�; ;�q�^ �4�h�����9���;5�A�~�$׆���Q@��:bs��Y���ׯW��w�b�-<���������>����<��r���"w�oCx����y���<�2��`�$;	hk���L���:�q���*8��p�LlLo�@�A�8����Ep�Zpl�a����!�A,�]#�Am�ă`C�����='�w��x��8�yZC˜���;L��p��~�1&o����)ov��������0/�<��NB�pQE<V4Ѷj�~m�m�=#�!���h�{��E�2"���A�<n�KW��9�5<��'�ǻQ\M��l���o	��T�ȥ�WiV@��>�?�rT�	�ZP��C2�|�����5�����i�����F)z��V�X��RU�\�tCS��5����\�1&�~e\�d||cF�n�ͻ��)�d�����b8�u�&�n ����5�Ԟ�Q�e�X�!o��$%�ѥ�w�ޑm��Ȍp�����쬓�S�ɸ���||�h�ag���	�v�^N纭�2 ��Q6�令��+l����M��]�v>9�fxz�نChN����\<���?�!0s�z�o��P��L�Ɗ��#���j�9l-���/����)����F_���n߹1���\���i�>s,�ܝ����2̾PFZ��VH�x�8�xT��'2��0�C��Pބ�Y�U���/Or:o�X�����EY����+l��n�~f��I��R�K~yA�Q�(_�֩�h�@���qoCW���i�� kw�K��� 4���O׋Kt���9kO
xo��W(�'2s'q����P��iO<�0R���*E}�WL�e�k;����s�||�uܿ{&A7���.��9O��4��%i<0��
���m������[��a襸j%�K�1��Q�>�PYhcU����ԡ�J!��uW�e7�W�0�;�LՁu��6d�&|i�[�	c�ǌ������x���8>[��]���GkƯw7�c�j+	}f_v6�̯��@�g�_پ�*���V	�� LE��{^�Y�5��Ƴ��mt���^e�Uu�4o����;:�QpÅ������g1�՘4ʢ�ȩ�ҏ�H��m���ҢsT�`ĩ��6�I&�3��+X�l	A�,Hۍ&f���o�Y¯p[�=$E��;����q1��*��Y��3ͻï̝��uF3�'7F+���@O�"�o��;�PsR��ٯ�.�5�:�;`�jq��O�f�\��3A�5R�n���|ś4���g�}`��wZ�.Mɘ�u����*0�pJ�En<����`�o��6��p������SZ8���Zh����8Vo�QXm���:��o)�}�siTB/�K���������Lo�U�\ǎ+�1ѧ��/fM�suo���C�y�Z�)%�}
�fk���WKc���y@�A���m��m���W9[��]}���|R�cuv��ިx5H`��,�|�����h9&\�O4�?��d�/c�,vR�ޫgr��m�����t���a�?{Cꐎw5p�h�+��$Qt�6��1����^PXX�u#=��nx�� �H�)]�O�|�91�J��˗J���U���]�e�?�8X���=��X~��ʮ��F�������������m�XnI�n!,m���Śk8ƺ{��%N�3��7��N�N!��7q�&o�	���6��>%U�����c��gQnh{(�֑�s�aw��q�Xix4��i�{۱����3��_#J.r�N�J��ￒ5wK/^q�ZV<q�A���1��4F��w�xY��I��zy ���n~~�b8�nJl[��k�H�W�[NA��erd+7Q�������4K�n�/=�xV�3mV��Qq�}������
�73��%Ť�ry`J�&������5��S7q���e
��2n�fyN8�4�8x77��ѡ�w�
�6"����|�zR�ⵏ�<�s�+�Q��^�����'|���隵�?X�o&|���YX&��x긃(�<��� ���a���VC}�S{�Ii�yߵ�M�]"J����^�u�v?EA��T��\�$�n����:;���wO���ox\f� p�ڄ��U����e�Ԃx�m���?l����������>���o!�z�R�q�0�T��aUqT�:+N�uQ�f�t�݁��u�Y>=��A�`�]�պ�:#��Ǻw��&�b���RH��0�_�)���q4�1���p ]�}nRޥj>�[��x�K:D�u ��F�H����+\O�!:?�[ȼ�a������J�u�P�Q~�Cc؈�ѱ��gBN���Y)�ڡ.6��QC�UU�V�����i�r�5��{`�!ڌ%����*�������|��v�h��1�͌	�a����`�'٥jF�z�8����g�ui��,���xx��nz/ؠ��Lܰn_�g4��)%X��e�	#��"�Fju#��ŵ���y�]&"������Y��� �r����y��Z�##h�$qss:c�]r�C�f��vMtZj=��Tc4�gxߦO�]9��Yyq�����JI�踡�����&S��mOii	��S[j�Cr��ؠ�Z٦�����b����J��'� �/��>&RD\Fla��R7��O��N�w阰&¦ �3����$�SL1��S��Ix�����q�É|�ˢ��r���n��e��/��XY��/��!�7�jxI[2���a}����)��^{�5�XE�81b��c@y��/�T�s�"[�CI��_�<+
��0�O��&�t��615�d<QF:��md�������p��c�~�3�~u�{yp�u��7��B����]N����H\�n��_���P�}�piBx�8f1�BT'^ac��^Y��i��/(�N��1�1S8�f��vq2�t�S0��2Tx�p�x��R|f9T� {O]Ҭ�m7X���G��;7����v��KJ��
h��\\_!>�b1Oҽ���ZX��6F#�GT�wc�u�ܸ������f�)2|�[�PȞ���_��6����}����c�Io��_ �AI���i�]��&��U��jB�%^�z9��{���m[	Q���h�j/E�2maS��h��F#F�)�.[�qjrg��嶐ܷ,.�K�J�h�8j@�OMz�S�������GC�����.��كc� nP�Fĕ� ��p��'��1M���w��U2�wMK�:g�I��8݇���ǣ�{��}�����*�kX� �s�;=.���|w󣫱ǚ9���R2����!�*�&r�y2���i��
�M.=�D�-+�%u�M�M����k D�O�-��k��"Uʫ��Xp�`�u���ʸ =�q��U-����B�� �Q��\����^������lE|�
b�n ��Ӱ�Jڛ��9�h�Ӑ<�l[��b��k35+6��i�I
����X����G3o��(½q�=��}��s)N9����ު���:}�=��2g���ׯs���ְ��rVoXXح"���垟G�4� ��F��Ep(T�~Q{<�,{@wR��%UA���2n6� ��2FD�n9nw�)��7�,uJb�U�b����ä��"�j�0ʉ��l��v]n�������dgz{i��\�ç�T6�3�v��ґ6�;vT�U�o��_ hD/;m��j��?��^JyV��Wi���*q���Q���j`�g����c�
�Vk9�kv�������Jd����P7l�3���x�놐;�մ�x9B3�"�U���j��ˈ�-&� KOlrҰ���A��T�s��y�<PuϱT��"�櫾;z$ʁ�'�;(��h�Lo��b��#��S��t�U��%a[Y�\�2�A�j�����6-t �vr	9��D�#έJ78��R���܎9���0�K�����f�s�C�J�ѵ�CR-���:�iG�mmn��v*#�7�9��FB95�ћ��př��뵙�K˚8��2�0��չ.*��]elɏ��\x��b��#�%�B�fr+Zg�q�����o���iY�	�!4��z![��§�xL̸ωn��2�%1��2'9�t�,��!�&�I4��7��\������k���EC��qP�]�M\	xǆ"�ګhs_c�1:��X���L�.˗�T����W�ȝt6q�R�So��#�8;m���汑D��g�����Eok�l�m~KS�N�q[xr�f�k�".�cm�;ó5.$������������m��3��d�Dh�TL�?���|�W�d��%���5���8}Fs�mL��@k����O�ҾoW���(�ʵWa`m�;��e
�ћ�{����i�6�p�P�����q{?�/�y�U��f�xgў��O�LD��A�j�M���:U���+�PUIc��8������#�!R΂��cN$S%����M��Did�V��8:����ns�R�xĳ�AT1m?�)x�+�^�C�z��ǡPwh��ǅ���F�9��{?��~�!�d�U�����)��6��p��A�@w�k��u�z�T'J.����k��W;�<�y�]�6�+���~M*/O��|��m��π�����\�2Co�h���:9k!��;�I�V���ou�Q{Sq��|���۰�4pȀ Ug����y)bR�j�:הQ<E�|f2���d7À�z5��Z�a�k��| 7���!���&yN���^��?�t�5}@�ԋ�X�~��"K%���eܧ����2K�Ճ����-�4��0iRxru5��dS^��y����2mG��]���	T<A�������A�3$�����*�]Q����~hcWx-e*aJ�cB.|�.X�F$I�4��]wÊ�xT>5��Y�gMBI~�)����� ��~{	��@�ywz�c�h���:�<a Va�x���������h�M�����+���z]J��O0{��h	�����M>��S� �0���M���X�X�X�u~�C���7^�v�D�-J8������@���)'l��é�w�It1��BmM�8	� ��Q������ZNL|U�U0IEih�Kv6�v��dR��o�{N����ƃk���^��6Sݙd5yD ��v£6O\
�k�M�b�E���.��=�T�R���γ�vD�X ���ɻ��U:T9�ft���h����X��*)�ν��߈�7���}�W�1�>~]{
B�^!,.B��_�*��j�#Ⱥ��ft�2*�����98�M��+�n���uM1J���5�����h��B}�ԍ%5���E�����m-����d/��&�4���*|!�����}�xv���d�R䅮|d��=�
wj�:Č�uQ/�V��1�L�p�� b0o�����G�ݝ������S�q�����YOj����Z��O~�f��|�s����&���;R�^�\*���q.5sZ�~՞''�B���j�6 �quvV�?(0P�s�3�^����]������+>[�j}BZ�3aT���u4-�޷���}�=�X��@>�y�+b_�W�=�[W��L�l����� �r���t=nW�ǐ��_
���͋�F\�aS��u�����̹-���;�G�8K�5e]�N'��
�[��fe�ZJ�6�{ � ���HW���~�}S�G�a��]�v��@͑�����}5�d���,\�/`��A��g��Zn�4yz2�q���Z���T��_�s�ш� ��8���Vb���䕡t��p�̹0�T��f��XU��O羘����<>�:{j"=7��r��ۢU����&A�N��_�Ľ�m����#ǃSlO��=��6�-�/��������g<hl/����ݱ��4���YVh�b)g)�������6�����20qd:�.��Z�J�*qU��o�,Zw�Se;�&�Xn�d*�zL5Uֽ8%+-�q����}��I�κ£4
q�J�8��6��3���f�5-}�{�}ݜ�f_��� :�ϜÐ��"M̍� �<����4�(��?�7��<�o���N�O�(Ȥ^��;2�	+:��c��i�[�=g���*$4g� Rq�M��n;���gu���u�1tK���1H��,+��#�b������nzp�n��Wi��q@	�g����V�������.��/�Xh����[{�H��g����r̭����$0�_���������ub�C)�G�ݟ�^�I���y�\�Ǝ�Pc(<N�Τ�����=Q��`�(���@9�^���}>�K!_�^�PQ��m���k"����ꯃ�*��D��c���\��}�zQ���Sc+�@ �X
�_�1��qk��6���u�oyU��k�tN���~�)��Ѵ��/l��Jʛ�L�D38�,��Zq�r�lE�i���ʱ���\����v�S �,ED����>��sz��°���������>�@�� @��k6�}��2��o!�\�yO��3�Fr6��݇��~ͧi9����_�5�Ɠk=���}���L$��i�Xa�|ݟ:�:��Y�����wֈS��K�1�KBᘓ��.��,��D�D�J��}l�g��'q:�B�Q�	[��� �����y��x:�o��K�5^ۭ�N�h�}1��΍���TQ�歙W\?��s�H���Կ��_p�q[�r#Q܍F���$�u�a�������;�N�f3r�"Ԣ�3����dn��aY�d�3�df��¾�s���Q�e�$��	<��x\�������P�n�N;v6Rfsn<�׾w$/�/]~ xb?	����������8�m�$��������b�N��"uY�vy�3;���� ��Z���G��$�OԦ�AM���(��8�y��e0��槷[dp��w������t������F= ���K�׿��H�o�)k�#o��I��z�}���������O���ei���!���*���ǁ�
� 	�"+�S�)[�Du�=��g6֨U�w[ �S BկR��i�
�����gC4�d���O�p��4�����H�x@�u�o�Q�����p��!��R�t]�L�c�dňG�QP �hL�� �فj��K�z�X�/��|m��3&қ ��qs]櫷o�#<���l����辢{�j18F���	����u��R��M�6Л� ��)K5���˽�q�U<'�ug�;�@K"�\��Q"D�8�~o�kzHH����7S�r���^ �&"�#�c'�H�Ks`�
g��ч�.7ن�.��c����4fP�c�"��GY���b�gU�����ݶ�aI��Ĩ�~ˠp���G�g�1�(�²<Phf�ǹ:>�X�u����H�^�t&���(Y5o� �����}�Sޛ+���7����`iZ�4r�*��}���Ɩ���@!���٧RdhB�BU|��i�#4�m?�ιѤ�4�5fue9��fnK��
�!1������܊��K�>6����X:�ހ�є��vF��q���N��;���(�3r�f>�e��#Efݣ�t
1G�8�6c�%{T(��Jv`i��7�,��39{<흯#}�(��Am�1@�Mz�%]��G3]\*3~����./!��B�>z�֐�% Wg���h����1)�w0N
�Q���n�>����~cE��@�K�|����S ��/�R5�A'T���J.̤������Y'f@��f2eBUy]ӤL��nE�b,�ދR�A<kt�:�WǨ���9���� lU9~���.�Lu�S����	j|G����}��[`죌ټ�QJ�߶N������OZ�1�r��i� ��4�Lplc��Ԍ���6q�'J�ò�	Ks�پj�+˪���=9~k�?�l���J\Oݧ�-���r��f�,�HW8hV�:�R?�����@�� �	�
��T��Q���ؙ0ft�]�~P�F�:Έ�l����  j�B&Ƭn��r��۵|��D���<�6e�4�H�k~�F������H���A��Cv�bx��k=��12���������;�7�p��<�*�Rr�\��ΩNX,�E"A�]�Ӊm�C�Ŵ\�x}ʭ�x�Ֆ/	}-{�noYY�5�����*�l�<c�6gQE�Иy���jTt:g�8~�6^����4���Q:=2\FX���S���$=���]��d��'J�= �,
Fc�}2v_t	쵩�U�Ll��v:H����_pK.([�r�#�0꼔}��Q=�n�=߾u��4T��s5��U~v����dR����/Y�Q��#�ֲ��o;���+��*�>y����	=~��eB^�&��B+��	d��C�W��ǝ��ϒ��!�탼.�����d���S0����w̨[��� �v������ܒ�Q�B�cwȫ���ޤ�֊�#4c��(�FH���el���uG��5[���I��֒D���q�T����Y��z���@�[�G��-�ט��_������=zD �5��*�u�=��8Eǉ��p���M��Db�ۉ������I�)�Le����y�E�64�=8�yJ(��[���۷��IIɤ��C���MV-���������HU�.-�ح&�?�9'8���!�aƎ��eң�yY%��E^��ު.鱾�;;Y���+��q���ٛ0��".�x<a�,�C >��%{�M�?|e��Gɂ�aSܺ���k��<���n��� 7ng跄�G��2������>88oQ�cr�Ҡ&U�p����T�
�.��W�v\�E�T��=wR���ڴ��Zg�)���Wnc��/��<
X��Sc�g���p�[��0�y����T����ը$�K�ߖ�,��?��^ܿ,J߫*�w\6g+�}I
(��@+E�覍��Sd?����r�K
>s�6QN?���q7��Y�5��k)K����T�9?_��>Aq*���^R��˵�CL}�Rm4���@o"y�7� #.K��P��+|~1hŹc�+���&w%���u/�&�� U��8>G)W�����Y�1��_�s%P��˂*q;_{Y�f2E�K�Π��Rw�7+���~Tz����� 嘝����h%S�3s��\�����oS��ũ3h C�;}�a>�_���a,P���íBi���������+�m&B��K�o��.��[�k�8�����4C����ɚ�kL��O4n0�Isݜ0�8nƓ�C[A���A����Ez�g��~|�Z�����}�.@��������G��ƫ(��ᶖ�$x��a���L*��ӿ)(z}d��Pf�����[�y���X{��0� ���:8Q�	��Ѝ��Qc�oY����g�t�r����1U�ַ���f��<8p����� ��8�}v2�|�����]jj�Ǒ���~�O)��<��N�L@��ͮ��מ���`и�����X]��\T���;�?�b���l9� �XB\n�}	�ʇ_����ms���9���J�w�s�7�sss�UTF��U�6�w���Wmw%�ɮ�5��h�I?�c�]в��ge�N�s{��+���{�S��2למSQq,�f��¢�]kkv	#���'}:+�^5��ng}B�Z���cn�8������Y�f�]=�HJ3�Si�	}&��U�&����|�;�܏�n$R������Q���u�������j��	4!���ZKbJ,h�3�6dh��ԯ#�Q�Jk�Tws��S��
�hc�Zq�x�m���=��~���G>�n�L��G�z�y����6Ǿ�s��):���:�����7%E��p���ߙ�ߊ�¥��B	�G���9d��c��Db����;9UJ�7�����3M�y�Jr�N���h�\����-ދˣ��*3����ѝr3����{��C%`�upS���1��)J7��~xe7�X���Gu�����9�D
�ۻdڞ9$������T�H��`b���$����o��������`����>7�15�P�{y@��W�Oxt���� �S��g�����_�)7�����I�{�8��(��";;a��Y�A��ߗ{��q<eJ�/o8=iu7��T���������v������c�7�οMe�qsu[R9MG2d�yB! ��M5�#������v_ �- ����1'��=L��y���[@2���ꍪ��OW(��n�X�8�F��?Jc�of�/2F*cʜ#�+�T���K��M�\��>�|��;����CFK�s�����r��2Պ���~�>'p�E����!Y���ڑJ�W�a��ap*uI��?GС���0��:�8ݲ����љ�c]�8�s@�?��b����P?b rz+���x���B��T�i�~
V�+��m`�x��~�KX�|��DY)�^K�'�tQ�/Ũ��h�����;���T�t(n�A�����c��|��ԫ�x��'���n��+�b�8nM��)����G�<�ỵN������td|9�ΝQ�Lх�29zC���궎�Og��>�>���q<�7���g8��O5	�qY���}������{�)�k<����"s� ������{#�Y�-�`\6���u1=���J����9 E�F�&�d2�_����k�ky	�����b���pt�8��pc�����У��A4�����1U��O�"a��l�����"��Ν��Q ��U{�	q�9�b)�;�����O@��=�.$I�c��,�	�!���0�~%2�J�j�>%��GL�_.֋��G�)�+�hia���s��+$5�ɵ;Z��(���񪮮��ꞈ팃�M�mN��*q��a�K[����8���&B���m�G<l]�33y���z�)ᘚ�$@
���[�ǟ>}z�
#�jp��B�eX���9k�Df��;����"��z��Z1�Y�gf� ���	R����*?�����+����]��P|8� �0)�`[��/vz$�jK�띍�S��궷�$��T�A���J�w2R*�ܭ�-�8�T&P"�
��v:3�4v���契k�w%���*Rv$���b>����U;e|�6������MDmѺf��S痼]W���?����|���;��Q��F����&���b.�}Hr��e+���(+���H-6�y�������jt)�a�1�I�x��Nr����y��r�2�
�l�혉B4j	ӧ�A_9�%}M�8"����b��S�#T���� ,���0B7S��R�K�x���ԥS�m8���/�2�E~���������B5h��oa����\a����`'������:�^{x���@�����f�����L���$�*-�V��'��q^:�y��ϵȠ�E�Κ�!�����6bQ�-%�Z15��aY�ʝ�E�������G��H^�ɫu���u�x����K77 ��U����'�%ee�D�H��ӌc�i��X(e�?$m:z��~�6�g���]�cH"�W"kM6;:N<m�<1�	9�\E!˲���w攵�l��>��|L�&����������sǯqc�3�U���@yU�M���R��t 7�Sn�+Ԥ�J�A_�� �v���`�p��G�	�潽��)��w��IdGk ޿�tgBo��B�$�I}Rl�
��K��$=4�2h���)�u�����][ ���w�\?%eK^#�=�f����댔*�}���\(�v�w��Zdl����O���U�/8�խ6����=�2�&�l]X�����W)%����4K� �Hw*Kw�
+]���*,��tJ���H7�,^���}����3'���߈�zxn	������RC��%c��c��p1�å�Pfط�2�Z��nlB���kT7M&�XY�GFN�J��_a�����k����Ԟ^�r�R6U�{<�&lL6Q����$EqI�#G�Fjv&4�5" �R�ֺ� ��!.���J�\X�������fN\���:R�(��C��L2��r#�tc���,466��~�}o�4޸�ox��sXo���P�3`$� O��<���]y���&�A�!H����[_A������8���x�Z�� #K]',���e'����o�kZC��ZJ�٘�w8����f��®��f�fYM�S���K���7����yծvF�C2J3����E%>��Wc+Y��h��>�Va��耡&���7�����b�R�1ӱ+ �R�>s�pP&���Pr�DX�h�<q�y0x��LNrW��v_CV	�_M�^*)(��bk{&����V|$����:�{K����:��屄��7�uҔ8^Cϭ碓�	�b��[)`|!A���g}�����^�F�����^��w�v�H�sK�+��z��ǭ��@;�D��|YWW���Ij���T�����	�[���sc����V�����;�׾ڵ����=��Έ�x.=��3P��O���WG<����?ZY��E�S�!��؏�O�!]O^nQ�:��D��^Y]]=L��T���_�܆���L�0���F��٢���(�L
m���K��>5�j�b�i��(UV�$m�k�����Z8Ԕ5�#+��l�.Nqv���DU�bSn���a�%�����`:v�����5;	�����(�6����'�}�nY��;��컩N����~I�~�T��4i-������ȉ
��W������	�S������>�4~>��:�g��:��˵i�29�"έ�R\4�#��dش�D����)��S��V��fO9�L����}�3r7�2w��Ja����yY�`z�\l�����m��4	AS���Ttj:+=|�M�R̡2���k���ķ׶�X���LoG�Ȉ^`��T	���Z�o������]�ñ���ӞG]����W  ����_Ѥ��W��^�J?����*���7NS�[%�]�\��D��;5;V#
bꪜ�~�(�S���R��~%�(�t��V��[�L����co@[k�J[��Qcf��3�s��R���=^��ՐW/^��/ԇ�įL�:���9[��X��-z�T`��Q��4�F�B��/
u�
�D̳@?C˜� �ٻ�D�$�E�r��(��R'�r^����sE ڪ��G*Q��۷�#
a�2�)��Z�����(^`��鿴�
���Tttt�s	e��å��W��i�IFbA��m��������N��獆�=�fg�:y��T�����hh����s�]翥���=ޮ����7���.����}d����y����r���z˗���K>	�~ީN{ppP`�:g�z�@�oB_9[j5x%U��	��J'˟�X?_���e�:2VN�}����ff����^��W������#�W �1G�����r�:a��b��#p˽Mlp��o�;�}�r=�#(H	B$i������
�ߺ�;�������e`
�?��L2Ͼ�!�/�:t������V�4NNN��&���R�A��\��$�PL�x��Tc�����`�>O��7_N�GU�*(�323�����\����_����_��5�oJ]CCԹ��]##�`�����W���S�f�o���)o�h��-��H]"�+��KH�?�u޵�������O�����]cc����]==��^����NLL�/�W��X��t��EhtDDD���u[�薌����2����+qqq�[[Ҁ�⿅0Qd*{l.����GI����}�
hxf5Rnׂ��u���f�ꎾ���֦��`]}}��/�r	(IeeB�Ô�l����􎯒����ߔ�x +ۚR����{���߂
o�����7˱B6A}}}fffQ!{�Ći�X��Z�چ?&�
$�q��&;��Y�ntt���b�W�`2�6775*������%����gZ4���F+vww�ݑo�� �vS�xp���qR�S�����-3��3������&��g�A �B����M��/t���|]�i5�qN�}8������H�� lH�Gh�ߛ7�������#X�9:�oni����(�Q8�6�=�㷌�o �P�o��Fi~�h��_�ffi�.9bт�z���m�V���Xn��� 8oB_�Gh����Է�����jr�r/��74J����-����cNɩE�G�n��ۛ��$\^�[C�O�Tݗ ���p�wy�4L�1��S�t���IX�^���.����{�/[�6ek$������rh��$m��?.��Hȸ�fB<c�"j=: )��AIii�S?:J��կcZ�x�	e&#���áW-�C�����〹�ir5�<�$$�ہ������
3��k�!�o�8�̓BϝU���C��-��<k � Ov��vyɃ��X��H�4P,�}�?�����7xs���������ۧc�������������i���x���%bb�u��%E�H��J'E�[��h^룗�:chsʯ�T*Ǌ̗���b��D�z��R�XT&D��@8`�L����-###��Q� �%z����}�����	��;uA �Kz��g%�*Qdgw&����!@��1����OEE|@a���9�؞O�q �,�۔z(�\�/�*��l.�I�U�m�ID/yt;�*��}٘*���ݧ��D7��od��y���N��G���������ʆ����o�F��w�H�j8dbBmLf7<�v�8��j�t�[B�5ZZu�H˽9������P�I�?�.�y� ��0*̀'chH};��p�HrW�f��`����v��V&��az�w[_u���<l�������ͧ6����\\�J%}�C1�����?��l��*�un-:���1
?�x���

�4C�hK��x�.��<,�uI#�k��b�A������.=�zooo������GW� ���l����U:e?+���;�+�Y������ �L�%��n}'1�����oݒ���ѿ�h��S�$�PE�R�֎E�Π�x+6dzkOUI���C*}���㑮�UXXXn+6h"�RaZ�	)W��9���4=ʮظ�2����B��CqBO�(���x��{���->����"���%%��F������ �+
]�	��Y\��x��h�_���n�=�� ��d��*-��o��H@�W�$��͸�쌌&����z������]r?9T���{�T%L�l�CP�0��\��kk9;�g�?�)��}�S�Y�!ƚi�W'f���x3N��6�J�ffgˊ���-�6�8˰�'�x��4��x�}LM�.�~^��CD�TVV�H�7���^߻{���K7~��L��xv���R�Vjʮ���5�I~ܧ@��a]ʿN<�ƞ���N�M6�U^��j�E��z����x1-�mKK*���[��G��	�'5�G_[JW=co�g�קv���6<k�m<<��=<t��$�\�ӹ~7���CU�x���D�8���1P�D����͇���><s�Lޒ|Ł�&}��#���n�e�S���@���R�VS�Q�L9l�P���b����~�k������F�C�v�I]���������z�[�Te��˩����� �9ؠ���z���d��0X.SfQ��Ж3�4@��LW�(0��p�4@�n�Ȍ�	���w�g�d�Cz���!��.R6MM<թ����OQ1X�m9�K�D?�Gn�����dQ�搛�;ۋ�<�뛛�����e�X���� ������vv��\e���@TLll�#&�3u_����H-�?����~���x(s��H�u�J_�OC��|��������d�*h\,lJ8/��w��g�a�w���V��nu'q5�g��d�����b����� 7������֞�(a]6���]]�7�3&/󱜾�F⧹d���-����b�歆� ��Z�>>1���0&�$���
|zck�ʝD���W�V��.ՙ��3AH��OE�-))	I��x�ߑ��.�V����Yck>�600��^�u8����5y)�?��	�����"���]A�������������𤨇��z�]>�c�27WNc��=wj���Q��>NU�ߖ��m���L�C�����8w��͎���lK��䓳<j1�Y�㣦�r�AMC���X���amY�eTTD� ���g���1bf�.���8	�������y	�O��z��d:Q�R�5�Г��E~z��7h��M6�@@� �V ����|��n�ؗ���sf>=���Y�^C&�C�%��W��*7d؉��K�ى^������S�[R�XpD+��?�K����<M��9����@�Y�)�L����������Mv��F�G`�c���:�z'c�s�tR�i��ữc���w�"T�Y��Y+5�vq|$�uư��}䜋�@W����{�������:��#����BBB�yyO�g����9���g ��2�I�S:�P��ǹ�睊�c���Ǟ�ǯ!^��_���V�Xՠ�Tˬ-~�!�yyT�U.��¿X1��H]S�j�r�y�W=��B4(yyٚ���r�ڍ��-���ytؓ�P� vl��4��c?�
|�D+?����(�d�LI�Ǜ�E�/V?�R��!��=�����}��h�8>��tP%|�x;��7�"��7AЅ���/�T���.�8I: ��E��$OB,��ؙ�lZi���1��k����F��Wx5,HHcz����jd���f	�����Up�0�w�n� 8���dE��2

���쇚��BDEá́�O3�u�.��ﮜ������F��tp�p�X����f&��|4�%�ij
��0fw�x4�]h��8���/A!d���~� �DMQ�r�Y����`����i+%v����u��d�q	љ���s�f��-:���:�[�?̥�@jME����"�b�е���w�#.{r����?��J>>�.I���P�q~��������yw�?����5!&;���^5\z��X
t��G�J �?\u899�99U�o���߷taqQ�����.���I�1�����;�p+�T�M��օkྼ׌�������d__�5:��� ����@)�@)U-�,��@����Ja��YUUî�I'q
���F�Y��߸;+uP�G�)����M1��/N��˷�.4��Ns�w���@�'�=e���=��٣�{��V�<C�k�c;��؎j(K�04a7![@�R ��Y�	�J-�'��S���A��_����ZX^Vc�Mg��c{���*9��aq��j�@,m�M+�����1q����hp��n�^�� Hmm����rsU��31���0�ZXl�j���E����ϯ-���d�b��ъ���[�ŝ�,N!������R��C6�.  O
ZZkFC(�5x�Ull ��b��^�g I���C�b<�v��ٔ!�2ꦎ��"i !���I�� �4 �Aa�?Tb�;:�k%h	�b��Jl�3V�?�v�3>���e�q����.شւ$�m����D����!# ���1g+��7Sɢ� �d>��Θ��ɫ�3I$��c�T5�RE�u���	5���x ��[M��uT�m2�� ���R�x��V�(e��ڌ�<TUWϮ��JThr�hS4����xg����|���I�~�r��P�MB�����Z���+�v�R���� ʚo�Y�^qԲAU�iƚ�}���q#�C6c�XQ�舾'l5����� ���t��̥O���n��@t:�	����OJ�̴4)�����W���j���k�dl�����-��s�v��EH#%��
��Е�)a-�`���X6�i�-�u��z���kHb$�PH�hm��5kcl�����Z7zp��<R~8:�����H���)�^$��`����:����*qZT���q�23�1QO+�s���9��I0}<�X�[�x5��*swn��mw��j�W藉9 7`��^������%�^�n��G�~�9/�h��|"��<�*���N�%Tf�A��.�ӷ�N���G�EC?^h6)Z���B�~������x�N.��եH|钙��0KZ	�ĵ�N\��#倇�O4�jw���z�0wuIۢ��m������	wK3��d��� ��r�s��j�U�&'i��VB��=}����y����q��=������a�v��ʘ�(>|���lUs��| �����ѭ��B^UUՓ�n�R<ğŧ�)���a�f@�ݜϢ 7�>{�yT��f�w"��}6�g?�r��A��+~��C���L���~�:�
+���;7w��J>�UyR8�YA� ��Ԡ�ߌl� =\zm�S��r�N������~Ȥ��6}I^z4�֡���U�*��h�!d�r3q|>�t�K~/�Cl���1c(�塿������@�[~^�ey?WFwUdDD@n ��N�MM8V�O���++�zaCG�^^5��H��?�(�}�Ձd�v��+l�Gf���:���u�i1^��g ��6�Nɤ��Z��B�D�خ��5Ͻ��ƫٴ���FYY�B��Ѣ� q���b�ٽ�Q]�s��M��ސQ���B����g��(l��2��:N.C�^=N�c/P��Y��Q�BN�{U�q�PìA,���q�2}�@��HT
B_KT=�D~��?�����;p�i؄p4�=��D�� A�Id�{�����z����A��J�J�c�5Em�V��H����פ���Y�B���Th!=w���ڽ��CV��,zw�_Q�����J��ڠ|������KY�Ŏs_�<M�7%�\��k�`�����Δahxr�(��?�8��r�?�`���W�S]H:����t��()Q��a�G��Q[����U�\Ba��ҹ=[����w��a޾�[4.��|� (���:
= �~�;V$/ۻ�]���Jw��Lށ��jjF���(�ԅ?�vE�� �Y��G�`vYp��(.�wk�M	��;����P����mL��o7�E%���6X
�(M-qXm��?rwj�๪"L��F	�^�9��C)��+�V��ҁ������ggg�J����E�~!~c���.QkO�\���}ZՈ��Z��\hh�V�2�}��~�P��M�W]�pK@�ٚؖmXb����@)�ԹN�ӧ@;�����}v�7��b"�����iI�#��Q;Z�e)<�8�Q۟zn\��/:���gk���6y�l�֋�$9��TB�-�U���.cOY�m	�O��j�IUE����^�.�_g��:;��3�k��7�j�Xk�I����P�#����Є�3-	�W�?�G��s����e�U�_�!z�\�RT��;��GS/	;}p���4�N��q1�YUg�r�����������wc;�fz��\��*������m5��q�l��������	���9� �K/�	=[-�m�RҾ�Ψ��B��U��W}��E$zGΝ�\,gV�Y�y����&��t��&����� �V'�	ș����v=����b�ϋ0T���Q�;�Ui}+��YݵCqRg�K
��&	�Y�^�9�]�s�Ǆv����H&��`�"w�kV)f�� ԅ5�j����,W��WP��Wt	���N=����˷�m���b�g�+��f�|�t���r��(��aƸ�O��v��ѝj�;81|�
gB}������ùSV#�-vL�AW�ծ���f�,Uj��`�%����7�A�r��JE6�N�P�LEk�𪟡f�T��L��,A�d��5¥p���z��^�2DnիM!�2O�%J�=8˙͛��H+㎗����[�1
���;��5����R><1��}G0����(�/	�+AT���>=�����s�B�����lf���fw/n:�\#9���-m���PZ�9���¹��%e�qf=�J w����C_v�S�;��k��
�i2�Y&K9wfګ��o�Չ?��E8�n��?θ����ֿ<�M�ƙ'��A
s�Ke����9�գ�ͰF>�<W0a���n�����5ˍD����!�=�7��}4x��Â�]77^�.��ݚ,5-��z�Ie��}:"���)�,S�A��biQ�T���oD��˹�b܋gp\i�6��}���&�U���X%�٫����L���B|]��fK��R���Ɖo)�1jѲw��<��\�s��w����o���v+f�1J�e��!3���[���b�A#gv��D	��(�� g�2�$/~�r,��U����e�sAS���QA��STXԧ�\_���I�^�bկD��K�F���K�W�?�
b����k�y3���j�z�~\�A���>1��ה���vl��ӭP�U`�B�2s�8��GLӶd�<7���S������L<�.�P�9`4��P��wd"(" ���!��2�Bh��~�����i�ͩ��Su�Aa�2�7FB:�| I���̰������"�l"Wl����]��9�:���rڄ�r�Y��J�ƙ!!��g��z~/D}}'70oC�)*e�;*eK���|x����O`���w����s:.f�K��+�ul�p�i�c��zu�6�}��O�td#h����+|ٗ~X%��d+9��mG�����T��B�J�� H��]��/�b�X�]���`�v�=�,���t	ۈ�LM��rC�i�}oʟU��d+�hs<{�Ԙ���R�mP��aZ�v�\�����j�z�Lq�!�	@���T£�fn!۸1��G���zr� }��_���s�rV�>5%!��ک����w�{{f��W��H(s�w��$����E��p��'��d"8rY��S{�����\G)��{�PKE;%�1���.*�<��!�����/)<�A>��!�ckd-�+�슱������m���*--?�N7P`ZXY�ӝ!+.5L~C&V�;%��:*�Uqf�a� W	V�fiQ�@��jB��U���H:2�����Γ5��1�V;W��*����	�;��p+��/_�����;G�#&�·���#z2�o�{���&��ϡ9T��¢ڣdE��*�v���KUّa�#Di�KRj7h),�5b���N��j�o��e3Rj�<ZM�\��勫��#��Yw9麳�.]��0��~��:�����!b�z�"l��"0g��Kɔ5�9̻��,w0dw�c���3V��߿�L�^�b�0Z8�	=�yJWW7�������N�Q���så�s=�gL~g�Ɍξ��t�����D}����kS�w76@�*en�%`�	x�3��GX�:i�AӾw��Ҝ��4��f����ہAA1 o�Qv=��0���{����l�=�F��55�����!q�g_10��-MwS����"?*��B(�i_�g��?�RS���yS�u��Nh+�۵��S}cX]ɠ6�i�#�(sr�P��tHt�/o�3Vā�4i��U�Wk��r�W`����T����g��z\�&��� C��UQLG�Uo
8�TK4�I��aٸ��b�����C�|�2ā�C�{s�@N�=��P�;�k5z/Nu4�-�?Si���W�C�f�r�"ʝH�z%�?[F��;ܖ9�d�U����  �}�|U�ec4�;}s��NҜRj3n9����x�A�I^�v�kI߫gyb|�BG�yI��if�ߍ�)ֿ
�E��teRl�����s���f��
�ْJ�S1*]:��{.Tk�O��E�ͱ�]��Ra��M�X��v0����zd#�-�������R����밴�_6�P�^�����InN���6�����k_��N%~�d�2�HN�MʦH��MW��M��.c�\�(	�2�;��9�-?�4��7?��a=�(*R�#����\��aܓ� �o��9����m�[☠_��=<���D��)��z8��p��~���Cyi]Na��$��MLM��⭤W���}C�mq�����MrC߆�\Ŭ!O��k���	��#�Сr;Fy(�W;ڒ�Ld�(�PP��{�e�	)��Iȉ�~ۏ���@E���[��TfH�������2:NOXƄs�}�8s�w���l�H�C}��9,u�����yi�)伂-�(�	��z|� ���*���e�t0����d�����5���4p>_;����c�U~�P�)N�떋[��q��*�m�v0������ϋ	���p/���2kk5~j�t���ͬ�"��O �JJT�+Ia/>����MI�WN����˵@Ft~i��q�Q'o�OM����8�u���p�SւA���ͱ���?.(��;�3���l�����U��Q��t.������<�+�ic�ذ��VVPNNN����n"����7��|mn�����[��Ťʝ �ாL SM.�oƩi"�����P�)��x�8����gપ)m��;�H�*9���ҍ�v��3�����0�%Ҩ�<=��W��Н�;z�t��c�r�D ���v����+��-���[}�
�P��Pf_4����|	���ܷ"]!�ޕ��@��\����%��<s�,�܎�fFb�J��2�cu|�� u�\�vY��9~� ��򟾜�Q�[U
��V��Y���c�,�q[��ݜ�vl��I�1�:��y�Ң�U՗S��z�b��W�|K��v �>!�)h9�l:Bb����Z�U���|,�p?�'�_��Mp`#)d̸��Gz�4XUR +�wC]`2%�������"A��+�eJ�x�;9:��?��Va�r���,��B^*�����"�;?*,ꉱ�v$�ѭ�7�M�h�D��bh��L�޵s�zSh�2y�~�ah�CK:K�n#)�~3nͭxǋ��>?o�;��(g��u9gx���-���	y��j��$�iiR�{i��FJgΜ���B����Უ��ot��>|������Y�I��#��GLL<�1`���dIKro������Zsq�����1&��͟���IM�AV�ep9���oN=�F&8�V��K�̖��v5�v��yl�Q���%xOgk)��3-��,�Xٱ]6�gZ,���Ιm�]�W+���.�)���?��UURJJJ���b釫Nrr25H$Q�G��S�Դ�=߿:�ܷ��EEK+��g9��nL���� ���b	1�[;�D���aUar�7�����-ReIW��-I����Y[�|�p�s�sA�E���R�-�Ĭ�F�8I|�S�G������x�>N�pd=�|�&!�$f��M�]���V9�r��k��!c�[�Nk�l����Wr����S�uvz�}�+�*��w�Pl{�-6U��f���+�	�T�Skk%666dB����'��W0]1�����RH6V��P�5q\I��z���|�F�\�����_��I��>R�X�"��Dr,�`�/B�����Zq&���F��`�˵+��i���ؐ���I���/���NS��-?�GgCϣ�7�K�e�������8�z%�9O.�,�а��C��@��4W��5Q}�7�rk� #�@;�y��_�A��+!oYx�j������gg/�7�s��ue�	LF?���vL�誫ke�!W���F�K*l�d1�_<\|ҭE���y����A�{�����H^��@��'li�S�{�t� M�F�{���+�/T&6 ���:V@0�/1���IݬdO��k���� �'�'�/�^-%�q�s?�����J�=�����xWT���g]����YV�������a��6�����A�b������#M�Z_	�c4�!X�.�U�)�M���)�%#=g��y�ˠ?Z8qȪ�o�l���0|즗��.��J=k��{�7����~n�Qr�5)sɹ��g�U~����0�VlN8��m�X�Vb~m1���謸��0���r��~N_��tj��&а5?��{�)���*����%^�&y���	�ڤ�z�WJV��%�s�����o\X�ٻ(�
$:��Nhfrˊ���vB��w��I�VU�zx햍��nH�5��+C�շU��Uc�����Z�]��$��<\&\"Y�h���Q���9�2�󬮎9R�aRI�=x
��c�]�-"_�q1G���ʻԮ�O=��)��#�	R�)�*�-mU�1c����07k�T���⥒$�o�M$��պ�)?3b>�?U�c)���W+{T��L L�?��}�Arşrr����,�����6S�{kHG�u�����<���7QT��	�r��(t�x@c�.��6mQb�������Cc{'[mB�A�pHs�J�G����ZӝpF̹��U"b8��b�I�x��s�T]��0�|u�<n.z~�+ɂ�H�
[��c�����t�
-^ڷ��I=���RW��/	��3��h�n_u}ǁ@}a��a��1_S�{�%V	�>�^KꤿV�x7$�KM��]#���#S˄j�üeHs�s�˪�� �&+�B��N��d�;��)�Ls�Z�ݺ������g}�����&ӻ�ɠ�d[�Ļ8hO^�h�]	Z����!�Q�4�� ,7��s��h��P]kԷ�10����I��y`j#��9�r`�,��t�7��u��Pތ�ҺV�����#�@-b&!~���йoY>���t�U��vp����\��G�jv)�Z[a��z��DI��=����hT٧!V�k5}������o���>�3]�[d�R���qǢ����H��!�c�քKb��t]K�V�:��`������X�U�1���T� ������"�+�=#��ڌl��䳧<a��Y�^����A�-����ړ�E�a�}�Ӛ�����%u����ݚ���Wo�#wEyN�[�a��7��]�l!%�<���b��TZb�#���o�.y�E�+�.~��D�Sd�d��O'vY1W���_mIa���	��T%8�U+#��'.#�F��2D�U_A >�4�9	������rh�\����2vZ{o�4�I�U��G0�p ���RHʄ+4�VFi�A��ha͵�s;idFZ��1��Z�e�v�q���1?}��x+�!����}����~JUo� ;'B��~H�?XH��x��pJ�=D�!䍢�h�h0Ԛ��ƶɹx��!+�ƚ�%wtS%p�u��ϿU+!�J|��튍���������������tMa���KZ���}40�=j�����%9h*�x[:c��A��d/G1=/�RZu��YBݞ�,`P��s����� .���98�^=KP��H7�C�_T�

	����Y9��7��Q��<ߗ>>H�ֻ}�ұ�ʹ����A=���2A���>��e�:�xt��Ѕ�8M���D���b-�����ț#�M�&&ٗw�ᔼ��5��,��H���}�I������s[�f�e��Q�|�*��;�6�;6���	Y�ܒn�D��;�
+�
��х��.V�}v���0w�>�Z���RN����p��2o}��+��ǯ���$Ӓǧ8x�e�-42^�-��N�9�V)�����s>^5ǆvk"�yz�k�]xoq1q�1���O�n�>��g�J������Du���$$WD�E�5&7<��5�����Q�����V�.�s�й��h���h���~�T�흣�j�ru�e��;�������ZD� �a��Gs��NG�鿖?l{;�$Q����#Ӓ:T;덾��Q��-��LQ�����c����	+���LI�a9V؂��+�;���>�C�vc�Z����~4d�8)N������������=��)�d�8���0jC�M�?^��+�ן��f�U���.��"%�I��QoYi���go�
:7H��뾻
I�����Zl�� �oJx׺����K��X��rg�UU_�Ғ�>���@(�?B�2��k:��B$?G�\�6�+���ь�>�N�P�c��ƃ�;Gpޠ#�ʵ��B��T-��>Ii%�����^�"I���=]u\�Ú�ƞK��,^cq������6�v%3H�2�i݇nZ��!��DK���]j���^A��ъ&����(���CV�����e��U���E*˻<V��[��}����]n[:%-����>n��E����$�&!���8�x>>1~���:���ײ�צּ|v�m�;�F�s�G!Y�A��o�m�gnX�h		n~�XJ�@:���n#���,�����~��ò�W��:~ó�ٔ�~'������g���Q��>9�/GӦN���ZWn&|��F�\��|�Ԃ�sT�T�2����KI����������K���B��
K���:�wf������;]�d�8Uai��(ϸ2+�w�nϻ��/�fCM�e���W[f�8w�fZ4�l1K#&t�S�v����2�^�59�
�0����ܱ�Te%1A'�T��e��8�M)���p�f��i訚ʪ��3f��n&��͘oy�!G�����g����T󦝇�myD"���"7��:ڻ��q¸�A[�0��dd��
���P��e;�Z�*��T�pC�f̓y}���A�M,`�D*��s��!=�%�A�<��c�O��1�Ru(�5�����'���*J�й�MB�>��3Δ�B�f�%|,i�PR_Q��9��sY�NǵG鎋�_����he��B���H���>̤zw�����+V��(��i�Ӻ��2�Ў�۽�zp�GV^�T����)��!��іS�,x�1E�j@ߚ�	�I���ß<�.X�����u�RvYx�ɤc<��۸D��QY��N㼆3���ÕlY��
�t�{p\܉���#K0��kL��
�n���17Ar�ҹ�Z.���'/77#M�����aʴ=ެɦ���_p�+���m���k�c��t˭�����=�������F���8� �t@�O1��te�
�#83|B��څJǄu$�����
j�eX��U)�s�1m�4����ؚ]�E��|p����:�U�,��X�氞j�U�K'������+ʎ���?�6�0'���	�=��1��Zm�x����8Q0��,@��AEo�癲u��@>���w�N�������7x��U�1�K�Έ��x�c��w�>g1e���r[���cȎ1�4r�t�u��$P.���Z�%����e�>!�s%������G�-���珛ch�}Q���m�
�i+�b��XX�B���a�i��l�oz;��,�_S��"�9���F�,jk�'�]0��f���n������ۨ'�+_�b6�̚����򼯠cYv�G�޼U��2�x[H�!�Axb�U͈<+�4"ĸc�n��k��0z����+�,��F�r$��	z_R��x�_�v;-a�i�3�I|MN(nn�Ĵ^7D�E��õSU!o��G��&>Ω�MN5�N��jkЛ�B�ý[���ˉ��iEK�Θ��O�r��T���嬅9V����y���HQ�C!D�o��^��W�?d�IM|����
��
�| Ʉ
f�=��$�_xG���Xƿ��$�&V�R�_L�b;�܉	�8�����	F�Ɛpb�B"��!Y�y�X��&O��}� ����8�G��u���Y�sn�Ee���	ۅ���tzmr�Q��(i�%}m�EoV��b ��yE�s ���so�������|��:����!]�4�l��'�KA	�:�n�3޹��R���h"�>��آ���u��k��,�zn�1 Ly�WF=��]#X��!�>Y 5��̓d��ˀƯLI*�T�Y/����T��a�\�q���6��hcI�x���=�X������Ԣ7� ��`���j��Obe�h)C����yQ�����������r�?�!7#*�U��_��v~�GA1�jm:��(�ꐾ�ߋ R[�Rk���pSLQy���Y�����uƋ�ܓѬ�Hp��d�8�bp�r������N��-�c�2H�g��(�]+|���&���d�H'T}T�U�۫w�����;A��_ԡw+�VUʺ�I��_�a��t�,�g�vDӪ��9ͧRF ���([��"�s-�k����;w�P:e�@L�x�B/'����o��3hn�,�IG�Kv;���H]ĶP"��ˬ�	ե�O{S&�	��3��ä]�:��	�����+ɭ������7Nl�����f������.�������2��z�1D�����ѻ��/D8�t��>�~ٞ-ɠY����B8�]�`�LxP9v0�9G�[���:��~JowO��'ٴ]jk7΁,ș��q(�~Ё��z�O��q��%�ڃ=�x�'N҉��%��$y'�k�T!(���_�V��g�)�r�.D@�GMգHk7�Y\�+w�)8��Q�/RUq!�<�i�N��Vu1�BLD�����_-$��F<ΝP�.ྑ�t�ցT}Tqޢ��L]����K�a��7��q�>!�6;*eF���7nF��=h�_z�U%���u�}�d�n``�Ҩ�<5���jB�u�j���|�E����"/MȮ�bd�(�"k�����|l�Rb{Q�����%K��p��[�G�H��n27[�����I!7�Zo��G�L�LI��B\$��l������������T�!�$���E���FXFG�#m�x8T�o[C�I�@c�\x?:y�C��Xf�M2����YN�cO��^N��3.�a=C�C�K������!���Tm��j��ô9���\��ڒi��匔>�s:���ºw��R`d��4//WL�^ʴf�_�Cz��]hD*� ���ԕ��<%��4ܿ	7���W�6���������K��}S�y�^���܋��<=�N����*o�(N��U�Ҍ�K?��x�s�|{l"4K4��u��W�א%j�p����v�`R�J�R�>=@#�j�^0cɡෙ\ωs�ߔ�
��gV&LD��zS�TG�����������t����\�f��N=�����1�$�=_)H=�Wyf&�uS
�l~�hl3s�lh�砾B�iq��H��,� ��q$
Ő���/��*�,��$[���?�Ye��z���Hܜ%z�{�5ө�i"�$ktYV�Fg��O�T��Oz�M�g߹nBF��<4�{v�z�p�"���u��>�5	��8e0��1_��n2gO�AZ,���̽{�<cI9Vi�@�?�B�b�75�ߧ[v������Aqu[ yyn�IB�wx܃;��� �K��A�C#�K�	��xc�6�����n���3?曚�*���k�g/y�>{sJ���u�%+��%��$��_��-薃���e�N[�S�<��
��W�����͓"(�^p�Kʨ�_���+�S#�Dth�'eH��R������c_]7O�-T`�ޓ�|{�ApW=gØx�M�~�ș��ϧ��Qq7�W�����0�>9�8`�П�y��qǴ6�\yG��DA9^��<��.�|�}"*|Y�y:�
���N���G`�k�-ז�:�7�����qk+�*��y����v���ߍ�d���"�{AY������8�j�o��W�i�ى<%����5�хE�À@�o,|ƍZg�ҢQ(FtkU��7�}%0�����aŌ�dwz�!���8��Z
�����q'D��A�:�Ur��IX��J�V���|Ɗ�;6 �I�{r 
V�j�!/��5�n��-�QQ��E�1�J~Qg�D�q�ҏ��ܲ��N��sƃW�� ���ǈb��X�e���r�c��(��C�u�w�O2���R�����L6�O��_yݴh� g$n=v�����U-]�>��M���}����u�- %�)x��ţ�u�� ^�L �zp�]��5ʛի��JH�]�j����@��ӖR��o W$}���>�;^5�A�ԏOa��j`!�-��]7��`4�b�F��B!�NG�{��n���@^�Q��Mf�Y�?w(A�d7s��fFšÅ������G��ͭ�|���~�ޑ}@��J��8��z*�e�R��'w�Z���⋱XJ�	�����-��wG��< )#�zzjmg*�?�{L��r����!��\}-Dj�­�w*�����]>U�0/X�`I��3���&�ua�xIa�C��o�v���<�(S5��9�?�.�t��U,;^$�΁�
�V�N��R��W����F��j�Ϥ*xQ��|)��N��?�#*��[4.2ɏB�m�Zt8�o
�<����W2�q���xIj�/�U��gK�X�,r ��JM����:K��4�F��7�q���}!M� "`SE�֗1PA`pCE���>�+m��s�#*�2~��ݲ	�|���}��3^��
8���`�p�����(|�C j6�O��c�!���Xa�+	���^�mU��q�c��l�6>�������x�Z�+����y�A���'JZ��ҭ{㌇�+��5�,��Y�֥��\��I��m�]_Fr�%��7 �a!<E�x�d>s;!�31��r�<�h�;�=Z柨
~���n�X��ٺ��*���p�;_ngp|_eZ�V���az�6ؠ�)�J����۶��+C{P��o� y0�h�� ����3#�t8�� ���͈ �]BP*Ͽ�s*E��]��xU�L`4�D�r�@�ԏ���A�l����G�K��'q�n>��]o�r�Pۡ��B	7��Wv(�s��;Om�ݏ+�8˫�%�@7p�}p� 4�����m�^�����?4�*�e���ϕ0����yp%����C���g�k�^ފ�8
�WAOĤ��u��QP���� ��  H�dJ�W!�_Bc�����k�'��c���q�+i$2�M黁f'�f����.֢��	��cݼ��qw5!F3jd/�����R�	����^�������E>a`��D���a %ۛ3�ͩ��'{]��~����fSC��Xʴ��%U�;�Z�}tل9n~n{���g�?obz;]-� �I�`�ڸ���<����8s����Ź�g�܄AY��_������!R�@j�b5���gK��
{�	Eof���a!�-�_K�Q.�r���gTUq���Y�lZj��	����UyhxޫwU�T��?�XV�#g�8<�v+��̆_�!�K�W�y'o&8t�T��?��	#�TK��q�Hg	�ɺ'B��)G���?}>42N9� ��� �3��OĀ��b���@���<�9r��t����oIsŞo���11��fW�ޞ:���\��}[�A���˟JR=,Prw���ӯ��}@�0QN����2���Ty��1vO�ط����!���H����<r�:[{�քe���2���z�eʣuS˶*H��/>+'�_bKU����X�?q�M�lH�̍-'�� z<G���Z��c��`�ʳ[�N^����r3	 ���L���Pr��Bd7���|)ױH�O*q�U��z�-?�o�y0���^K&��Mw0�� qe3]�foF�*L�|�*�b�Aըz}��̞� *O����m䝜(O'�iMƩ��Hʛݥ��%���WP2�T��jb��T��`[7�\$�b����Qw��Ѓ���V��%2�f��e��3��]T�}��W�D%���f���S��MH��M�ȆZ�&�����{�s^�cP�\ɖaV�pސ�Xh`gS�����M�]��N�ne "�D��PQ���&�O��-�B���ZN<��MB�ܲ*ß�#�v�X( ��F�e�>�|7�3��0鍽[����0 ��<��S��9P�v��ă0�/��l��w�ܽ�9��+9>��z ]�N6c�L~��W�K�FZ��xZ�|���G���=��������1&{����˔�_�1��<�w5��=�N9:�u�W�r(hc�8�T3��������Im�&�-�U��?�M� �U\A��� �cË�Mgy���8� �t����͟�#����?Ӗf��C��<��`�a��9q��z*���ê�eߏʀ3�q:$*���W`�4�{n��V?��\�e��t�(׎to�����Ɏ�_���ϖ��QEA��� �w���F7ƚA�N����}�Ӌ\���R�����q���Z�>�
���\ȣ��3,m�y��ʁ�U��6�w�����e����/��j�}`�+�q�ȷ�zi�އ@m��w� br���z$������"e���?̻������R;�#��=��ɏ����˫<�u$���AY��U'pa�`��u�}�;rb���N��x(��-��QϠ"s��d�]����Sg�	7�'���q{���	��rT�2�5%սx�Σ�Ev��[29��``PtK������ٞ���b&��*�%��Z��&��!�����`��tQ�� ��l ��m�����9<qD��g�����;�G�ؕ���̻�j�Mj����C~��u �����:����(㓧�b���p�ݬ��R�ͺ�պ:��2K��}@�)����5�&a��b�+�z{��v���	�S.s3���ܜ����}��j����syA@��=��<-�=�@��y95�;�
�ïO?Y�E�����rp��Z�t1�m�6������3>1�XQ�-QQV��%u�_�9;x�l�����
%/O����>ew[�&XgP�B���"�$hS�	5��v~ԩ74�<����Y(6{#>�	'�.���VD킳X��o:Q����0��ܙ�-#
NɆ�	ȃD��H���;��zs�@�|���o�Fg��'�Eu~��(;��?[�u-%�\./��Q������r�k�϶t���<��ݲ�d�Ո�57�<����[��5i���Vb�<`Wj��tj<���d�Ԃǫp��1 ��m@�uQ��� ���IR8X���T]�C�ÙEK��t;�g��d>ա"�����-�7ݰ�<K�c+�!��Lq����y�}���D��B�����<}�<�;�K����L,߰��G�Br��JZ�]	p�"� �t�u}�kw��+l�O�R n�ų
�u�~�a����y밠q>��a�@���=p�t�
��G�C�x'w�·w�L��<�d#3���j+�۲#�DŴ�`+�#�g5�1�����}�{T}J�)��@@Z8yO2�7�`�Ra�����=�i����U� o4�Fq��Tզ�:Yvؔ:��,��X��|G>�4s��BK���Axs%B�"�h�O��L�<�=�Y��@��ݫ��:����s�	6YK����$/bp��n�;�U��p��kA-B�B���t,�.��u¹o���w��;�(	�9��Q�6xe�L.%���~k�WK,���܋�H͊
`p���R g#�Bπ�½)Z��'A��P�Q�d�k���p_q�Hp�9dc��mD
je�52���_�?��KZē
�%�j$�1�D�!�����d����w���)����jT��������
ϼa�@���~��Y
_��*�l?�8��bV��\U�$D���o*�-�@�W3ֈ�v�ߑ4&�<c]�d�z���K�Q��YQ�e����GtN�U�&�28{6)�ƕ�O���y_�yd��S?�y�!���������^�%�7����z�(���6����o]/��[t|�@K]T�����G���)\ǥJ���(�I&���bZ,�Y����RO�_6�L��ۼ6��\���zH�	�~�]j��E��[�6w�	r�a|n<�2���4���E�9GΪ ��Z?�d�aN����]��{v,P�.��%�L^{c��� ���ԽϞ��o}f����d�d={���5�mM3k�N�0�������p��~��w_;�?S�␵��z�D��̫	��ŉ�cw�n�aVzd:�4�o��ñ�[]�t9�}9�Gw#=�������Ի"��3⃱
�C��V7ȯt�L�Oi����p�9�v��b}e�\���e��+�n�ɓ�.��p]�]�Z�}��~��P:�A.Ф�ZTsz4�D��3ġ��ps�e+x�z��x7c���3vS�q7�l��Qb�%G�U�C.��X����y�^�>#�?[Z�]��_
#"���#s�����;2����?땯����C����㍽�#VO��'ⲝ��>�Gw7�n�E���%e�de*i��A�cc��v��X�ϖg߉+cH��D�A�G��p���)O�J�6��]�#���"&V�Z�zԕ�����O�������l����]��7�
�M����d�|�a��I+��K�I��x�*���nY2�آ[9�J��2Z����{��@�sl�㧉�p�N�yN�����qU�{z=ru����8���Ԩ<"�����^��w^�Y�'f�*����9��ml�5�X�Uھ	�|�T�ž�l���`���e"�X�3��ن%��	���d��a�.�Ņf�H��)�ʥ)���$��	n��ݷj^BS�d�h:��Ъ\J�e~��3�i��q��?p�s�-ꊣ�BD�Ȧ��46�����:���H[�u�h�ǖ6���Sύ�Dʥ¤�kMfE|؍a��ϔ���"��u�� |��1h\���ii!s��7X<���;�vޤf�S�d�dy����͝<�����uŨT��\'q�3��hTIUt����5�)���z4��`r\�:i�G����v�����fD��cTp �~H�����m~*h���6&�
�����>]�����ŌG#�Y_��^D�D��[>���z��M��)��������ۛ5i*�太1��N���R�d�����?<��4�hI��7{�G���j�= $����r���K�n�(3Q�
��6�$��՟z99+l�w��~y��q�wCu���ĉ4��3�_�o�J�-�$�e�r��aÛ^,����"*��B�԰�T������'�]o�EFK͜���E���c�Þ��?;B�H'u��&�X���Mb�;��2�B<:Nȭ�:Ǧ�tέ��>��is���J��ê�Ņ�����T�sm~�J\���Me4��׵+�֭��D�N���EI1��|=m]�9U�1!F<����Vr�C�(y���]�jG�o�!?�k:��Ξ�?���p�l&<S���m[���ň-��=�K(l���İ}�7��#O~~Ĕz��>6�̽����(`�i�q5�~�>bW���fM���W��S6]ɺ�� !	�.��s���
�)�X�Y�D����,��EP��X�i:�b���H����w6HV�p*��O��M�T���5#�_^K�??J�X,����>����Ys�n�����o�i#E��.Ok;TJ��A=es�G�a�x���I��!�P%���&ɰ]��o�%{�� ���C&5���P�V>���j�c
)^�H)�N��P�0U�G?�oX(Y1,4���6ʌ�S��k?��HkMs�T-����p����C/�QNb,�a��kI��8������B��9�]q����HB"b�K���$y���kkvVrbC�%�[�����6�ȑN1<�i !L��`J�"s|��,YI2�T�FK;K�k�<I�ї�q
��̄��r7�{������%�����<��mc*7c�i�l�i=P:.2����l�fě��1��Ǡk���}�6O\�L�D�O8<�Κ�U/-��zy��P�|��mNC�|�
[��,cp+{�b�����~v�������!e!��;� �-��j��޽�<LO��ӍuY���f"Ya�9��Y
ᅹ�"��:-����\	�����s�����fN�����d��܌{�����5R��}�k���=�tm�c�+����<4	�����"S>x2���/�!(���rR���Pn�����������4���X��9t���6�7�����3�Ju��LT���觊���$鋊+6�	��N5�k�+��[���EsdhK;���]nˇ�<��ڟ�y��6�ii��R���_>���	N%7��uԅWrEz�gE��&�U���-l�)o	~f�2�%��*i�#�rB�.x+�����`KO�<��F�q��ܛ�uzW1�T߿��s��͟���u�Uhm��c�X��#t��jbz��ۇ4��~����8�r/���-���/t~<9zJ�a�$��TW��w,�Uͫq�{��綺��}��V��6�OX�]�Jp��*��g��9�XD�`�������<�iU:܈�6O#l;�*N�w��+�' ǽ�㬙~T� �l*I�\�NyBX˹!&8ޣ���g��J^9���~�b��Կ%غ1� �:�V#_!��X�����<s�0Wlľ5� �
|��2h��~1瓙�xK�N�����}�F=m��_w��˷v�D��*� F�a;��& ��o�nL2D������Zc�T���{k7_�a�����h�)̼����d�R����o�sC����Q�2��r��I%=I݋E�u�H�����8��N�='�W5�s,|����Ì�	�og�y�H���%?�M80`���e��I+������1�:R{ޟhLj|�=��Zd{mz�����Y��PS��I4����l��.)��U����(5y�$ܤo'�챫�^>���X�z��X𻶕��o�o���/���O��9���n�l-�9q{^�]s\��c4�U�ly�g�t=����:5� {	a�sI���̄roZ�{��0��OjP�9���j�Gf$��ճ��y��~z�o�o}I�� ���6�-��&&��:o��eU����z�_O� �}q�L���󭟟?���?����?t�1�,lՇ��p�i����{J8K��ne�<\gx�,��d=��lv>.��l6G�R���3�u��JVI��c���r�K�(vqz��/�;��ۋ�Z�&� ܏t���Ǳ��)
�?>fa�����\s0��E{~�A������\5��[��#Y�d���Ƌ�Ze h*GZ��2�]*c@����?g$.K$�j��o�b���#�kt��[[��d"���2�	�2�߸�أ��閴ħ$+��3��-��ع�+�%-��[�X�X�薇�vˮ�Qy�ɣj��ҩ��ӣ\��Ģ�������|
�q���z�D�Wa_
C���a�2�K�Ƭ8�;K-�z�^��Yv��K��rh�� \H�A��"�oӺ��/{yv#>�v��Jf[�Ī�
��Ӏ�Usz��v�wO������>V�T����+Qu�}�c>�ݚ�f,�|V(z��� �\�=���B��ͼ'ѻP�������]~r�����B0��_��	ɤY�Z߷- @a\#��b̛�`��ug;�#�e����K6P�XZ$�=gl�9�Wy�Zu?��,;U�A�-���5���F�+/��Ǩ�����f&��L&�3�F'��7�!p>@:8.��/\���
A�'zW Z:,o�>=�>_�p;�?Tר��熱'�n�Νk���b���%R�c�m)X{��1�;W��g�`����7{8�4H93��>"&�u�p{�������H���N>��}JԶ7}|(L�L0�F&b�ѤU��M����2������W����N�y4���t�}dB�3q�g^�[�؆]��:��Δ��尻������N��1t�%�q?�a���-�60Pl��-���)����asĬ����b��m{K��x�]���(k�%���qF�NC∼���C.\��$)/�ޓ#&��~6��22
֗ �l�e2[����ȂO]s�hٔ?�,^t�`>��L�0�^N���\�~>�c���I����EX��t���g�~sl�,�m/᭽��p�!��F�G����!� (f-\Ź	��*������f�)nZ���C�Yg�`�+j��9C����;���� ��a(c�PҴG�3��ʁ3��m��e���@������t�X�Pg��%5���%����Ń�~��%��  ��@�\��/����3"~t��EBu�49����E5֬�4���v]��&��z�\�T Yr�{��g=Ք5�}�\������#/��qd��N1>��6�q7׳�p#6B$��oeU���R�71	�4�]�,���j:'H�{Crh=��P�Y�.V� ��l��|LI�%OJ����5�eq���w;��$�y+�-�r�z�zλ���:�`�q�U5ԩ)�Z�o�)W@���u�GKP�t9�z�HA��E,W�0}�WO)�}G�hk����ʫ��6�K�ݚ�3[+�ȩ�o��j�J�)eS�M;SF��p�l[{��{,B�ƪ���'_g���
�+�	@��|�:��ݧ�K��+7�S�hn}Bp=���o�.܁���> �hH�����;�ӛ�r�n�jL����[:��b�w_�;Y���+�,Z��\Z](�,�×��DBp6�쟵�w�Ѭ��8�ys�ק�g��T;���?w���q���2^AP޹_$��"�W�3�4���M���{��{G�&RlP�����F���r_|�=�`	8����wVP���������40�K�}}QGl��-�<B���'���/	@=T�S�l����	�sy��l {�f:ro��X]f
�|����^ңJD���OZ���Mg�� �_g "Q��CPg{8a��z2d�B�?�v}�K�a2�7�4����?�A�U bYf#���痲�	��N�g_0�X���Iߏ:%�w�It���3|�/���o�(q����p"|؛]ƿ=���@m����;��-ա[S���yo��1�S���yNJʠ���B^���W�i��Wf.X ϩJ��hcQ9�ґ<��m5�J�#��T��ݛ��!��
�&@:Z%���+�BK��K6����l(�X��u�(ݝ������7b�ջ�P�g��Ͽ�x�@���c�䓴��?�o?G@¥��e��O6��#������U�Y��C�Xo�el���'t��Otiqa.���)8J_��l�#/v뺃�����g+c���g+���5�G*02�6��c�E�����)��Ap�5;�����ؔ��H��o�����Y&�=1��m�F���M�}�=G#��`b����׽�ϐ��q����2	q���v_�_��(��O���At�C�/��C2��W�k
�i�|/[6)�gf�:�z�;I�&�!��#��?b�/�������V��O�a( +��<*�ߠ�rz���9}w�e���m����k!���kYc띈�u���&~8�3]����g<y[ZQ���~�e�?!�o�p=�{JE���b>G4C��Mc��/��l��G�yR��#f�,%�����g"�Ďy�� 5�i��N��[k��W��#*��kNr�b���۩t]Zz���ݳ�
�V)���Wo�L��zK'�n�>��	��_k����%]8�E<�Xo��8+7D��n����jB�\V�'rRԖ��ZPԨag=gE���;cq���~6Y*�p��1�U���nބqM��+wZ�NC�j���HO�m�� Fz��]:4�a4����묇�5��dM�0R�W�1]b�4�T��v��:��r�k��z�T�Cu}S��h����VOyT̔��8�! J�ƽ�Bދ��I�:s��y;
"&���WiԳ|8v��-��[�!T�I${6^'��Q���[L�^�v��,7��|������S��F�&���2hO�U&m�6��@��Ĳ��AjT���A��j}��i��OP�|]g5=Z�}�^����:a��������{f���)� ��x����7]�a7Cj/���s�`Ȝ��'��%(�n{`�ˀiw}#Y�#񤄃�bS��J��]�f�2��a�u�Э��c5���\0r60&�?��{�?s�g��5Z���P2���4*���)x��j�z�WW(;}�mK�H>S;�dwd�q�4�rr���M��႟|cG�酉չwx��1e-������E� ��6��`���F_�x��g��]����o�GR�4e0�k���o}x���W{5�;��C�GF�:n���/�'���Rl�������j���r��a��`C)�B�/E�'~�G� ����Xi �湕���I�ܾ+�&�T�a�����@��>����e�����8����xz�Xz�Du��Fvl6�tY�J5(���_��RȰ�4ܪOp�S!�:r��M��ũ�5�H�n������v��2���.OuH����xn����Q�ϙ��w$E"�y�J���_EyU���Y��UDӎ�ED�;D	��ԍ�#�2����r�Djv�y��DOk��s��}(.vG�g��dP{��W�0�=�c�>��}v�C�a	i�+�uqp:j2M;�zɗ�&���J��,�)d�x����l�X�j�8ůn�����t|+��gSp𩘉Hw���M�a[�^���i��Pz�/ه�S�'�\s?k��N�#�3���٬qO�-��iӃ_��0f�B�]g��_����ʨO�����b.Y܎��
����A�pT`�qo�Ri�1b�����J��b�i�®MF�H������)6"�H�!�5*B$C�2zI	�#�|*q�LJ��4��~Z�O�2��qk���cj�8M3G�ӌ�����eg+��~:� K�X2筝M��bI\�QP�u�H�����LÌ���}�kxp��*���^�3����g�4w���w2�_��N���ḇ�	��Up$|�s�����bHBrm�����$2.c_@��򞣎4�~-���\ќ5i��w͗jPGTQ�0Fpd��)A����[#��g�.U�_8Bߛ(Eg���־��ģ�����LM�v�
pK�� �}i��Y#*���v�u��?�Y76t��̠g�R���{"KŨ�'�S���q��	����~/y��">M�`��F��,I��J�)y��Z i���k�wo`pl�,�vj���\�^9��#8T�����k�����(�3�r�V��N��<�`����#Z��ŅR]1�.�,@
���7�/�Q���"�	��Vv�L3sVQ毖s�r�o��w;��Fe������\�zj�(�VY���<�"zS�n��C��݋����!�+X�>��UU8(�^af*��%���M<��ޑY��0�.��jMW�)�=���c\�b]�f>g�1���+��>�<1�K�*�D���C����sO>k1(�w�M�E���$���-�r��f�Y���<�F�m�=�����	N.��u�J��c]�8�.�K��Xg����-_��&J_��SKS��*���Wv2�뫰?��1u�M�)\���Է]1"U6q�����(�sZC-�*礂п���g��/T�^{ƞ<��UË�f����?�"ס\���*�����eU��`�ΨBZ�����O	����;M�w��4�����!��o���çYQ�(�hǢ����?�a/��~�j�ߵ����j������cc�&�ʧF{R݄�{��b�mb	^C��Jխ�V��q�AUp;Gέ�^K3�(ݭ�z.�#����y���Pml��<y��Q�=���+z���MW}��Z��#���p�(ԯ���U�*"$��)�"�ԃo���O��Z����ݡ����~�M:dY9sȯ���2a_91K�!>��Z�s�q!��q7��Q�z�P��h����~O�DbWt�vX��K����/�}?|%���I!�ؽ��}�C����M?��!)T�0j{oRR�2>��N���Q�2��I������v��N/&T�)�GL�5�j���X�iA.�Y�)�Z��_i�7�"S+�U{�V;la��ޮ�c�3Bஂ�l��MOk�FA�e})�URC���1I�ۂ�q�OR�V�\/'���%��|��v��`��\E�V����	��Wm�*�i���v5�ef�Q�koC��j��h�_DF�cޖ�����+���S��)An#K��*�R�jiSF'�[�;�}6���³���9Xr��'wI�W���6dE^u-7IwH�k_�o��[+�D�n�c@��t����\TUr��e��_�ԓ3hF������w��	�ղ�h�45V7�I<"�]O�6vg�VP���_T�Yo�j{;i�)��AO�=��*�nE�t6Q�}�ۛ��q��$$�ZE���1��}ٗ�=-g��d׎PF����VNR���dO�Q���`6�(4���6�U C=��	����7�q[�E�-���=k;
/�4�nf�8Xd=���̬^�xW�iT��֦{�]R&L>�lUR(L�VS��Цk	 .���l�A�ʳ���>M��6�#�z��R�p�,�bE� �Iҵ���=�r<��I7D-T��s��X>z�MG�>j�j�O�+!W�0��5��.̝s�S��w�XG�Msp���ȝ̮3�k��j5ڽ/3��,N{�����7�ʏi��W�I�5�7s�:ǧ����=�|敏�,��]��L��~�S��;�h*�%�=�-K�"Yvh����ʿ�~�}ӥwh��޻�����_��S;�s���(�.$��w�854��Q�C����k���f���V6M��]���$�g�+��8xL�NFN����;�R1�4��=�Q_������=:<H�%��~�v�������x�c��Pݣă���hni]�|����+��=�|��BcJ�~����a~�5آ�4%R��2ZK�����R^[][�#��=�FE�������{���	�*�����_�Iy�׭�6��%�A\�Le)/a�9��)�/{w����%oR�)�	v�=�d�w���g:��Qj"@��:�O������D�UI��id�`��Xn���u e��@�����W�Wx�+�*�/@����g�B��Q7��7�y�W`ޓdƱ����c3;��蕘:� B�I{��~�~��޻�`��������X��l��˫�>x�Ζ�(\:�V�Se��pN��V��v���Uo���\�.^�yO�Ց��>-]M�$]�7zq&B��YK� W,��-��EmT�1�k������A���Z�88o�I.y�CxU�W0�5����z\k�|��.T��${�L��fC�r�� knQ�'T�5~����9TC��p� 6��.l,{�c� n�?���O��Y�E$�Y[��CA�J���%<�u�5�H+�>�����9,����7�Mޤ�z���f�����e�:�5��J8O|����2�=��kU� |6��j�XË��adn�~�����M�(�a���Pg��C���<D�� ����_J�U,�i�����f9<�5v+!�D���8������zV�[�k?�>�<S3�#��c;է�7��'�Z6C��$��u��M'I����(W]I�p�j�3%��R7웣d� ��_`�Li��|�6�sȶu� -�v��=��o��s�����˽h4�����_��j��t�!o\g��b�c_=�ö�D����}���9&9!P �Q�D���w���(�L+��׺�'�k�0�`��Z��8��(2�zB\©�2��)��Ga/K~;=���c� �A��~kdl�TT��kn@x���y���6I>8���)B��%3F�L�~���xAK�u�i��N�H�N�<��;�@5��~�q��?%�EX��0���ÿ�[�^����w/�D��`���J�Oz�����(����p��X��+�ȴ�toG�rT�6�%^�[R���?��oL�qe�rO��n�d#�7�K
�0�V���=�߱�	������q�KS��������0�-�tk����E ���+��&ʙd����ߓ�R� $f�ץn98�v�~+%q@,���U
d'���6�Y�����qw[B��%�+q�$��)�e���o�E0�c[���ń��R~-�5��*}k;�!v;j��ߋ#��D��3N��2�o/V?�V���8���0>��;�C{�."�6i<z�o_�MF��
&�0?e�u�&Z:{�e$�5g�K���S����Ie��O�Ͻ�<JZ4ISc-t� h�ROK�)�����M�K{*��yQEPH�K��d���s��i����g�x�&���k���r 7)1D�	1-ܤr�����N��}@�mQ��܄2R��ڻ��&�\o}�ߡ"Sk��z*c��w:�Q���=�ǵ��rV��#�D��B��ᕢ��f���ұ����Ϥ{��Tc�cYM��E{���x>??��5~�k��I|ff?��9����$�b�=�#!@,xzǖ&�*B/��V�������'Q��'=Q?{?�~����������h-{8ԩ����q�����q�K��un�斡���ESW���nC� ��{�f)�j-�� I�c
<���\�˵� l:�{95.��C���FD���:#μ�ߋ�G@H�ղ���'I{9{�PS��L ���K� �	P�:b�ݏ���(R����|si�K3~�յ�}`�zK_0�F�+�:�ޣ��b�R~-��މa��p��n��ޜ���V��aZ�����.��X��ҫV�����F3š|���%]�L�~E���B �֪Svg](��7F�ș4x�!y�~���� �KR��eﾯ$�=�#���e��Xk	s�R����� I�Ȱ�W���Q�§��Ԩ��� �(ة�����A`��t�o� ,+��-���E��$���ޫµm��m��ȼ����J��g����Qu�6VMR�����dH-���փ�������p(=o����~},7�_��`�7#���Dzr�ױ�����Jt��:3����M�UVdO��U��H���+}{H��g�]])��:�o5yW��n�Z���
~?�3���h�@���GX�յ�X|�_ą��M���k.�;�L��<�4����/�d�x+|�G9p�����LNu��%J����-U�
������ab�ELQ$^��G�	-�E����U.[����ɛ����(D���B�i�ߊż*Q��*x���RzA>����b�C~�u�y�f��?��>S���m�s/4+L�D�qRU��3�������ϬQ���e1/�E���	|Ƴ8��*<���~D/w���eumY��щ��ٷ�b����]k��͙�I�tnm�b�]����3�u��jjJ��P�хG���,{�ܛ5k���St����-Q�����%�kH�w�O;��!Y�be$�5w�ܷ^,>���ˈ5����un��O���.���b��}wc���N	�h}�[%��\4�����2v�La�U���lU��ն�^�G�O9,l�c����轹A�aN����B���f�I���6����1���������.'�3�L�ug��b��ř��6���*+��k�#�`�N���T������0�Ϟ�ƟJ���3}�����������L���PL����}�g<�	]�muϝ�Z��w>���ot׿�G ���?������ ���7ٱ��4���%$��8q��_z���;�c�w�?��{T֥�z�v)/Us�֍}H%��o�l��x�Ԯ��d���b���d�L�O�gB�Q���2���G���ņ^ʁ�o-�U
�����3��J�S�LQ��e�?w�gk��&���[z���o���� �f:X�$hy]�q�ӗ�g	�0�wFT�+�3;H�S���G��$����Q�w�"�б��Sj�3�NM�׍��n�&W6U,��U֨3�(����%���#�ǒzo/���Q����mp(z�+K�:�ܟ98�_Ӭo%3S���� *�R��V'&~mə�[�)L�1A���8+\��NY�.�9,RK�n{�v_���~��:�b�_`l<`ȤcP�b�dFUH��X��!/3Hf�v:l�p�=u�l����3��z�J�����Kvm��#���rgNe�މ�0�-oa�����#&����;�1�=CiZg�7-Gȓ����%w�����o��L�i�FP"O�Δkb�R>l&Etx�#�¹x0s���	r
_��X�M�S�~�U�G��zˆla������͔�)���IeD�\ pϛ���ޖ�����ΰ��H��g���ي�s]^���r���Kͱ�7��3��շ;9iZ���:<�]O�Ɂ��axY�5)r��ST����a�kh��.�,�u!<�D�d
��J]D��A��ڻ@魳��!E��7�%V'�l�_�{��������+>S���������i����c�8C'w�\�����/_x9R�⍌��n�xX����]��-���2v��� k�$��ML|�Lrxa�;?<`��j��?�2ÞƎ�hx���U����ͼ{��iM�ᑼ��P����
P-�.<�uBz+w��9���8~�۟��<�Sl0��Q�eB�7;��wT�Y�7�<<#*
VP��*EZ(:"�Q:���L�Pt��JQ� ��HB�t�AZBI�=$� $���� ��q�Y�;k�X�{_e_�w]���ݱaj�Q��%�'Iu���wi0b��a�+E�b��ĝ�_8/)3��7�h�Q�����Ѷ$�����sgGdz�0:���h�l��ώ�ZhM������f^���|�NQy�h����e�+�(�_��f�lV��[5/�������풬�nN�,�����ð;o��Qr�.��4�4��iΠzZ$i4���h�][u�'	�|[�j�ө�9:��Y�]NMu=����������P�;�D>��Zw]���?�z��m|Зc��*��v�����D�巍@�x���D�)ԩW����z��AS��H��d6`�q�F�x�5 ;͊l_��(Y�|=weԦ&KK�qY�����`����Y1����Ip���<�@�W>��N�D��>�,��3�o�+P�u���/��.�]ȥ44�}�Z���H&b��z+�m.�����L�Hw���v4��<9+�W�d�*E� �2�������]v�mE�F���Z{[�K�s<�� �K�n��|5�n����@Qo��-���f�U7�[rJ�Ԩ���$L��8}G1OqHFf��:-.Q^ѓ��?�?�"��,X$3�d��u덖��l��a����bn0�`lt��0��lx�:����������CX�x�&d��E����RH��%�!N�S8ʧ,%�j��x:$�:;�
���;{̬��ŧ�.��~����z'G��Z�W3�[C���Ӄ�^��l�|dظ��ʒ/D\�y4x��S����UO�g�J1@��j�9Z��2/>-��v�����%p�&��7H�#tRWɜݮ�;�K��T���gb�c7��������\���ni��Upi���^�
+Z��x�.�1�q��g9���ۄb��/�aĖ���2�WK�T��5����¦W�'@�qY�7��{����b�m�Đ�:��dY#���x!)he��瞇�e�g��0*G5T������:eF�+��Έx��.�;��7�<�f��*�Y�lwp��zZ��'�e0̊Y��Hv+�#��j5�������^���j�ZW�-]�$U�Zy$r�п���
Ez?c2�
^Jq%wr��=�Y���vr2�Ś� �ז�1��	s'h�-�͞����Ə	�s�4��V"'��p���/%������?�;��U��7��}�����]=��ld���C=�f�Kq���GZ��������;*�F�i��O�B����$ӡ�����!/��6����,�&���Е�>��&��o���\4Oa�9H�t',��77�,�~��]�rX�_bI�G	��X�4�(�e�����ӂ�6�Q�E#n�P/�>{ďt���M�w�~�E��:�l�t5��(։ڌV�ռ���{�z��-X�y1*7����?�oc�|��R�O���&_L��T�D4{&{'�\��;�T�R⺳�`���&�Q�6L̲ƶ.�b0%��-�İo��4�0h5����)�^>v�H�W��d،�Y����E�c�m�-�����.L������}rr�{(a�:\�Nq᷹8,G' �dbK����]��vw�j$�03-�8�m�N�Li)?�HQauvS��͓�<6�y���|�P���T��{��iC'@��_[Brs\,A�kbs��C�Rb�i� I��t|������LF���X�5�.܌ 9,��V�������nC;���7{�x�������(V�[n���|Bh������j��u��j�3K�ylol>�����kc5q�x���]yzS����n�ֱ�V�%��}+/V�� w�A����R=�8$Af�����t�,65[[fk�BR�̒��FPgQ�Eu� ���u	���(1w���-�c����¶��Q���o�%��i�-��I׌�!8��6��B��k�N?�����%i�jʒ�����%�'��6�'h5�Eɤ{��x&a��ȳ�Oh$狡Xu���;�J-�[�3�N�>��g"��	@��Q�K��c�m�6^"�1N����JR�&רȟ�T�pO̽P�A=�"
��k��2���w�0~O"j�{�A��9K{b�p�I�a�*��
�އLH���A\6~������6�N���.�T�b�B���JN�>/0�;W��8ӳ��v�i9�������7�0���r��;}ۡ����E��w���Kd�6���o��Ռ!��6���뽝A� 4�,�ɘ*�,��BP���cF�ي%�ʋ$^��<�E-
�Z�R�;Cm�R�c���
�p?���ufaH>���l;Xg��6y%_˄�׏x��A�Գ��JFZ��/�2�Ԅ�̓�b��'�5쨃�5;�LUh�3סg�#�H��ck�H�b��B�Q&bT]��NŹ�MX��V<KI%�%�o��4db��D<iݯydk�(P>�LnKY��;!"��4X6l�v9��	���G�A;����:�`�-6Ll|��;.1����oE!�yc�����=8��q��]���cA�ٻ���BK\Ѐ"�����n`h��V��	��S��\�9�*F�%-ĵ�.z[��N2Sy5���z�4(8�v�'�%R��_�N"��ǒE����5�	t�U�1!8�I��D?�~���NPLg�nyw�:�wڰ΋jB ]��R�aНB�`�q����F�I�aH(���|@դ!���5m%B1ld��Ψ��5�<9��<��lJ�]m&�m�6�3�^:{���P7��vʲNgؑ�eW���̳.����눌V9͍%jtT�+;#+�FԐ��yq��2�"z{<�,��e/��¸.�CIC����R��ؑ:( �W�F�p"��������B��"-�{�nkh��y��Zw��i|�v�PT]Y�� (�ejaC0{�qW,��zAX�k*��<�I_����֯uf��"i�&��S���0�;9v&�t�n��^�z��u��ۉ0�0FO��7W�s��#�.�u�"-fu��Go�
�2B����� Sˬ�5�u�����H��C����؛F�C8�ۡ��Ob�]�Z��)��R���803��������	���_��Nz�"m&����y���}65��*6���{�3�F�u�QØz�н~Qϯ��>��`�(����E)h^�����e0n�G�p�����i�&�lB9h+��;�έH����=������Hܛ˫�y�t|H1Nq�rWF�u��	��nL�r*+5�VG���,d�C��/�yb:[�x�1�r� A`���2x�{r���xs&CP.A�� n����a$��+�˦�N�JOp,*ǹ�,i�!�B���\���������V-�gp�PȌXߔ���I���`ހ�г�XB=3�Q�r>�a�h;jŸD�U������	�|�p%�$o h�+m�/vapS_�\:
��Q[�p	�e���6�x��4�1t�K@[��%@�L��n��@K"z&�+�i���/�=�mM���yxs4+C�-�]F��&D�z`�W���Έv�A��mt
1G���/�.�=\J��h�j5(��b���j`���}_K��]ص�Z5/W|���$q�:�
�`����m��V��Wc#�D�cZ��-��x.�ʩR��}��'%���l,���`g׎��������U���
�����?P̿H[�������ߔ�Z�~�5�P��e�k�I^�]z������I�v���Aʿ��~f���	R�v&wX�?�6)*X�&O����^\�&�{�����v�� ��B*���/C��?p�M��z"�	����q!�*X�猨p��R�[GX��Ϡ�s�6rz�ˀ�����bq�9�^p��ZeHF廵ۛ=p��;�v0��@�ءt����WŢ�>�n*�)����w^�����ڀ��M��u���2H<KXы�\��ݨ~:��P�6��ɄJC98�,�v��':�#�*��\A �(g���b��<�ٶ�ȧ+SCdM���s�)�x�Lb?V]EmL��>�|)�Lc���a<��2��
L�Q<���5~%�}�O��(�P?�������Y�:ٵ�6����@�}�Q�׆lf�K��u���EKRX�eJ5���0//ϭ�S���	-��	G�\H1�=�8h�c�5��U`��ow�E�j��,_k��'=�.|m�\���}Տ��g5�|�1,I�g[ɮC�Ê	wc����Z���J�&�6��i���RB��	�mm��|�Vf��kN�m@E5�ƞK�8H��Ϊ?+MTh�R��#��z�r��b�Ü.����WY��d�N㢂+��,M��DQ��>�vMsЦ�{����#>�u��?�WY�㘨G^"-�m���]+�ou7���S.O<�]�6�M%�BW�� \�k.�C9���������h�4�����r�E���ej#�#	��H�w6���V��/��!�� ���~�l����4?ҏ~�� ��LN��pB�m�QI�s9���b4`�^��E� ����n3�/_���k�R�r��zzg}�#m�,�!������'%B�����HB�� 2�h�M���8w��L�h��A#D�(���Cq�}c�w������&Bqy�����yx_9�w�������G��d�G=�.g�D���f�z�͕��fV��.�>*��w���\�>S>|)`z~��~&�7��L-a�]�����z+�C=g�����C�Y_��b��&��#�Ҏ�^���ŹŶz>���w���
�aה䩁[��u|(������-��鵅[�z0C��gk���<�F���I2�p����~���Ca'�;xxd�7]��1�ꗂ(ȿ^�}�[jw���9Д���"�;�<Z��q�k�k�B1�x0��1���l��4`�PC�����QF�o����=S���M�~�1B��d��C�)]��S[=�A��#� �_F�G�7��{��-�x�YU��X�<����#{d�'W?�Yu���a���{Wp���{���V��:��ьwR,e �$��mD���.t�}{K�(��?ź=,����s�� ����Ә��HO�KG�W��=>?:�y���x�g�Yw�h�T�~]GІg��������&�c�ѕ-6~T�x�q�U12z!����q����4������<�ժ����Q��o)����Z�ܷ�"�%��+�i���������e_U���>6f�W_֥�N���Q��.ķ+�wng��%Bm_����2�Ym�u��8�-3��kM�~��(�D�}�O�!�}t�孝�Z���)�c _��6��W���>j�.�S�Dj'�|���'}Ի��<��$��q��
�9Ӫ�1z�!L,Օ�����]��V���H ��E�ћw��{��Lz��(<ůORZO��O��)���w���+�8���$oس����U+
�r�^�S�D7�s�Y8�u��������wT��r#�Mk���*2�0��9�ڋ���un���P�T��P��o�z�������MM��{�(��~�����H�G�dɱ,׸���}�ȱ�b�*d��I���]��;�^@D��vO���~pujN1��]�B_5^��4�q�OYI-�~��k �!��I�U:e�v�ƒ��Q�\�>��w�]� ������9�Ԯ�`g�r䥳=
A	�M����gg�_p��r��O&x�9�X��g2"lz�mX��So�<
Q/Ʀ|2�dj���"І�E'���C~���+�	V�WPL#W)U�3Z���A~ rKʛ��Ƣ�PS�.KZ����C��[�f� �p$��I�ZF [��w�([����6�,P���WF2Y�� p�vQ�o_Z�nd/u�NR�¸�I�B�i�E-������)Z5���ɐ�������{���'�h�L4��/�"�y>ҷt�n���#����ƺN�Z��C~)2�m�^��6�OPڑm�� �%�|�\(��� X�n+��;z��Ф���ԟ��5�]�ҡ�Α5Ė~�p�k5F�s���w�o�)IV��W�C�]�g�-!@�)Ԍ�{�pۦ&`l�5.�.>4y/M�w衅\uNq��$�e���.{�? �����TQ����w�b��8�9yJ�/��#J���!�~��=�~9���(j��7וjd�!7t�h���&����Z��  �t��:-�sKj&?A�MS9:J���?7�`n�K�o��D'�`>�ԟ� 8/�.����E`����_�&7�0���h5������g��:�@�N:�n3��|�qz��BG� �����00;_�bJ�kq�åC�`%�l@�2ؙ�3�g���Qנ�n?%Y &e� L�Ia�t]�mfc�%�@��^K��- l91&��/����3�7]�4T��jK�z(�z }�t���t� e�<�+��M]�b^��,�)m�[x��>1D�Y�v���:(����m#Ȋt��ZY ୤���~'�,�c`�(*'u��k�ͤP�{Z�����2�[����(���G��٤H��x]L�(C)���^}-�s�̯3O�,v1���{�/>��%�k<�1T�U��X)[�,�.G T��N�P��,��Mho�����+D��W��XfD<���e�۰��y�`'R�K�	6��(��0p\0�����{  ��5}a�伝�!c77�v?X�V�}C@�XHt1��s]H��0���v�=�V��t2@x�^�:T45�W�Z!^�U��a2���
�?}St I����.1Ǧ�e����e����놀�f�ѥ���}�ȗZc���jZ 	�x,\	��=4�B��؄�~G ��;M ��0���LM��Q~�X��`a�m�y�hf����wޚU�r�̃H͔�$�k>�3ʳ��4��i����ʀÊ�E����)�[�gk w�'-J�>'������g��t?`o^r֎O��(V�ō��  �9m�[,���C�	$r�t;��k� ��9#[�z��Brl�M�1��j5���н���w9L*aV�Y]���E������KU>��h}�vwW�􎇺k&3&{j��.�W�И�͗���ǔ5!]_S&����&��hjG#��^��I�ۅy�Z�G��;^tKJ��P4@͡ڼ5�KR�	 F7�=��	�7W�L�>�la4�~����B3�eg������z�{屋*P�����^0�♸9ͪQ"��չ;_��)�D�Q�����K� h�' D΅"�d�G��� ������ő���'9��p��Y;M�e��P�IQN~A0֕����s"E�ʅ(�.^P�= <�F��.a�|�y�*6lcN/�˲�,~}X�Z��r�M�y�hgi�;@�g��w'n�����B��^��F�=�0K���;�-�PMe�yT�*)����pfV���maDanc���҄�6���+4�e��KGw̱�3Tp��kO
c����
t�M�]��ʴ��	�
d�/��x������m
Ta~c8mJnO{��η��v,nSY*�I�%ۖ�,F�q^,��~w���QM�~�K�
�T���T�@� �P�d,w VX�l0�x.|��a��P��22[�35��K���/��4S��xA�r���vyC�2<��X��"zV�zp��q7���}�#�Y·�?�i&���\���`4�]v;�E�	��̕"A�'Fc�vr��q3n`Xq�Z���(����⧆/O�_����]�������wsbH�vO���u��B������	du%�l�kh6'Y����V��-u��$�`�7��Xo�"A[Xi��d�o ��t_7΋F2>�A���6, c�r�hfE��fv{5M�c��Z�G���	���Rx��Ii����9�hjl����/���k̼Ak$Ԍ�L\�À�IN�L�Pm�xN��r�E��ȣ�F�_�!��w��$�B,3���̛�	U���Τ��U2��f�:W�!��n���P�+�(���������n�k"�� r�e�ʂ���EدXK�N+Kt\ߞ�n��Ҹ���v9�a'��3c&:�*�6�3�=պ�赭�fZy&����@	�:���jlP��������-�>�W�@x$�$�]{P�ڍ���QY��0}R�-�VH�����~Ҟ��W��YE�&�8�8ɹ�I�AS��&2�b��,Pj�<��O��dT)�u�-�w�,�[nJ�� �n�T$��/���c�P�Q>�<��ϯ���.h� 1tM��2�d��w@��5�k�8��h�Ch�jO;_����㺙�/��/;�&�V���>ˍ�W��K���w+�s�f������i��A���!%	�}S{]�o*bL}#+�sVΗ�Rc�W&��N
�7\y1*��K���Z�}=�^�#�M�Y����A1�}ۜ�T;�1�{�����\��<�#�^�x@�0���tK���sCA8����Ws�o|K�6xj�M��@�cKoל���IG|>����1�}�C�KlTKʡe�%S���$g�@m@�H����zLA�d,�|�>�Z�ԁdyA��1Kd�@�Z�R+y�l�	O���?�;�f�ܿ�T�s7#�CJ���A��*��9H���"�����s�����ԡ�(z4��&�y/��|N��<����n�/xd��9�F`�Mѥ@��(���x�0���:(7Gӷ��>��^����\~�Q��碛v��V�΂9���Ea���lR�Z�Ĩ8�$ A�M�9�o���ګ�VX
q'�@��ASO��7qc���&�<��$��g���2
�i�a"A)p����e�_9�0O�Z�{��ZM豂+	�&���������{�D��0�z�Y�ND�X�K+9�|t`�����C�/��o��rq`�N3�s��!!]��¨,B�,�/t�=3C�r�:��ۢ$h<	�Ƀ	����$nɆ���Ֆ��g�4FJ�Tޖ��t*Ϋ�����ˉYk�K-�� ��۔Э�MZ�5�5*�A[�z���yb�}�K�� �9��ëp�狴�E�p)�<�?��Z��E=�������`BlY㐊E�ح��aK4����-_8v4FB8��j.@���M�K���oJ��rzv Ԅz�`��IgՋ�r7��)Z�$P�����^���}��ܭ�w������D\�9]<�=�yzY�H%6*��XI0i�tqHB��I�jcm˝���.�w�������Ў:j,���k���q��{E�(AZ8�����A?�T�������ɝ��Ob�o�s8�x���Q�Nթ���?cx�>x\���xaT��=2"�v�Y�'��SD˫T�䰢�ReI9�K6�GVS0;�(_
�a�����dEO�?_�˖�'5\�veF�v�20J�>=�Q1;����iMd�v,��
��^�3���{@߸U}�{A�X�ߒ�U�Y�H��m�o��/�p��M��� �z%���޸f�ps}�Y��'��J9@�Kɋ�Ui��zW�|���&#ݜ����Wt��1 ��	��
#R(���i�(��!J�W׭t�Za]W���9��	�Χ��j�(Mh��f�<�g}0��|�1o��5�Gm����+�8�� &��.�<�p��!@���5ԌHW{���!|��!�0�L�6�yBL�c���!�/�T��^d0(�Ŭ�i�W��.��΃9�������"��'���C2o���J�1�-�[jC[�Ӄ�ea������dYN.�Gh�������)�'��;��k�b����W���C�ȥڙ2KEV'O��������Y��<���XB�TW^��6W�\�4�-��!���31R���琢
%S�1�)?��h^�N��(����Tx�U��.��KY�C��8��J�U���]��9#�Ī0�Q���K5��֦��%[�#"�1i���τS�L��>�BsS~'�0�Q܌�����@��F���D����9XKbg����Yė�1��hN��r����M?+�i܅ī�� ��cΓ OF˘>q�j;c�lx�Y����9�~8rJ�Rb,�0b��7'��Cwz�4K&8��}߁lf}P�o�����~��"����
t��/?�%K�I�C�Vל�&7�&�(���7{���a��e���L.u	p����KAW��\.*�-�[�r��d>����q��n�m]�am��L��"f�h��g�����A=��9(V�TR�Te�E�C�n�ԃӏ^r??v�N���wӇr���o��/�����.pu���Ts��:���th��#���!k��q^Dd�����v'cq��;a�u��]��O��.��n���`|�<���ӥ[{�.�q��zwi��%������,I �Pԯm�F�H�3@yn�#�����jG�P�r�'�]��\N�(̃ �?���lm�J^)_�J�6�<����i*��j��K�Ksy�r�(s'��u;&��pz���ki��R�RyKc�$�$�Dت�%�^����;���ȱ���-9�rP]d⍏�>k�Kz��߽�����,S�
�6�X���$�������4^��t�"VM1���G6L��m�{�ꈿ[vz�"֢GS�4
�۞��w��Ud�B�'%��iL"���:.ثQ
	��#<t��߅Y[�(2���xu�e��Dz� ��Ӎ0	O▌NC�;�S[8J�Z]�M�[Ec�('i����Ĝua���k�#����G<>2h[ZG��2�l�|�Of�;�!���c��R�"�B���]��i ��6M%	8�P%0�k�TD��_����Aw
�8���l�i�x������p׸��+�ޙT��.��>[�����&첚yr�\���nC�*��"(��p�H�`N��\��u�i�]Z`z\����!�6��;�+t�t�f�������Tn�~�$A�1H<M5��N���q��?��`@y�N�C���s�j ���.F�O8ٰ�a��ҹ�Ӡ]�ql�3�ο����9T�p���=������S�&/cI����ᚬ����9v���>M����5����=�Jb|(�wYMY�y�tn�r�(9�#H1�A��	���o�0UW���L����|D��<FVxd��r�a�yQ6�X1*�Q3���s��uQ ����0v�� ��$��.���d�Yb��xe�0�W��c�*{���(gW�F�/�ɰ�e1"b!签���Y༤+0T���a��j�zx�q�sUiq���jy� UI� x�M[.6"��5��]��t��p9��h����"O[��N#F��8����hf��]���Q���(T�e�`�Ĭ��Wcv����'X.�*�S��*�����1S�%l���%omjߌk��Q�4�����^�Mл>�震�U�k�Q��1�J��\�����jp)I]>� �7�nzz�Eͷ]E�)�H����Ļȅ�dB��E�IFT3�XD��vc,���T~��0q.^�&N_F?r�ې��Ww��ox&��W)}L�<�k�(�T����_Ff�;�f�/R�[ݥm�}~}bA�D5���ԛ��Kr5���
ȱ����̟�]�(nQɮp�B�y\��m�ƈ�q:�(�S��f`�I �g�Y�s�^n6���g�������WH��2v�n�I�^l�,��yĴ���고��f��a�BU�� ���J8��esq�qt���ǂ��������}�	v�Q�C+�7*�� ���}H��0��.*G��'%r`��B8E~����׽������]�g2���?d��l���|�� ��i��\~�p���I� O�8k9J�<p�t�)��8w��U ���%^{XԼq�UPͷ^YY4�E����M[Ϊ(3�z�|A5������IL��~�K�{��ȧH�� �����*�ٚͶ�M�W�{�5`(f���ڣ���ׁ�*ݝH���B�Ns����?�6qT&�����a#�	kS�������U�%�\�H��C��퀜���̠��k��>�)��@=e��V�����W�m�Fǈ�T��[ʇv9�Ԥ �W=�b#b��[>����Pg�7�+A~#�Ź�Qi�ZyH����i���e������%��e�$|T3-�`�o	��3b!�I:�s���ր�bF���4ʜ�|�ƱBa�}O?n�Y0���z���tT���bZ}�����0,���*���NPu����	����$�M��Vx(����m�vׅ�dI�?<')��n�݆{�#5>yu��Aqw�ecc��%(w���'��A86Z㔣@�롴ŭ챹t/({�G��X25�����i���T����������tϱ�̑��u��)��8��� �"
�N��މ��ݧSqq�%t�i�D�0�ڂ��`�_y�7ԓv��-�s>eM.��8(�zo�6��Y�IL�?������k�z�{�]�q��PY�z��e׉��^�q�����Ⱥ���yo�8`�_B>]ѩ
�=P���k�'�unp^���5\KS��=��t}��ړ¼k���݅ͮ	>Έ��K��H�I�w�,�q�����e�)�l�Ű�w`b����bϭ�+��g �T9��ݮ*A�M/
ɏ�%��7���KH/w;u��Q^T. T�z�yS�F��͈�w��?Z|CH�+��2S΁(��y�v�����7�[ٹ� �M�[�~�O��ޔ��M���\u���Č���[Q>���a�R=�5ӎ>�x�p���_�tx�ia�|��������!b5�_8ޕ����"���a���N�G߮r�Q�]�7U.��l%\���$?4�N_v�-6<Q8i|G�4h�TQc�8����Ս[�ֆ6�_z��3d>!;�>z<�Mz����2�%���v�=�Χ ���(��;�LD�L��h�R�p���� ���*��"��/or���b����:��UR�����Z��O���w����R����wew�:oUy8���sC��b�,O�|�+֘���Z7�a�<я��>N�����|T��y���ap&E�1�BI�~��,���a6ÍU/Z�s�Q���n�u��
�|���:7P�]��1{M��1T�=/Q+���_��CZ'�Y^�>�?0"���w�4�O�xJ藮0λ����k�K�1������-��T�Ae�F�GFĳ�ˍ��&:5����v��[gg���Ptڷ�;�������}�)�4�hD��:�8d���'vA���}��Ȓ#�,�7�!?��GG��w�@�`Z�ŵۺ�!:���k2���m�����v�_�3���,���V_{��t�{VҲ%h�p��Ǵ�O"�c�.���cF� �=��mIE�޸k�O�ɁR�
�@|�)����G�0�x�K�&�]c���S��D7�2��N�����Tu�����5�sַ����&}n�/�P��"I��>��J��L��>s�+�X~RK�]Vë���>�y}G��G����q%Ճk���p����9{���Y����K�ǃLJ���x���㞮���C��S�[�$B�;�'�sc�ϟ������̧Ge/����t�E��9�{���1��g��EOU�ܺu��W��؎�\Z}
U�On�T:Aذ�����ɨ��r�c���������;4x��?���h_��Y�2����. ˜?f�^l�VsmI��ۡ� ��;�?e��j��gm�����,�"Nk�ZC�㖹�B������6��0W�?S�g��L�>�� &}�\-7�����(����7c��;m7Z�!����M�#E�T���$@-dg�7dn|�K7��#N���q�������g̕��v�'��d��Qg����������Ñ�e�Ѻ�.��r�H=t䟢E���м#���q��D���ŕ�.Zs�׏��.�gUm�?��;)x���骧ǿ�PС�'��������o<��:�y|}
��v��1�ŘU�5���]���N� ��$� �"���H��r�a5��ǫ�^/}��:r�,}.�.tX �bP��Q6��"�Z�Ǟ��O��V��kՁ#|@���q� ��G�1~����3���S�����~���J�8g�w��{Τ����H���t���o���1R�}bf��7��*�H�-��k(=�#�>�\����R���H�������]�,u-�P�;��Nj9����v}{�R�=���:-�_C��^39����D��^����?�rT93����
���S<���zn����#y��[m�4(�A�3�DsH�@P�#C��O4gG��N`\!f�Wӟ��b8Q"#�"�e�ؗ6�Y\�������1k�i�_��oH����6Iќ�\y��SK��':w����>�*H� VL�7�,cq��?�ų�p]Ra��D��xi��Y������_u�b��~���#�t�r���Ma	�\����n��^���*hM.�=��0,�W440�%J�x��;1��-Wy���<m�����j�|C��E���l���\��:������wzݍ*=,"ҵSٺ�v�Һ��W,&xb���A9��k��c�Q֣��S�S���	A �<u�XW}�;�����X���Ek��ȴ�K��S�TV���'e_"��/�R˵o[�C�+�pAs�gba�x��]�/%��!c��^\ǌ'Q矸�i̜���!���=RSU\���2�R�\�9�T>���ߞ�Z���a^MC����j���>a�Ã�ŭA�'3��3L�򀴓�߄�ٸW1da�O�_���F�����3P��_�~u���R8ak��ZWnm&;�.�w����X�����Y_)LP��	��k�{e�nH���&�B����xJ���T�~P�#��q��S�S�<m�5i�qv$��ק���Պ�PH�J���sc���U�$��%�5��y�:�^��K�|*��7*�����ֲ�g�JK]��v+x*5�вl-	Gt��Uש��*��K�e�L������r�]w
1R1*��?�yb$vp8 *	u��5�	�L��(	bF����P�."��k&?N�4<q"�2�w�D��ͮR�$�w���ʳ#л� Cv��~)���d�جy vj���ņ�`V��K_Oj=q���}��M;��粔��eP��l�bTds�Z4;f���9���6�h�;S�^�5��X?'�N�IE\H�HϪv�s����4޺�cM�{V�:�q=�
�O��r�>���g�B�B=Y5�#)������n�4	&� e���UW�+sLn{$��v~h��Z�/��(�ᳶb�,����3H	�<�)�.�{��e�����M�iZ����$�j"ً����ol<�Z�%\�����%�_�����GC�NL��2T��(&�|(aG�[�V����;�����E�D��]��@� H��u�ʱ+V�	�|��t-+�����[[ۜ�:����y�E�F3?ٍK-2]E�Ҽ�#�̾��s6��6��DIY/Χ��o�]Ag%��	�(��5�T�Z�+V;��˚{�X׀��b�c��T/�RH0�t��˅9�+��dm+�@�46Z��ц�Hz��h�V��2�9;=7=����T�F}�JLd�ɨ�P{����M�+2�j�dw&2q�ڼ�ZS2��@��M9�LX�
��9�����!u��Ov���j�%�sM*����@=��Ft�fB��X�t��6�����2R\�L�a�_yl���__"�K��nm_c$D;���(�B��,�i�rM2r-����ދys�gQB�H�r��b�JG��,ia�:�Q��mw��]��㥐������G�� ���� F����k%	�ф�}���0���P�W8|c_� (��eI"�0npL@�吵(Y�^��m�7ܝqY�YK��hF�΀���S�5������%ӄ��p�S}%��������0aQ�3*������%c������oCI�и�����tw�b׸�Ԉ��d�y���Z�aD��&O�&�#��Vzn�T�F�FT�-h���a��9�ξD�͟��Sw	����үq�icu�_ iŞ!WC��Z뷩�3�r@^8��R���q�[��?n���|��P�/L|`/�����bj�^%ڜC]q�
nl����jM�VoG������-l҂t�H�ͶO�_'<�cj�F6_��T��珮s5��.��A�!]��J��m������̨+iKJ��MO\~y_Y��"!���kTZV�zZjj��5}!%曇�w�9k��J}�ۑ�t�0�j�WU�\��I�R�Ҡ�K���:�2݆��$���^ʭ����y��8.���u:[@�f��p�׬��]�F��t���s}��n;���p�<���H����6^k
�>
<���sg�/��ϵ��Hy��4q�R�&�♬O\�a�UsZ��X�O���T�D�A�#0Gq�S�F��Ћ��=�L.��8�L�VY���Lζ횞�@�{5_�FFa#7u���chSO�V��>����w w"�,NF��,j��??`�
Z��+;51�I���/o���:�v�����{P��\�n��9�62��~2��{	"�;�oPh��)�[�C�����H�Z�!m`�G<�uL:�����Fc���ɡ����ɩ�_�)e� Qm��D��ʡ"p���X:|��5��
�!QߙQ��(!>���&�Q�gQs����4���	���H�㢺���۾��A��s�>&�_`<O��(B;�i��ݡ�<�51�I��W��=�ڎk]Ea'0n&$km�#���Օ��Aas#��˽\�2deH���X�I����:9�^�֠���UV?c)�;�"�`�5.�+�][����-x)�]۹������y.���L,D~+L�O����C��.۝E��@R�o�Y��7>A!�5��*R�((���Cٗ�L�� �k*��I�>�-C`n�酋�0��v@�	��R�����1+}s�G3O�Lt�7ȹ�4M뜷i�J�����{G5��}�x8����"�
(M����T�JB�5B�MS�J��"5��IUj�5�P�IHB��.�>[e�q�_w|�{�x�p8�bΧͧ���5�2�+��Lhka�G�t}Z.E�B��r�iw:�S0,�Hs3�� �������z+���y~�2ݪ�ńЛ��?V1o	�k�����֙���h8���8������>`B�})��H.�L"%��sS�l���U��}̪����k+�V���L��<����6�k!��|���߰��˅�=$ο\�k�Qf����$�J��4[���~ԟ8��Q�~2�/=�U�B�I��/�E̩�����!�LA�:)�~�-��% ��$�q�i?M-���iU9���S�ʑbb�1��'�#�2l uFś��K�{��K]N��H������4!��i���rq�-ȯ͆d�����^��0t=����p~K)�W B1\
q�t����'�>#�z�(H@ҏ/-�a�X��㆜c(����]�u�'���$�d�l����A@O�D�!�ȳ�)P�ӳDw��O�
4k I^��mј���Ǘ�(�1�ڏ���H(�d����'�������c;�r/"U��Z��׮ȃb����9��u,3�Ғ�N�pb��`"B�%B.!(q��h�i�%!����O=�q��P�P�#�^�}/���@}`��F�bM��8�*�s���Hi��e���N-qT�v�ke.5�y|H�{���見�4�G�};v�`�c�Y�Xh�BJ6B�p�;
�>a�	&?׳kP�=(UI�+�뫐���<�V><��\G�q딬�Ʋk5�nT�E��^)�e�|�9L88��q{ލ���}~B�̫M��Ő����i�}$T�\�0ݐ��/�0�l�M����Kopu}�\��f\�%��e�J�/�d��!����Я�,7:�!$"��nD�'��Y���>�*���Aγ���{�T�A*FL�@��x@C��-������Đ��N_/3Bd!�F��8 �0�ϩ׷�is�&�Gw��,>�����k�1��K-��{��r^��0��l��Y���2��g��|�t��������w$s�~�%�׫'�>w%���?椈�技�O��\����v�9Un%ÅC�7�=m����.]��l�1��W���6rM`h�( z��XQn�j�JM킑5i7<�	�$xw�&���.F��Џ$V��5�y
0�Do�j��}P��ĺ�J���IXcJ��n:N+��B�OTx-4�r�3VD�>1��J��n�Cm�Ł�X��*݄ �+i�,���X�b��1&S�wj�u� }�H̙=���o�����,�op�kk/=�x,U{�r���u<�	�= ��Z�^���4B�zRX��tE�*{ֹ�־�jKdAp2?đ���Voϰx�X�{e��y�����X���Hg.\���2��rc��GL�kx����)��Z�^b�_�M}k���,�RW�@����w$I�w���:
��J<F����%��HV��6���Q�:���A�쯭Sq)Pbi��@3_:`�Ur����K�)�ɘ�^ݖ���DK�VH9JO��h�q"@�5�QFU�N��>����Ϳ��&w<r�vV�T�D��%�D�قFҧ�\�h��o���������,AZ"��qM����g���M��mv)]Ũ|��ϋ�>����a.�����ģ*X�rl0��1�=K�D:�t�od&8�CFhq���V��GS2�)�!$ޟU��w���-�m��V%Pov�=!��g۾�=�Sb�p�u[��e�[� �I���E��Ab:�F�Jw�������ĬI���ӆ+x �ĵ��UNv��3����k3�l�I�)ʜ�;F��P�lEhåX~��+�h'� ە?�w|�X�j���
m��2o�K��}�|k)��=�/'�Ww8���/�`9��i���W��[q���5#�? 9��: OL�Ǥ~#�:"Z��J��L����鍫�J]����M\D�m�[�þ������a�
���ɛpfs"V��{�[�!B�G�q�i�!� �{�)l7��vc��%�)����I�__�[[}�m|)r_ze׹W��F=�p�����Bׅ�!��<����a�|Jc��`�͗%�ʼ�߫wWY�mm�)
� "�-����H!�v�	lS~�Ǘ��[�!%����5��ƥ���T%C��+�؟�"u,v���Щ ���C�!�G���ī���Xv=�,R���aP�D�����A�	
/G�=�)|ֿ���.�v��e���~h��  ��P�+����bto�f����߂�j�ku\S�gT{K�v�nv�C�v^`5U�1�V�D��zX�!��EW?�FEh
-�E���\&Ѿ_^�&Ͼ��	}�?ɾ������<���D�<JR�z�+.;��k��m��E�/V�5����p
���˯/���@� ���%�ǜ�Z	�e��a��+���.����? gM����/ u�=��s�� ����4����������Ə�_�J��M?�F⺭$DS��'��ѡC�ſ��M���㛳�e�U	g2
z�h�K�g�� ����n�\���Wg����;cdd��XM�u�a�z�F�ֱ�o�9�Y9�ԡ��2J|4&ꎎPI�?��Cq@aD�7 ��������Եoov5����y�YͲ�&�)zW�LW��p~���A��g}�?;�7�	e��ubK��t3�ht!�r�oh �d���Θkq+��?�zY;�UZ��&��%,l�g�5's8�b�Qߘ���3:���"mʭ��oQ ��ugߑ��X�b
�߹i�����<�ϥ(�E)�ͻ�Y���F0��1~U{êaB	e���� @󜫋�cJ��Jl`vW]����X)W�M�moۚ���Ur[��Іq�������7!������.��k����'�� ���r�sHX_�?; `�K���I>��ߞ�I~�w|4f3Af�С���3t7�H?�������Z�-tJU^���:%
u�I;`�eZ�ǘ�13k�5�!�-Z�������B���GI�^{;�Z���e`5�
r����~�e��Y�2}�|��r`樯҄�孬\�Ǒs�su<�RTT���4h���~î<1
a�X'u��Zt0��گy1��%�s\5���Dw� s%F%�}�����,_���򾾸��r������:Q�U��\v�	?�zm(�s��m�Lze�� ��<�Y�l$�09N<�rZvA�򓚧&�mr	�]op����ؖ����),������3G{��u^�Ǿ#ߒ�j�Ȉ�(�UءWO�ϟ�ZިU�Z���,���s����d�s1��G����3��~j^dR������H�٩�:���3$ރ��9^��3 ��^�;v�vN�d��*��|ǛB$ħ��V@,9g�vf�ZP���+jNx������;9V�>�k����B�7�w�(bC� �L/	�c��f��D!��98Ny��!Hʢ_�C�s�t�@5rl\�26JU�$��`c��C���G�d���f&5�`1&��9��� �(hw����@���P*lnh{�J��vz9̫%У����K���������T������Vf*�hY���]�7OZ���Qt��IØ��G�;�vƈ�m`�ȷ�7|=:���/�My������(w�jώ�6�: ��`�6=q����g�����v��[�9_<Ro2Q�*v4s�
�e-��[Ԏ��Gk��K��w�(A�G�||�d�<���6ޏ��T0��iZS�7l�����t#i�s㾵�I�9Tb�qG��[�|M�N�p�~*׹�����kY�p�p5FК��#��xj&*�z��~Y�Lv�ȍ�铐�ҳ�!P�B�k�fZ�k�`� �a*T�E� Ewٔ�f���s.�P"�t�
�����������%��qG�j�;�'&q��a��^	2���TR��I @���m7�M�W۞
�`�wA��ϱe�X�g#|���ے+�%^+���KqF�@�ʳԒ������w?�ׄ��{پ�z�>w�ԏ���'j��C����;�B@Q�J׃͎<Y��P��r�}��{�����ψ��7�B�����qɧ~a�@�R��m� �羠��.9��6���v[���h�C�P��_��0��"�M�{�e*#/�W�e��
k1��Rz��y�E�G�S���p�(�Y��x,CIK���!���.�]߫�o�|�3 &7�f#�SD�Wm��ܶ��E!F����� �K�il���#9��|�n�f,�N���s�����y~^���->k⬍����u�o���A���ͯX�*A^Xo�L%�,������%y����:-�F0�F�3oH��X ގu��q���e�Q����O��������HD��_) ��>�X�}�aO����3{�ݘ�E=�4��0�T;�`��y��o�YՃP����è�7vf��^9����5m��i$�?����`�Vj���z�@%a��=�c����Fq�:[?�2�m�x[s]�}����[����
7�����D!=�oب�^+%���=B-Wעӫ�쇫$-"�\	�Jb��1�o��0�1߶W�z	b�q�f��G[�1f��i(�s'I�/}��� Yp���j� gnÓZ�<wG%���X��+/��I��'��bv�H�����y�ԁu�:�$��硙��/}��Dݝ�ӍeN;�WFi��D�!}�@.UA}/�Q�_��{_��������� ��Q����8��m����b��Dַ8��M�Z4ql�o��.��-�����Ę���sM�����՗,3��{;�n�W.U��ۑ�%����"M��H`F�4�&׿m����r(JP�PK�� 8�X:�ߠ���m�v��Ό �� w�"��Z9'3(p�sW1�`x_A��z�z�z]�@��v�k��f7�����Ef�ʚ�^S:��8*�?%~0h&��eos�d4�=�A���5GOmKXT~���Z�VJ�ɍ�u]��cq��v?ہ��`�(��@g��ɯ]�H��8P���C�}{*|�ѹ�(u�?!l���R�K��3���ȁ��L*w?�6�<\�����ԓ�'P�1$��l��5&�a=H�XmPW�o{v6�66���g\0dаj�ݬ�PCŃK��j���' ]3�c5�}�Pe�����Wt�1<���F���p�=y�x�´�ka�����l߷T_r�Ha
��r<h�f��x�3㿙/�M܇�@9�vV�f�n�%��:����>gl��xAc�����Q=ح21s�-F䚀jy�U7!͏ˍ���5����P2oP�X�w5q_֢ɞ!!�(3�	�\��|�,#F�W���t���0٭)�mI�k�t�o�",�aDLU|z�����1��¹F���Ċ�w岲�E	��9��{�IdP�( �GS3�V.`�X�����>leD֤\IІg���e�4X�������\LZ��e<F�7�c��7
f݅�,4K�btg�Z�|p�e�a�ֻ�tA�~�3���N�������7��q8:i��Aa*vS_���t\OO
�,.z��tg���
��2��f����;%����n ���pۿ��3���	�mD��׃Z&�*��%�ԛ�a�)̐��EKgB�J~yAy�%��
���w~B�$]��N z�e���M�x�7L0���P.$�sI�H�Ȍ���B�D��[k��6�x��U�/�|i�X�E��0����r���@t[��|+� ?�#����&��Z�yZ�ȨE�fx�.f���n��`7E�ѱo�� `&T(C�fg-Bls=[��nvx��w]�|n���d`�@��xbl����~E��u�r�M(,V)Nk�����a���a,�5���,7o�!��E;�����c���&�Ҫ2kX<�G��X�/qR�͇{-K�*�E�Y�2^��f���@ݔ"O��cW>�r$�h7�{|n��R|+"MŠ��w��'�Dyz��L�\����^��U���"�p�"z�a��9��ӳda�s��m���#Q������78�؍�@��{a{����\A�p#�=�<u�SKQ]�:����v�����F����0�]�]��F{�����t������A�z�(w�i9jj��?x�p�yY�]�~�b�nL��ꋷ�����|�s�5��Uܱ�5�w,�8��`�x "� 6����O��<�]��f�`�ePa�֛gP��k%u�7�����'�@�5��.��rE�De0�������`��X1�#���KkK�d���U��N�*�՝f_R�蒁nvc�1S�Q�+/�6IǷ�~���ߠ>��#��O�������v�E��{ZH�,7�1�s����|�mt�:���!�(?�%��U��lpe��V+��S�I�ΐF�A�=ʱ��o�6j?�O��~,���mbu�s�W���+$հ�JQ�ff��'���|;{5�ّj,w��s�f	�����G��ט�qN�Ǉj�v��.8��<B�|�y �����t�K����jnv���U�� v2��z�z����Kx���i.|�Whm�.�����rFv2L���4x��a��N2�!�8�Q���Χj��#��u>U f�Y�N��+,%O`�sJ��Ŀm�,��6v��")Ö�g�'���`��}�KM�^" |
����b_ly�困1R;,��V��Wk���<�a�D��᠊T���V:&(ѣ�������d���1VD=^c1��ȣ�fKH��E� ��X�JFVڔU~ed��En��8r.DH������B�� L��$��خԿeV_��h?�E�ت�[Z�2go��n$�L��b�$+3���4�[�2[�;�� 2��"�K�Ap��%Խ�b�l��ÆGv�C�U�]�A���U��@�Z]��ӔD�����pWt�5���j*J�6GL��aZ|���R�ĸrI�w�.	|d{���G�JKyI�Fm.�\�b^�J���ռ� m����W����4��	����o�וP&D]9�h��h�~�޽����0�L�
Y���n�2�uwB؝���u9B����2fI���b�x���8���%��B�ƌ���*d7���z�H@��C�� � �M}������i�x*}/�*X�W�0o�*>�:�C�b����Q�{��(��	�XF�d�_��ٳz�jя�2:�^�b�N�x�n�NeYAU�~2+����z�c�`3���d�{�L��դM�a΀-����f|�2���yij���M���I�sI�
>^ݾ�a~��Tu���`�ࠥT*'��ϠL/����Ȉ:��y^�P���ያ�������ݟl�?̒�E�>�צEVy<�^�VGe�)w��/v?���0����	�M@p{��PW#�Ƅ4�9�TO�t�;�Dq9��{��ñc�����v�ug��*7Zڀ��*���<���IV�nq�be��;�ߝݬ$��y[�d��lT%���Ae��W}�ׄ��f���]�<G-:}�e+�����A��,��f�$N��QK0ǭ��C�3#@}&8���~��´�5Ş\� ��ڃJ@�(?Ѓ��_��p��"LBc� �&yh���qfpCQ	�C ���F��P�{�xk�,��\&�
B�2�N�cJ䫎��M�-��x!�)�P�i����E�C���[>H��^��j8���"������Cc��&���yr�?Pm��[�gH]���a��!3pąBN  �E�H�?H����������S̠���s:ˆ�UX���J�~�6��|nJ^�=�z�PEQ5�a���&vw���0�|��z%�
��p���&t���r��am��ܚ�J�iGγ�
1`�j�!�T��j0����#�\��o�Z�!�vD�>?���Jry��kY
�4@XwD{��6��g��-���>�i7ZO�+?HM�������������Y7J�F�Tuv��0�҅x T��-l,|�Nb���؄�����|ܵ��1P���+*������_�N���[KW�X��/"7la'�%hh�}-`��.�С�\�x[u��.j��`��*�~�ldɖ�wp05ȭ�9��[��"�N�Nu:�e���ݕ��=�6(U;������5��.��B��N� Ƈ+��X|���ee�8�
F�����.��<kNRG^���"�|�m���6�I�>���%�l����T���k���g�d��OI�ɇKK���I��o{s@�G�]$����-������u�rӲ#���j"����_f�C�9�
$�_**���o@ɺ��+	�ꂔ�v��I�g��u��oP�2��(�;F�%lxmϖj�a�v�78��1�,�E�����d�����.D�4*H�m�Ԁ��K��s�c#��*a��)�<�Iɢ���B�,�.���͐!F����5gB�Kx��-��s�ZZ�Z4�K����R⹊��\�L�X^�7�PFA�V�''USY��VRp�՛����R�������{S;���w�[v��	8o4�8�	�8�L��g���2�{��:袌o�M�E�a�TH��d������%�5o���r�,�7��7=\O��PFC-�Jb�t��\�NC�e�`�/��>��M�HiL$]vf���p	�={�T�2�b�8�)9E�+2w��.���"��ē��>6q�C�=���59̐��7/�����Z�88���v���C.�N�:y�����VwN��9y6����2�O���_���2�q��#�R]?����ڙK��u�������-4�k,c6q�cN�Q�;���k�Bh�`�:�	Q��8n���JO#/���ɧ��G�Pr����=b�����`?������P}i!��m/m+X���vN��|����]qU����.�L�'T/˜R-�N�����p"�u��9�S:�A)�#I��9J����]�7 rE�����!ɧ�
U}F�R���"瞛S�3���!ԇ��A8���.Fh���Ј��;�9�T_��XN8��\����,��ꤖ��$�eI�J���`���؟e��[<��O��)��eh�m��e*#�\���J-�ow\6���@O0{k7�_�Z��{�
j��o)"�'Ѵ�?�#��r�( ����:��ȤW�0o{��DNQ(!|y�{~)�9PhB�C�,}Xp+��0cQ����ܱ`���X�цH�jNHSa;1�6V%��6k�\�0ޚ��0#/'L��_
O~�k�y�+��M�� r�˂��-�۔�ڼ[+��@>X��be�E1x�{����s�@�O�?��m����U�:<� ���h����24��[���I�q�;�c�ߐ��He�>�c��J�E���ꇵ}9�ǹ���e�HS�e�)'�W�`��a!����Ӣ6�`�ߵ6��!���2���'m��!����u mf%M��&|6����˛ o�r#�qrBE�!�u�� �j-����/|t��q��׎����a���$y|��BW�n����v�����;J�\�@�v�i����{������]S�R��X��K����s�Boȿ�*��p�,�hP����c7LDP$�����\���:V�-MPK�F��x��Ѓ��;��^�G���o��Ei�� '����CKXr�Z��0��p�����`"pb<�HuK��`�a:�5�fT�p�d1��wU'���U�8|
l:��;!�!��'����o�����2�_���1}���wH9�+�����fnBwA�v��VE������+Ayjv�D"�<i�4�З)��X�.�`���y&ݖ��Nz~����=܀�#r����q-[}���[=.�	���	ư����8	�~��tvH��30��m�jy�R����ك����Z����.�4����"g�Y���d���&��-��Vğ��li��$��S,� )�,^�.�eG���
q���3`�*�x�,7�c�"' ��@�k� NZ�.�<~`*��W�Z)�Li<H���܇6��MB��%�J�s������������,D�>��-��I��Ʒ������K	5o�k�+�:�I����sKo�Q�3m���z�F �����>Je��||k�����Q�E����\�E�h�Le�z�a�M��2,Ë�ɳ��: ��t��п1 P����0�œ����+���9��{�SAF^"@�t 
=���AV�� PF��ȏ���K�X���1�3Z�q���obqg�.�5,�".YU���^H���
0���O���e̹L��V�mu6�-��&�Y����f���NM�_.�?-Ks��W�\��,�����9e��$d5t�Il/lxb��3��Z�>/�<��.�����տl�ff�n��S~��}v��Gå�9fN�;�2F�'ࢌ��,_�[}J�<�)�Ex��PT��1�9��]G���H�|�9𧞳zx�?�B+Gw�ɡ#;��:�Ò�V���l�s�k��~�oN|�ҁ$��uGȋ���cdŅ���$v���B:���J�|���*���j�[,�^�fߺ��vL��=�i���1?���ඵ��>s	L��E���������=�ҍ�G��a���!��2,�7\�#��^z4�7�`�+D��6�"���� ���#��23�}��(���0L�c�/I��ga22���w�?�-�~��G��߃'����c��1�Ӽ}�f��뎙��}�o(3�[������:A�!d �#�,s�+���jy�q�������.�Y�R�PMPJM�3�j~��6��u)v��~��?��IBw���۞�9��]���7��)!��z�]I9
�WF0�g~���� �ph麱� ��l Ud�ų���D����S������e����a��-7�m8:��Ǽ�R���&Fs���Z��i3��ܠ��&�ԓ�\�g�zճƲp�v��n��E?>�Q!?1��3}�ApSg�� 7Y7j�8���Ym"��9�1�f���1(�Y�{�c���IG�]�GyI9��FN1�b+">�m�J�i�����G6\y<�w�x����|7�16f�]bҧ �?����� �sb�o9<�G�Y�m��(�Y���Gx�<��0?���~w�J$�u���۾?���� �+O�|�-��
�^ѣ3��f�M �[����3ԦN�(���������8|����_uj�Y���b�B��8�-\Q�wM��ZNԉYd�f��`���Oc��C�R3�o��9��P�34� L�NL{��1��N���˧SF�r0�jS����Z�f�Q	1J����ӤY��)f�z_�jd�q833�[�q�X�#'M�Kl�ع�/�y3Nk#:;��\&�M
���6�6?z��G�o�I;�Ƅ�ό �Ԭ����u8E����}̉��-�I������V����^h'�i�AĒ�n2�C���m�;�y��~�jn�O̒~���s��g<�s�ɢ9T)>��J5�g~��r.�r£^��\0�t�Z��E��r_w��-�2�(NPW��Ihϲ���-�,��Z����-g�
]����@]����>݉f`��D��oc�H�٭�s$2}�).�o�\_����C�����E����1�z��P�;���WO��M;0�̶
 p�e>`�*T���,R5̔8��s�XT��3����A���A��?��� �~�s;b��p�6�!��4+����V��9pG �Q3��h�:ԧ*����eD���412���?Vu/]��6r:�BW3�/�~o�` s� ĸ@�f��(�L����8�lՑ��U�1m��6[[?	ׯg81α=C[�=��瀜tڃ����rN�����o	$�]���|gX�QT��ۙ�*+g���9π��ׁ�=���g���/v2��}U	�y�|@������M��:v���?���y�����S� ֤S�����4��"���5�6�sN%��Gs�y�6��O����n���V�|9N�����7��TT�t�����7�F���%���V��������xEsV����z$ne�L0q������@�i�U��9W������^ssv.�?���H���V�9�B��h�C:n�����=5�,^7�n'���>H�>�V�U�_sd�W@���E�\Wqk�9��jh��7{������aq�g���#�e<-�x�#������;��5@�@���l_r�O������s6#�[	LΗu{oi5���W>��S�/#�P�G:C���)=P印{*c�`O�b��������+9DgC��;�HX��q�e;\�����=��a�9���\t��ZC�!l)c�_�K��^���<����V��Ay����}�\���05��F�*{�x��3���]�](���27
�_�lgvL
���,.�y�
��>R.x��5k] B���(i/y��B���7�T�J�T���E�X�D�X2z�O���
��I�5�I�7{���Żo��z1��A�sa�<A�-sH���d��!2%�}�L,X`�uż��{��q�����a����AAT��ƅ6���b���<Y�Ve�WJ)5��>G=�6��0�gl��::�J��-5�;G���f��X�e�)���|��`��r���<���O���%�W��H���,���R���	�|��MS_h��/$">�s䲰�.eFݙ�5jOd/ó]��|���Ա/>�7��h��5���k�e"�U�� �	��ѩsZ�jiF��|b zڷ`_���.+����+�*�H�]s��?��]]�,8q;��M�,#ڌP�3�8�l��x��x?��A�j��T�]�\���0���2��ގ�3���]���G�^���7���o�%>O�y��W��,O�����l��IQ��\�n�ս���t6��0����^G4R{�*gJv�[	�9�⇢��g`�����ބ�-��D�E=��%����t�����ܼ����f�F�ͮi!�^+ݽ��m3u�2{���t(�A2�7c�y%�|ߌ&r�Bu�x�8:�ù�L�D����֤���v׏q��=��"��a�8[��msW�:����\5Q�{]�_�>er V�}�)�5toSn���@�������axP�P�����Q���*QR���P?#!���3���챭����ѷ?���qQ�}s����,���Y�|A�:5����D?�Hfǀ�Mn���0md��G�������Y����٠�m�4�-O��94�n~q"���;zg!�1�'��:ccA=`��W����4\�@����5��\�=��A����çxUX���ۮiO��������,?�������Ѣ�nfw�`a��rU�}&V�fȵ����[�aGQRE�g_�쎞����4L����O֒�-%��G�Dҧ��T������@cq��z��¢C���v�)���\ԕ����t�F�zp�����C�F�Գ�Y����o?����?�Q<�p�g� $�+vwr܁R[�����QtS��X��Te�����*�ǤӃ���������mB�G�v�UQ�oD�'5���߫5r5U[��H@�+_�0��iTxv�7��<'�s����Z%��X����t}=�S79�R��(XB�e�d�@b{̮x.�\м&CF6���K�)a�QĽ)�o5�4荊j���7-	hV�dݣT����s��*�;��$���h�=�lߨ�;�e!�c�G�u�Kmm`�2�����i�yA<lb�]<i�+�W��m���.}D�{��,k�O�P�����KU�S���Fu���u�{�h��MN3��M��k�1����E�F�$��MH������id�zV6%�<�s������^���8m��OV�{��h�\�)4-NXN��=���}��������u/�\�x�Q9�#h��J�5)�!�'�!�)ˮ�3�A4Qoz�f�sL�6����oՔB�b;�Έ#�=�Û�zLw5�>?&(4�A����t������&�"�#E�"����0�+�����j ��3�$��U���)ݠ���]ž��¬Uȕ��>�}���.��?&??���KAC2DL 2��r�qkt$���7�;	���n5�F��J���V�6��:�-���K�U|L��s`c֘6n;{��Ln�\����vK�4��r=��"���=�Q�@@���^�+@����HT�aa��[����8qkl$�1����-2�u8['�ͧ����Fը8�tH;-�
[��G��v�U}#�7�"g���̣:�>��7ne�߻�ݞ�o6 �D���`v2=��MR�g
�}}r�u�T�4�Q�ܐ����dE�d�;}!�\�@�<��c��5?��Q���.ٻﱜ7����Rq<ҳٴ�ʟ6X���T�Z������I�ln�����w�r��	+��֕M."�~P��i1&�������Ӊ&j�Y{�B�\���C$��{���kq�_���UG��!�L�Qå��e��4�+��Yfژ��?<V��H�L[�cO�D��
D_o�P)��Z�C�dʭŖ�6�tRB��2܁֘E�qv��s��_lVU��ya�ȵ��I�����SI�zڕ,~yB+G�?���7A�3�}�M�(��`��1�)�$G��.K(�x���)���6�n�,4�(�o��b����I�5�m���N� ��"<�F�S�>])i�o�t�[ׂ��P';�ڛ��׫$���b���L�zcr����D��>�;ZœP7M�Y$8����`��Q�����n=�X��6���Ou�����^�?J��;���(�7w�%}��l4˯������D�ؙ��_���5�����^�?ub�H��恷��'}7�Ԓ��P��W�_��)"^V��-�1O�	d��^Myc�ʫ'��-�f���P�M�ta��'g��\���g�J�j���Dt{� M���R����E��v��� 6O���Q���y|�Z���q�i���n]W�f�X�;�k�Ş�S8c0��h�Ƙ8Jnq� �]�f���L��q((y%E��~�������P�n�hda8ŉi@���\��V���Z;s���(q�P����h�|nX2�\�F[AT��D�M�2�W�����Q��N���!������5�@�(j�u�g)�+y�6��A�ϒ�i
³I���u�ZDU&�l��$D������Y�g[�R�A���^@�|��C/G���zH
�}~�FmH�����+/�oܺE����C��w��߸z-,�M}�S#W#=�����w2���` �Yp�H�>�������U~(�4JH�T��CV�>7>��N;�v��JZ&-W���b��di��}U��׿S���*%���Z5��6�y�TKEf�R���\�Q���~�披t���
�kK5e+���8��3��Awe��=J��Ǝ���/uJ��.�����=ݲ��C �r�ny�g���<����5��vO4�wt`T6J�ǂg�܆�TZ]�N�ܯ/Cղ�ق��m��)�,�����R��r�l�u7�L�M��z�_���Ww�n�y>qS4���-�J��y�
q�g��L#���f����X��,�f��I۸k������9m�ʉ"�W�J����q�x��&4:}Y���>�ܩ���B������3>���z��������`� D#���r�l�B���f'(���C̈��֪����u�ud�ɭ�sp>4��F�S�wH�0��5:ELq�;��]������!�Ç�[ ������
�f�!/*�O:��O��w�>kԒ&Fa�/���(��o��#����������:z��<+3S�����b5_��vds"�>��]ͷ`�Ʃ���sa��d��4˥��@��y��e}z�Ґw�N���z�F��y�rx�Q%��O&�����Z�ph�B��3&��5v�Βq����__�(:
+1N���I>Z�ҀNv�����8��A��b ��Fm��N�v ����3�[�+}��,�z�Q�?++�\���^cs�r�<a�%~l�;�E��� wr5OM�� �(�a�D��B�{��@_6���`p[5�9 �tK��-9�ԚJ	(I~� [b���4fN�m>����^����9�9���]?�Di�*���a2I[G�����m,=���	�t��9����7y�k�,^ӓ�K�.���i�&q�^yxj&]E�u��+>r����7��'uR ���+�c�}�/��
���eW�?"l�c<7'�7ߊ.(ڈ���+B[��vOcP#��,��k��R�,e�(��УU�L�ۖr&��(Uk	C+~���E�{�ad-��Ks�������������e^�ioi� ��Ro���G�ѕ�,̕Z��P��n]�=�oeq�Xm��mJ��j�ՄN��v�/>νa/ΰȫ�|�ᧀ0��M�V6�6{���t�("l��q��(������M{o�l���2���>+#K!���8���d�v-�kp����실�/饸N�"5�ՖZo��N�i�J�\���!��פߐ��=�QG�K >�VHR:�@T����(�#sy��䴥��������� --b�����tV��4���_�ϱ�nC��9�9���͍�Ld!o�@&��&�<��Jl��3]��)�3띝��{9�M݂��j'7?�;�\@c�� �|)�������vk�|��%U�'�{�weU1��nI���`By�a�N>�}H�[i�F�i�cʊ�Qr�!=Lxq�Y���Q�	�6�k�>ASt��#�Vx�[�_����rM���1�#�j�D�����$}�&�^zhCH�8G���$ߙp�u��2�鱘�	8�w��5��n��K藪{��5�U���,�y�M�ϫ�ԏH�l1�%n��W3o�G���T���S@�w�9���L���^���p���\ݜ?̎�RWk�lR�v&�1�f��J����t������"7R�}����~�[_ZPx���0��q:'��N�H�ƴ�޾�0����6��=]b��oʼ��T��3LŇ�y� 27���$��B����Df��Y<,�����8���+��,j�qF�DltA@@@DzSQ��ti�.�@Bh��#M�RH�D:(�БZh��-t�'�*~�����ȳ�^�^k���k�XSˍ�8�˚���>>�4�sD�������jp�d�����~��g1���Q�E�''յQږ����1tr�	����tw�P���%['�2=��������������E�:��܃�����%֌Xk���<Op�W� M�K�O��*ś�@nx�#P�G���P�tm�^Ng�0_AJ��#m���c^�zWH0`%��@�%y$�iלP��#`&��h�,CGQ���b�'�9#:��|g����6n%�l�in���ww\&�0K�I1K>Ϡ��3D�eM�������l��_�:b/?+]Rz�^R"�mḩ̌l5���A#˯ uzX�m���C��L��0@z8䬿���J���S��M�Ge�N��G�\�T�EV� !ex���e�#��P/Jf��� J��,<v�����D棤W�?&�'VT��p�hnG�kly�d�"��ɝ��Tk����d��)cQv�	+�!������r�C(M	A�+�r���O�3Y/\Т��a����� ����8�^����ߒ|�Ȼ��sHR�����b[;b��m<NȦc<�WNɾ)���)<��&.�Ȟ����p��� z~n���=���x2J2�@���	^�Q<���١+��T�]��j�q�b�6˫�`\e\������+��}%~����=�<�pƖԑ�P3��B�?����pw���ւ����[����~t�R$g�g�զW�db�⩕�CV;uu��?aQ�d�{�eb�3�5�@@|v�d�҇�y��[%3�o#�N�����#Ȳ�;ճ�?nٚhW�� �2�#v-݉�苛��c@�A�V-^�b)>�;hm�	�U�Q�c՟�B���ik!߱��v��X߫�ͼ�ŷ�8�b=erY��,=�xV�ԣ�p��z�־<���/t/V +۠Q��?������Š���"�\�������=����c^:ۙ1&��l*1휧�	+"��W)��p�c��Z`]��`�dfis��O�q���7��ٌ��|͓6<����ՔJ�����zY��t$�m�?��Y��i���2����#-����\�^ͬ@=���
��� ̞/�5��A��۟-@�tAO{`����(m���K���gS�A՟�F	�����t����Uo��Ip���{5���	� ��,`E�oTֿ����0 F{�L	j���-���BGs'�\��Y���n�_�,�m��㇁�ř�2d�q�M��.�Z�O�jrt����R�US�� ��~��Pzɥ���.D�*�6�+�u�u�F�>��~�ɓ}k��j��Z^�rrPׅ��V7��}��J��h��k!qXd�)s.�%�(�]�늠��,�kg�ɓ�P��t�}B������2�H�*���2$�񈿜plN��\�k�#k�ZD���6:+y��+0��ТЎ^���� 3Xm��6�U�7q��dH`���D��y�徵�_�.��4��(3��:���	�dU:�����g�t�P����i�v>A��2� �(����/�z>�6n�e���!e�����pg�"��ͽ٢@d>��|���˚�L@���A�ϐY%a\�����΃*
�������V�1R���[�҆jn��e��&���i?uwq���W�ϠZ�`:Y�p����z��2���p���l�ԍ̉{�̕��ͳ�#�z�!Ry�{��tc<�:�X���w>C��x��E#��[p�#�#�|u�����~^�����t^���H��,-���څ�;	��֓�e:�h��������0&�/��m�@LY.�K����?�i<�����Aqz�lOy��U�S��l�]�ۑ��%���čg��r�3d�7��}z�NG��Ǎ���F0'p��y��ѻE2����� �]���{�з7�%���\�>�I��v��/o >%<�Taƾ�y�f�)�9��/(���-��kf*�y$_� vI ���(Y~�q-�n���&ɡ��(���jV�?�|�r�kk.x��,�<�oZ�%i�f'�@g�~}q��!�#�GK�:/�H�o�M�o�+�"K��J������C*� ��G�Ј���lkZ�'I]����;�,^�w�hse��E��9gي�G5�����4��x��u�� V�B�z(D5�44k:�Iv� ��ҒX�|��s}�������'�б��7p���ҹ���2�?H0S���x�_�t�a�i��������Ӓ�q���W���~<�$i\C��bh�ju��_H#P�a�ܖ�G1ނ���m��D�3������qW/����/��G��)���ck�*Q�&'��dG�[Iۇ%����N���k����c��g��r�����#w��o6:$�\�h�,!
���2�o�%�ɻ�w��Z�cO,7��b�g(V| i��Ts�ȋʽ4z���ѬUv�jt��'H1�Qk*O)��<�{��|֭�u��ENI�5����f�G-��շ���v�a��Ǵ�u�C�\���;vߟr�+���$��׊5�=��j�����u�@{��.����L���s���	�Ny�B>�����טYF�+�]\TR��� W���\$ae�3L.��"��4�E�#W?<ɞ�Jl4l]�hI4�˝jU7��>[H-Dڢ��;n�|w����:����#n+F��l�D����r�Į�S�؋�h',:8�K�	k����d�J �������髿G�u��T�F�>Kz��ϫ'�/��ˏ���+�;]����|M��x`)[Q[K�~䪦�E!f]
$��SN����E�)G����A��r��ړ	fA��9憉Ձ����B:���kH�ǽ@�C���
� �Zj,f��a�UO_����c|®9�v�h�c����ev�]{���׆1��;�5�u8]3�,�f��y�ێ�K.�oiLI���?����Ox���� �ol����^q��9}�-��|��p�,I����/��K�gQr_�p�1�|���>��|K�iӻ�/�Gފ�l;���Ħ]L&���Zk\'e��ݨ�~bVuGdu+���V��o�*�{�!��M}_ R���n�%!=�U��3@m�2A���e����U�י��j�XW�N�Jl�-9][��K�q�B���,�*���J�K�A���rĽ�H�9���E����I�^鿫�̋N��$LNM
Oy��W������~����oFW��Y� ��o�	�v�5K�Oڊ����Uڌ���u+�/;9v�n�)ޗDw�6���]Rx�<�?�M��}J3��#�I�yOn�_�1ę��>pف�Ұ���<�uϤ�nL>Q̈�ڟXͩ�5�^�s��qQ�M^�qY%�/{�BT]�7W�l̓�)��P��H�����7��y7����O��;t�RixB�j|��K�2V����ń�̣$�.XX��0~��٨ƛn������ﰪW�Kw(i�n�B!�����)u;��^:�n��ą�J�k(�sˉ�)����n�'�e�� ^�ǯ����ڒ�`Y�Ij�Ms�Aō�.�kĴϙz��6s�͵�������<���H�V[*P�z%��L�(�v�V���R�\c�93w�D����u���p'9V5��ۚ��FF0&���dZBgJ�9W�^��b⩄W�ho�ET�"r�QY�':�5�5���4'�S����u �3c)~� ��3�-�eq�8�g���СJ�����6O�Z�FZ|��T�o� �y���� ���#yJ XS$Ie\^Е����� {O�c��J�Ҕ��g ;;�Rӣ56�t�~�fS�+_�+Y[IpsC�k���Ý�u�c��,C%�<|~�J��7����Pu�4�u���/��	<��/��K�6����~gm���/JLw�׾nl�GD������3�#��Rw�Kn<�>���u�D��"��t��{(�*tcZ�D�qQ8~�s��\�Da�S�;*n����ݤK�L���۝њE�Gݴ_�Ƅ�^��~�ǋ�b��4Y����N2ɒ��Ρ5;��n��T
V=5h�e�����,�y��HF��}��}U���@���h�#]�oƶ���VMUEŶ�����yw���������iE�������ʏNH��q�TnM8%���>��z��f|���B�
���?|�F�׆���j#��u�wn El!q"�ϴ|
��{ո0v��{]В�A��H`����fO���{����STP�[��w�-�[�a�Y'���X����6�,�T<4{Y:����o)���>]@ �;O���ۯ`��p�}��X�w�}�Bh�D�|u]Y\;�{��R��']o}z2<���`L�,�粈j4G��^�A 	6ddR=�3�4��u�yb�`qAN���m��]�i�:�N? J9����H�F!�y#	��[��F E(��	�j[���S�����(���y9���<�4z�j{J���;W���s"�ƒ�c� �
��ɚ�}Y� �n���~η��f��k�8�s<�&����?��Ҹ�����Ilg��5nñ���Ľ����g-fW�V@H�Ϋ�/�W����ٛ{,���ZR��{������nvL�e��uwmDU������~�S@��X� �X��zRl�v��9��ݙ,��q�Y��Y�E��4%��ps �s.,�@96L�Y���=~��\���8�� �g�8!�]H�SD�%�4���|S��E�);wїz�]b��;�6H���#fꛦA�V|A6df�~1�����v�V�����C��!&���c����"oZ ��a�E\Ɨ����jS� �G�w�tekq�����m��<죾���e���ۇ�/:�7=��(�<=7�|�p��	�]�9�������'nAGL���[�3�wrތ˲��5�_ѢxD�?n>�/��d�]4@��4��v�/X���%����w�t��!�o��*gL&���a������B�G!8�8a����-�z{��(���˧r��QlJ,�����P��������Nnej0��s�����a�- �-w$�����NE��x�HKI�Q �����Yĥ �D=�N�<ٷU���1x_k�3�ë���
�u򄌹�ྞ@�|O��v����ˑOp|9s�q�O�Kq�<i�h����7y�k"R�@<̋DK���)>`�v{��Y&��#�x-�wR�?�a͋hd��ow�w��.�s2�����<�n?cb��0��b.�t�X럠��}�9���4�*���|͙��f^���/�1��C�`�ke�gwjzc>9~uu�"i�y���>�����l�G�LBȢ\���s
�ԺjKR��`�x]��IխǓt��g(�R�o�= v`�N�� ��m ��P�@�5�������7�;�FD*�V���++�(�q����@T���u�(�(��h&����Q@D�	�Gʙ.n~>2
Y��v��{�UΘ��X��Mt�cM�[Uidq�	��b�Ź�4��yo/����S:e�����z�}%l7�y�z�}�>�.;���2�:���Mʿ���wZ�d_rn���aiڅ=ܾ�qvחB�N{ۗ�y�MOϦ<���H{��C�����y7KC-��d�.w�)�|����-�^��,��������֌�����D�~���@��v�N?�Ԓ�fV����oS�uw~�_����ѡy�/���
~��}�#Ӈ4�d!�tHȓÔ�s/1��G9w�(�e�SG�u'�Mqv��>�feqc��1-|����v�J:<U�*������2��+�h��<�u"�: ����k�إ$48&��	)��\�
ٕ����͞����Q�V���{���������/�s��oC�>$�n�.}�-k��D�oJ�:��ɟ���;kJ2NGqs���V�&��r
��"���B?N����@w�ኦSt�|��aY�Xܺ�JmN}/Ͻ�S���䫙�:�R��Q�z|l1Z�+e��j�;̈~)9��?�#ETz��!TY�
�ހS�j�O �xmE{>V>uFY��n;�L�qnݶ6��]3ܗ1�|��g���4�G�|d\Z�X&�W��%%�dy�ֿx���E������|)���ғ�v)(n�X��Jf����O��M�ۧu�&�;�������w�����H�b��xBNש#ؾ������1�B��j��c;���4�9')�l�T�ň2��ӡHIz��oE(����G�N^�(d(�_��n1�T0o`�_2帰�F�Q��qQ�x<���g9%�6|�U�Ã1( �s��>�%���U|�O�g��]č%.D�Y�Cr)�ɕ�z�`�er���<�5����Msh�79`<��_�л_]�Ȝf�����OM�$���s~o��0� ���{�h�T� �RT��.��
���%^���K9�٦�K�{�{��-�P��r�C'5@3�dOt�ª.u ��%�8����Fֿ��w�|�y.�q��U���G��^T2���<�J���J\�p0\P]*��yKV�-6f\�d�6��0���X`�?�?�P�H�O���	vЈ��_��N�VH�\)�!��8o�rx�O�R�߮�|gہ�rI	�p��՝Oj�Kc������4����^��c�~>A�G_��P��\��A2��>��0P�]���T��>l���+E��Kڦe����6��;��]�'��ȬvO�f����ɹ���y~&O|�g�em(]���"� {���ʺk������*U�am;o�R�?�9���WpW	O����q��n���o�ú��x����s�����KƟ�.���P��(�j���L��^��;�����ގ���s#׺齺Jo:����؆�G1��Cߔ�VD�{��x�l�`�ȳ(��H���W9ӳ��B�1�ծ��
\}�Z������ C�������#�$#_ހ�E��l43�5�Ɛ���L�5�æ׉�U�,�޷� ֒W� j�t+������ p�G��t+�4��ȡ���2�$X��k�Ύ���1�l��ɸ<��� �Ɛb����y{�G�߼���׶*}�چ#�_��P��}���R$'f8*��+���!�R���8�<��x�����yO���l���݆O��fm.�)B��$)C����>���Ջ#���{>Jv1`�xUee��' v������!����	>����W{ޒ��ZQ�����ݻ_����ߗ��h)e��2�!�a������^�h��f�B����W���?Y�#�1&5eX��>/1~Eܚ���Cj��^v��NDke[�bz�j/{h�l2����]��nu=�C��m41�)B��TQD>-�݇w���� IM��ߴ���
H'����L�߅�5us����^G6<!Hi~����m��f5����H��2L���\�1�-�a��gnƅI�����5G7W2L*po��W��ɛ��4�����c�V}Ȳ�
o���-H��"5����R6�0&�;C7� ��{�l���w��B²[��d�$���Jڟ�Z�z��k"�����3{-�~����N[�T��qR�74#�]�;�
5��e��{sj���9^e#B�x�e�]4��*�B�V-����}N��fTx���:E��1�'+9��⌁���¼v-����v(�N��Wx���@`7�MfY��]2K�v�1���^�te���Z9CDDv��cV�n�[������@���7#[�9�2�:OU�42��{�-���c*$EY��A��y���c�^��~^>��������Y�1�2	K������1/ٲ�S����2����;떗�}�I̚�n�ѽ6 �hV��Ҿ]e��q�y��̗Q��9�(|9#�#l,,r�WK�I���;|��e��"�����j
,��| �oTba3�u��KҞ�ظ=5B;�T�� �5�>�#��j��Q�N̠�nEM�ʻ����h�)g�
��o�dV��+�(*bI��W���^� c�͏��$$�+]������ˮ�~�C�u
�F)����E6�'I�z��S�6*^Bx�bl����V���c�FW�2�!���ۙ�2�n���M��v����_�v����G��䭄�jv>]�K3��;��l)2�7���e+���
������p뇶l��w�M�{=�o�N=.iF�Ԉe;Q�v*E��*��ᓗ O�#�4�,�U��2u~�|];[lF��b��!�9~�oV��%x~ebo�Bq����6I'���&1Yp+�F�W��lc��c\r`w��| <m
"�o:Jk�X<TP6>�����s�;�W�,w�������}��������kP����ԛI]M�4��Z�O}����A�8���澥d���`2W��Ȯ�^jŀm����3[$�	�t ��v���/�6Ñ��:vɻ���{d��ҏ�^�-$t%JED"TQ�-�g?8�9��"{t@��Mh��,�ڮ�ݚ�6R����5�����9�TZ4�\���p�e�2����N2�w�<�4�o��7�;�b�.��*σ�c�	�����~���ÀC����l�Ҋ��#�2�A�l��X���d���J%��k�痏�>�A��={��ۛ+:Q0�����>[	\iY�2�5g(���cS�� R�0�x1��t�-��栕%��	�	�{�BJ�`F��y��b�����|�^Nɻ�a���!���i�7��7�$#��K�����MQ]{�;�^�H�G�)��D�������	�����C^��	�p�{��N .�5i��#"v�Yt�
k���L����.v�U���w��{��Fj��� ��(6��M0�X�W#��hWg��Q�H3.�5x�Z��W�V�ri��/�<t��/<���>�ɚ	��0ٳ�7����BE�L�I�N(�ǘV���HꞳ�R�ܤ�z\iD�]"�W�1mPdn-�W��m��?�NF%p^9&�mX����R�I�t� ��:�hJ�VԘ�'ܩ�Kg"��Z}xv�ɴ�eC��;u ��,�y�s��"׵>�b�s} �9�������`|臯��3�]D��#��rȸ���T���}�hEfs��4�ǖ���{�j��kB�L�Y4�'�?\?�X��UW�a/�7�ks��2T�ݯw�ӂ�m��cK���8��$�ܝ��O�$
?��|�j~�#�/h^�����2 �@�*����_����YMw�׍��K8{*p��\�����`�����@��������c����^��E�^��b'^"�S!�0(9�Us1���� ��I�krk��z���-^��k�᛽�1�ad*���:\���� �q�ܹ����}G�}�+�/�i������Odk1�	4w�����Wi"X|�ݵj�x�yh�F�|ߨW�|fh#
_��_R�gd��MnaVhY'����#f��J��}4�x��TD�&�^۬��@)y�Zs���t�xw�x��n�#M�����:�d��4>�����]�x�>�7֒��)��J�B���}o�h�V�X!k+�/���CT끡��K֡�K-;���nx;��1����|˽�c�ɜ�P���X��JY���J�&HJ"G����jоu������W=�����h�]d�{���֤Ny=���F������2�X��&��]I�t��8U�J/�^fm};���(lzS�E)Tܺ�8��U��DO�H�*�c�{��l�PF�C���Q�I�MY�s�lV�%�L E��(ĕ>�f�6�8�jｊ��A�������̆H������bH��p�˓pM�̧�X�¶�s��|%�|�Ȝusc��@]a�#���w�RE�嶽i�|�1e��eA���d��NrĄb4D�$�8��Yl4�qd��^n��0���Z�j4փr���so����^����^�	���}L�>�+�,&��Z#ӑ�o�/g�!J:GP2�V��C��l�ƕMYs/_�%'�X%��EV �Hd|���UR8�	�=}�\!�!y�M��أ��n�N��/nƧ���.�(ź�r�h�]L�xSSP�h]�(f *2聽���@�p;�w���ķ�&�Z�C�m^�\��D��Ț��/��J����OOrw-P���e�!���M�Y��"sr�>";ԥ:�ϐ_'fG��N�[�rY����\���e^*�����i�nn*&C�.E֬U��ͫ�Vt^���Y�:Vbߍ��J�(+�[�!�?C��뺏�H�E4�eW;ʖsŅ�7��v�,^}w.E�����W��h.�u���5��Vr����}Q�A���212���̙�M#s�&�q���d�:��f�W��S�l���`�ė��sk��#|��麋�1'MT(xش�_���A�廲�F�f����>O�^�W_����o������N�Ds(Ją�">Ď�[tT��e���'���u/	��OӐ��h�^�,���n_��lޫ}���4��e}ޝ��V�$&z�c�S�K�-6��bv!l��p:�^�ǹ�2�~�j|��^M�ػ��}��D�8���v]�\�E謊a&�1l�ˬ��4��~�?�k��|���Y#"wi�I���/˖� 2���Gѕe�R?�Yx�D��K��2��(%EsB����f��]�ǫ�"_��R�����:7we)r��ً��vB���׮Wc ��h�[v;��e��oS%�N���R�Aη����8:��r���j�m���=���,N	��ފ<��47
�hʼ>��"����T��&�p�,�f��y������De��\gu�K/YIn��׽_�E�� @w$O�^QW���2�@��1F3�􃓟fd�ܹ�P�
�hٟ��v�������+%�Q΢���d�;�x-��t�w�TrE�[A���N���F��E�`{_ҹ�_&���$(�n�n~�XL܄xȍ���w�M�n-}Ѫ^؉��[��U�=�����_���J�l @}���b#� s��k�7�����x��Ce�w껇˦v=wH������E�cϪ;���������]owP�W�,5W��|t��i��#8iT.s9�}�{x�u�&�v���l���}��7��GPV�zc������p$�5��[����vF���[ʆ�gj2u���U���-.,I��x�����c��|��br!�ËoY!5v�c��p�w6h��r�Z���49K���:���p�w Svy��-���2��� �{���"|�zRa��*����G��&rl���S����d4��.�>dd�H�"��)�C��H_	�l)]���ś�1%�VHl�7��&��j�|��k�^��>O����ɇ#�.�Q�;d�H���[]������XvL���xjc�H2���K��.K���*���Eσ���=����U���d���v3f�I�}V^���׹"�,�y���a��o�0����u��[��L��%qG���wj_y'� mc�޿DrX���m���,��2��Nn@�	Q�p�R�_E92*���.{53j"�ۓ���d�lʗ
^Vz<��R�<3�/����!�]���:��ľ!b��D)k��P��nw5�4,�#d���
�����g.YU=���vu:��0�	u J���� me�:�ZI���+a	�F���\���ߵf�����Y/��f�5��D��Z�'��ӥ��o�DJ����^�YeM�攗%>{��<fN�'gTV��1\El}�$i626��^uԪ(힔�$XDNn�#}����I���
�_f�ɽ��b�C�A�&�h��[�;F�r�����f�t��B�wj�M����	(�M�!�dYT��dZ$=!���ӻ�C65T���֥�0���}���lb�|�_��;K�r�Q땦�s��� ��o�1`�j����ڌ��2|�ܞb��K$����aG��ꊳYn��R_�)zm1��b�Z�����d*D���t�>�������Ϻɍ����#IN5G����2��5".5�0�./b����D%�vX�N(76���U�7-��뺲Gϭ��y���{$I�:��������V�ƍzF�9vǳ����9c� Z���NYrb)��'�¶%����w��/c�ݠ���G�%CM%o N�;"���GH�[C���A<Z܌��|M�����2����S���Tr�������7��sQIѐ��\=K%W��Z����K߰�@]+6�o.2�']h�%9w]ZJ��4���&6�X�%ڧ�V�/������2��@�]VF���k3+������˨�PA�ʛ\"�U��
�]��nfE�y�i�uC��l��뤫��]�����e7�&��r��[痲��>�y���D�K���NX_�&Ķ���v&�׆J�s�hxw��]\CI{�|gq�� �������V��i�b�_�bܪ�_�;A���4���J�r~�>��mW���c;.�.N����c��0���+�Q�z�_��U�P@>�j'� �ti4�r���e�p�R$��=���m��'��8"�w(���|�}����ʣ��G�o%��7�$4?�?���S��U�iV���MQq�'24��y�s:[æ�\��d�1�c-�T^~�N�k�	 "��g���}F���~ۅF�'�sױ��s$d�sy����̗��٢7���� �k����6�.j�ܓ+�H�)C�	D;x��4���p��"[�x��W�5�;���Q��T�;h;�~R놕�&$%�=+�23���N��]���\��.F�胚VĉD��v�A2����%5��ؚ�'� \��v�\�����F���S���<l����Hݍ_��d")@�Mę��`�T���Oڸ����{++�i���NFW�5��r��
�*�&$\Ue��k8w��%��)cW>@d<r��I�l%}��M��Z�R�8�a��
q)B�@�r�:I�����J}s|�`F����EXa��[�Ee	�'2<�.)�5������	V=�<��3�W�
	!o�>I�`�J皋tm��cl1�1v��Rc_�4�)\+4�Uhz)
��%��[���(�ATd���MF��I`l݊A���*>���d�b����Ӏ��`��(�.����P��U9���@m��)˟�|���S�V����@��{a�K���e XC���Y�x�ڨ���.���{��L?���3�z.d�)`� g����ZI�P���G��`� �-k��K9��WJ!&��L��yb,�ᅬW#2�^�:�J��LW��1*8&0GÒ�ͦS"A��f�=x�WD��*==[���{/��T(Q���wˏ�����K��ԡ���@�����:U��r?�����@�J�<�0��h{gnd��j삒���u���������xۉ�v��ɭ������O�1N�tC*����Q��������y>DP8IU�����pO"�@ї4�g�Vy{Z���8�'A��D@�Ce�^�S�	���}ή�H$t��-�GE����?���W�'/��Kbm�╩+7?hx�hU%N�V�)���#`���:�;^}��B��ϧ:�+���[ؘ��C��KXb5dNMvS'>�2������q����J�����{F'7���QK{�M.��Y��1"�>�e��s�h�\�����_�A��ӧ�kd���Y*,�Ҧ�ɌN��_V�j��?��>��y��2o'*�41>o�_\�@<c�wU����ڔ�߾/R����ԕ�l7	`(��	͗,����%Ēu�ߺ����|�t�+Z���d؄J&���ΫIl���*f�}`�+���̬xç��<.��L�(�\�����F�F/���w��˄��2�a���fe�|�)����Sj7�y\���`e���Y@�N�����/iΚ�2��6�$�bΊ�*2�C7L���y@7��,��p۰� ��@P;��I�o	ղ;a*�` �..��<�0&|�e�-Fk�$z����R\�a.��U�?&Ӡ]���*�����G�c��U�N7� �/�:6R"
T匈Y�^����W����>�N��*�I{�ʇ���в��� y�"k'%k�8�R�����6,�MR�5�g��i	��j	��7NU�<�Y �����5�U�Z��=�ֹ��/A�`ݾ=)�&O�ơ'����u@��0���SA��<$��K���8���� ��1��ML�_��#+j}jz(c�"�@�+��ǯ���%)��k�PA���7�S��[1��t=�E�:P�_~��T���:3�QjIŌ��D02�)�Q#�3j��ٚ¥��|���A�E:�9���N*;=���>$������ �u!��*�?&��h��M�dA��st�=QpKX��h�7@K���M��`��,���x�ύ\J�j��J��Q	 g���y/�r�n1à4G ��4(�J�!�:F*�$�^�g��cVė�eۛ-?e�J����\	�<����������+��1�JIe�j�σ~�rIn�$��K�J�PKv�Aq��VD�c��u"����W�1�G�����5!�nWx֖6#F~410A J3�7x�R&�HFG4�(��b���w��}��[̈�f�t)��g��(G��s$y�Dw�� Ee���(;�QB6C��VL�~�[�رf	\���Ɂ��b �H��8��o�"����&�ߤ���*72~)����Ç
�Hb��z�1�ʡ�b&�wJ�S"0�?�V��i����XM����\aN�+���+w�V��J�݃��8#_�͊��V��_��	b�/:��bB�6�s�1�<c(��O�!p�HPm1�w��oZ���"7i..�م���}z��ݣ{�����i\�c�"��|�=vhj:�z���al��¼#���yF^��o��|;��1�h��'��=��Z�'���|��ۄ�XFJ�+g,��@�P������PX�+��T���b��mݖe�m�w�F���jWÂRZ����W�"���SϞ��/��w��ߜĳ����#-,�������l��������_Ϸw���|�_��O��� �_N����K���_�}�9����?���} A����Ƶ.Ϭu�)氺+���z�ؽ�\���\�����K��C������T��n�ogg�́��[���hRy�m�$O��A�Z:��W�_�FRfT���"�c�'0� ��G
���(e뱉���7�G;�%y.|@��w{A݋S��T�["ؐ�گY��h�:,��:�H3��OىB�?�,��0���>��˝5����?�� ��r̀z�62�a�%=U;�W��
HL\i@u モ��52������)��������Z�/�ٱ��̋�b��5�+-6G�
5�����mUv�iU�j���������ӷ~X�y � �8���+̮�R��6��buu�#�w'2�����,Q�_u+2Kʹ)�������e���-���mDҥU�2y�Ld�0!���V	Q��c���A2Q�N��֠�6X5]�Jx�M���3i� �{��F����}v�aoq�BVSp����BHe��`r�����	/��ێoJ��U: ��;:R�u��������u�eyx�a�0�+R�T'z��S��ɧ@����9>`>��(_Q��a��Q>/vſ�N;�R�7cT�^�����1�s�)\�� Ȥ]��W�t7w���@�h��B��q�VG���Q����ny@-�g�����)Z�U������	7¶b�j����7�W5ͩȠ�����������P&.��=��V�M�]��Udh�y&N���w�?N6
�� ��.Cm�H���� ����f��3�I:8��������T�)���.pN};_�#�'�hM�Y�&��[;��潌����P��4]W2�D�:�R�������I���X��Oo�(J���y�륂>��K�����!vI�jyfgק�m�g�/�N[��� *\�/��ч��nY��� ��*�v�*��D�%�=E�^l�x�qB�p�%KL%��_|VW���(9Ww��:�G�РO��g��3�T�'���3�RHj����'�\�
�nZQ�N��]R;C��/��Q�+|/i�q�|Iw
ņA���������.vVsrp���X *S^V���������X��
�8O}OL�=��]M	s�D	��M���C�#c�뻀z�L�!�m?��9�)�n�{���ي���0d���^��m�����M�jxB�y,�nH:6VJ���]r��&»��k^���6Q���b �O����Q�\�sq\��P��Y����Z-B��v��P�d/���V..���fwJ���Q��G��ռ�X�(�_�#iQ׶e����7E���k$~���!$f��h�d�x��>���F:� �l7	�Y�0�6��Y771�0\�Lmq��������7��i^���:�슢+�x��s>f2@�z���r���3�*Nl���t]�VǶJO3WQ�(�7^�Y.b#C��^�ȕ�52��ɒ`�M�W�4^?AU�iw>�(\��q�ҡ=HjZp5�|Ѿw��2����w5�h��\��|�p�ms�f ȝ�D$�l�D�������)H��CpW���~\i�9ŗm]Į�5�����a�N�#�ty��?����v�h��=�d�����+Л
|%����~��~m���\��W��N��O���Α|}H�����
��f�z������Q�Φ��GTn� �� �J ��Oz(��@I-NLp:&I�:LB ��H��E�7M���IL�����W�3YG�~���#~�f�~�^�,��}�c A�����}���E�$6�'�D4��1x5m�726iu=�}s��DA	h����C1c��ws^/g�:��@��W<�����G�n��鏔Ñ����A��\�oR�*� J[K�v8d��K]��V���+٦~OkgLd�ifXh:��]W�D��bOK���P���a���=M��cf<�\���L�>�����
0�?b�ii���a�WBs{6I��/G�z���)hE��p�&�P����VE�}{ۅH�ײF1�dɾ�������Zv�Q�mP�gƾ3!�����|��?�t'����k���u߯{7t��@�smT��s�Ǿ�7ý��z��Q�xz�7C�C�Ǚ�*�9��j���Ů�t�����k��������XIK���쫍�"���*�\۞-s]����N+��#E��}R�}��^!�4A��~��2�	��K��"��MZ����gFRN�o�j}2��&_?�Bja���E5�G6�驶�Ȃ(� ,b�gB�FA��/돓Hn��`�넷p�-~�O�$�&���K4��#�K�B��2r���LЀ����?I�\�V�#ɵFw0�lS}'P=�.#�����p;��Ј0�"��h�����b��3�)�Y#�Tw~�Q#�� �x�}��-��"gF�
����{�^�Iq]��(Vi���O���4�b\d3I�h�/���ۓ��O�;�# O#珄�V�o�.е����J;F+�3AKE���u0B9��,��URRY�A��/��t[q�a,p9�H��啕�U7s>�<S�����G�����4�}j}���$�a^�ȏ��4+O�Vt-V��*�x�',�%	����J�hNr�5����\pnL����5G1�3x�'�Pl�O'.���-�ϜG� ����wR��PR����5'Sӝ]1�܇'.ԏ�i�XR8ACM(#�H�)���Ǉ�	���*�(����?qW̟z�<m0�"�i������p?|X'�;�3�[�'%ʝ�Ӻ�}�s��b��H?�ւ�E�ԙϪ	[��0M�nH�O �h棒�ְn,< 'R�vC��d��q�J���	���-��c��vK�o>�@�{����VL��L]����z�����ia�<���/�J�c)8�=��1"�ѫ��c��1�F�߭�}�[�������p-�6�������!�H�i�W�am����h�����yJ��E��do��í����V���+1]��=����]E���'��um�;κ���ɱ!pK���U��0�z΀�X�\��PՔ�T���i4�7�ۗ��2ϥ�Ҝ�����p$�35�@��,��e���r�Y�Q��Ћ4�a�a�5����0��LU՚ͷJO\��L��3e�%�^�>�׀���;p�@�"�H�����Ko�l��	H!mjE����v���DT�c:|T�*4���I[/���g���`.@�?��MHmX��x8Q�6�9�hk�"�=�����e3dW�0.��|/Y��w^�PѣzCI.ح��짐!x!n�ЏV43Ӫ���1N2nw��۳�]�7�)��G�35.L-��'FN�("��s���M�-��V����5#뫜��-ǲ�;�u�7�a�5Bj.�#��R�cbzn9&q�Ep��}(��D�`�nw�6���e�1� n��������L�?��T�Q�ԯus���昖��4��đYE؟5�b�����6ұ����.�ẾA8�Uᐚp$��n��H�ظ���O������YR�b���s�dDƻ6�(/~
n^�)���RAp����U���Sdd#O���� �e�:s�$��c�f���U�j�Q1�����F�&���vզ�|���D�3���u#��vzNQ�-�ٍu��=��6���7Z��c-��dk�)���f�?���b�Q�&[���-١� � H�7�֒��(����u�s�@�g�k�wĎ�M��~9�暴z�76���&ǚ�襆�);���
>,�����s-ĮdF� ��I�U����b>W�М=���J�c��m�XZ�_��M�J�ʩ��M��;�"��3�m�OT)��E�K����?�wYJj6!����I���a�Q��G�
ԈteW����0��W�WT�5�������A��E�"�*1��T�T���A0������t����xݒ�ӞՄ�3Xa;�8H[��nZW�؈;d��D��:6w�;��ݳ)�ӛ�&�+�P��1�a-}l�drӆ߹X�2��1�"��彡���k�w�a����H�;N�H�J9�t�����T���!yF	�)��Ԧ�Nx���zm�g3�6��o��Lu�(����m0��7~�DL�l�P9$p</�۩��Y���l:0e���8��R+��t2r�q1�A��`�������k���\��f���v�;S���
�2���@��eR��-�4J��KCE�G�W�r�8�V)}����p�lCs�h��>����F�*��	luh'�x�`'�W�v!y��۷���L�U�@`�d�����*B�i6��O V�b<��F�?�-�>M�눌�9�b�	�2�,�tD�E.�Q�z�f��c]�{kkt���[�=.܄��8�o��������k����np�_�s�N�I���o�]i!��|�H΍&�H}�J�3&�s�� �ܟVa��#O��U�3�#=)������6w�+b�"�!C�բz�R��:���)z�����k޼\�l�M��ֿ_��eN���&|���l���?�"O��EeL�&mb��!G3˾�G���:'r�������r���y%�
�uw)���+/����b�ޚ�`���ղ����s��b��jD���je=�»��"1�����	+m�.���yQߨ��\�t0x6.]�����/����
�μL�t�s0��S��Ö%+EԜ(�?����ձ�k:�;��v`��mg�x.���������"2�!���'��0�~��g�!e{� �l����m\Fqs���X�>Y/+0��t�ct<���� ���N���[����
��3E^�]]9KmW��a���N�r[�5!M�O���z�Tbnkұ�N������[6�=�NFf�U�{J�v���"��Et��z�рl�[õN�Y���U���N̚���C��q�k6��<�}��2�=f�.�۲0?eL�]�@��i܇5*ح�&?����Q��6�tWLd�V��Z��z���>��"����6��E��:��bV)�D��h$;Q��\$�Q%ρ���I�j��Ww��M�y�%rwV�W����F�x4��k�,�M�t������=
��l�����?�~�>�8\Z�O?��#H���ݠ���@�K`c�[t�
���4-�ǎ���KWK��
�uA�¶��]��¯9z�y䐗Q�>EESo�70%�8X�T�[6١
8bG�r������ig{�����>K#���3v��)D5�c� )R!��յ*��Y��KJ��{G=T�V{�9� ֫Jd���u�̧�+-��;�N�p:Ƴ�5���/�{��/h�ↅqCV��X{l�k�"@�"����ƱEb�UU ��\���-H�cq��2��\���*C���>���F2DP<�,w㏕5ew�qc���T��j��f� ��mG����Wa�1P�Dİe�2��h-t�
D?醉�GL��]J���~��ҶC���>�H�[��G5h���8t�|q��o�m��tu�%T��f�f՟j��PHzٟ���mZ����h�^���O%t��\M�6�zGD9�{2�����ɧ�_o����^�~��"-�: N��?(��4���$��Z���u�6 �A�bxW�r�P��<$�b,W��A x�aG�V�`�������Ůڏkq����(0�v�E̍�н�p��e]��ďGV������\<X"�V|�! ���}���
d�ս-�Ñ�� �[�Q�`
��nbU!B��	IͿɓr)�V�5�2l	��?ަq��|>���zb��������p�Q;���5#�Y��ǹW�������Î���3ck��>��
z��ހ'k�S�j�yy�znk���M����lu�)P�&S^ZJ���[*>~2>/�QaRՒx�yC��o��h��^����`�[Y�XU��ts������!�hL�l	����@%)M��˯J��h^���w!���6��J��'�ax\P+��@wk�\[�=Y�?~�%*�|�̞�Ș0��2*�۪x���Y�N2a���Y�d#�#�~*	�>�6N�}f�o�@��9���k�M@�k�Yάel������k��4���U�]�M��3�\���ǂV9���̑�zSZkl
qfo�jU�e���,�/�B?$
�߸��C_v��KD���D��S���(�ù@mߝS}-�ma ���ho	DZ���>���0�Ր���3 z�1����d"�~�/�ڊ}�Wc�"CPڨ]��>��q=���Y���nA��yl!ߚ�k���}O�ɢ�c� ��v^Lٳ�7�e��ʾ��k���I��T}����je���P�P=�J��w@᷋�5Fpj��گZ֖Z�����q��Nn�jR��(R3K����8N��"�ntD-,Qb��6�ʷ�8�X�^�:��!-�';�����0�)�n2I���|�@EwN�!�co�ڝ�T,���mTW}B�� |�&Y/�+�z�֤�T���Rlwg�̶��W)Z;Y�nT�͌�;�!8�9��Y=�='��%'�qI^�X�So�k��Պ�FB��K�o���%����f�r݋��D��̼�����	d��
����R%_z
)�{�$9���{K�)�ɹ�8�����e�L �k%�������`����S/�өZ����uH��Knbc�"�7������t���ѐ��Nun���g�˽�Ah���^�by���5���19���`ߚ����Y�DD�Jb&k�U�B���8~�Vh��2d8OZ[�����?<a���x���:s�R�D��'�uN#�k	����?����b]N�­|R��������{��m��d�^C�05MOW�iI4�a)OC�\���:����w�Y�8a���u����}S�?�|X�H�(I4�}���'4��re��]���pV�ԣwԃPp�a�B���CUl�w\�������F&anT�]��4(AU�Ȣط��A�(N��lrZ�٬�.5�FD��S��f��2`끱P�oŝ�m�}+xi3͞_3k�2��.�>Y���Kŕ:�~�W���3	���a�ԧ�
�*k�r���WR���,\'{}�ϗpϴ����/j�^v��?|׫5A>n�KU�B���o,tj/��;���=
oV9�mޓ\����kt-S���P�k���s�Cg\9��Q�j�nl	-�춲BI�����W!�k�-�����Yp[�Q8���xU/�����͞
�l"��ݮL�D��,�X%��#���B�����g<��g�ጝV���M�)Tcn��Xy�^�-*X���dծ��]��^ط��� t`O���k)�5��B�5��M����ɵ�����7���bT��S���� `��J0]�P�P0�����P��/u��OOVu.�{��j��r��,F���\��6!!*��܎N�����$�{\��ب��<�I߿���'���|�kѯ"����q��:.����=�o=�]FF�nR��e`1,�y�s> �.��sb?l�tn5TP�[�^�䉃W��S:�����J�+4�o���{�&Y;���  ��k��s{��M�����_�y=�t��*�Q�>8w�w�QI��\ց(��@��y�R�z�MJ3���?��%)k�^^�U�$�i���l�A�	�r�� e���nC��|qX|&y�C=̅q|��3	�Km�E2�B��5W������I�͡@6�f�B��SX��}�QT�s�#��v±�¡�q���a�	�.�%]J�u�>�ì@m�_ÿ&+&Bͱ���'��[���
�Z�Z9�)����
7�*r�׼TŶP֠�7�*���I#ب%:����pm��ހJ�}N���U�.��u�^;�o��K�,~-��F��~�S��QgqN7\M΅g0g��������K�F�ل��%=[GA�b��_��15�R���/	���ڗ�"P�1�����@ �ș���%L��M�Sy��br<#5U��7E<^�n}ۀ�(�[#g�:�J_u#�p%xj:�"��.�"3��UL�B@׊Ӻ8U���tk>����nb/�5��|zKF�x;9�T���r�H!l,������e��4�/����o3�@0HK�CK���.X?]5`���l&��BB��(���������9٭\��,ӭb�_���%|ZA�I�ĶrR͖7s��Eҁ7`����^F3�ŏ�:�{4?��L"����L��Ǵe�|l;LB!"�"�>,�w� 2F�l��I�3�B�E�7P��n�7-v��!����];����p� ��pesG"�qv��)Q�����h�U
�!F΃M'�Z���)�Y�{!���C�>�����W�qh���Fڀ���=�[*�D����o�Z�`���c>�ȱ(g�܁_]�8��9r:�XU�zw�d�3�ݢ��6��~dDP!qش� D�q�K���#q��������^��-v�8B �6kPt�xT��T����N�
�7][�(�g�U/<h�5Ƭ��;�׬"�G�� �=�M��������I�iO���u�]��>����"���#M�Ix�|6�v��@A$����
y]Ie���^��I�C�j�˭ŏ���"Z{�ް'��һvΓwn��ka<�t���t�=�?��m���7h%�B��D��3R�Z!#v�nS���U:}X����y�{5>K!�U�)�����yYI˳,Q<2:|�	��0����w8Υ�/��.b����Y 3}�A���C�`����t�����S��W~�����;��_��r�87�#(rFxj��ĺqE3և�B�wʘm0������O:��:ǖ����z2O)E��N�� ��r?�;����n�fT��l*{�w�$�*�GSV=֦/d~t�A�E��T�q U���Q��Wϒ������>L��f�b:���(���y��g^����'���T���i����oN96�
OPR��
���b�>E��>z0�g�����S�|(B��տT�?3��s_���>��Y���O��?��900��[Leש���� �����#X�J����Ϊ�4��1�5�q����բ�����}z@v��u����@M����KC�=�����Y��J����`��It��)�sCzNvQ�*2}�scttT�>M��p��j뚤�TU�ߕ�F����o
/���V�N�4'������ȵ����U�P�;���'x�E�OO���IX/�}d�-q.�hBB����|���-t+2�ĭ�i.�=�L�!�# ��Q-�<�ޏ��(q�0(�γ�th��*�ʫ�ST崚�6���M�Hb��'�'��q�g!:�y�8+�g,: +`&�r�Y�d'f2�O�Sf�"ѳyZ��� t��@�'��d����RQlv�S����-���7-�++Q*S(�?��n��v�	��Ýo��*$(֯��?Z�Փ�5KZh�o���k�@	��i���~���6g_��3�8�}����×��f��8�a�,b[�'m]<�M�w����a-�%`z���0,\��;6���n�梻��YS}
{�t���NAי_}Ē�j������B�^�}&�b)�G4}V}W�6(� l1c/��{����X�מHP:��M�A}�����{��@RX&��B�~2�-�Ǥ쐒f�y��Q(DZ���o�z��5K�)^��\_�uߤ�sA��v��#�| R���w%XD� d������D�:s��?=��=��N��/w��O�39�9�+�l`v���p��1e[��h��"��@#��Z�ow/*�G� �^�0KKE���w��ޮ�ٿ���yO��V�Ǌ����/Ҍ�L*:7��{�O�8�Z�nR�������.Vb�o�pm�UU�b�sd*܂�ސk�/i�2��e
}&���I���y�u�zY�VB��������f-�6V��Hq�!��X�����p�N�Ƚ��cP��+�0��&E:��(�~��ƍ�Z�E6x,o��{�H�cI}^�Lx�̿��"��,���la6���"�c��㝃ݞb�i�!(x� �N�69w��a��!�z����8w�k�dj�D�걗Ì�-�h��?R11EeWX(�5n�^;���sfR 0��ؘ".N�Ȉ\���[�u��@���xv��'�[��&�u�IK0b  <���X�蚘�u8�{�,�:s�0v����v^�a�
��h�4�}� �,�Y���"Z�"Z�7��Ӹ��ru<?��uX+��_�m���ԟ{�
׍ c#{�ގ���z����:`��+���*D5EwKqXQ9���\�Q�pWr�Y{Όg���F#�����|����9y�j�X���D3m�1���";�U�J0ݸ���*G���&,���x'y��V�`����_���S�q��e���F��Z����m��:���#�q�C�F���}Z_f���:��B��xw��)c�'��%��+!�<:%��񹡊�lW�4Q��U�k+u�Pמ�z�X.[�j{�vv��"�&-\��]q�`���]w9;�^�?���h�]�W���oc�kV���}���T]-"�dQ��8y�$+�1�/S�g�����S`�je�<d���G������QGu�Ƃ\~9�}r��"����PW�1wVE]��*���� ���x�1����S}�+�l�wC!c�p���s%�`����JY}�*����D4r|�a}4]�X����!��}�)���ȸ�<''��5�u��m-@��!%γ*�B$�Y�a��nH9э��p�Ϗ��gf.�����@넅�Zj��Y��D��t����b��J�̽:�����s�㯛Πq��"�q_����$Y+=w�~�Ϩ@r��{�U=�����PO����K��U�����i,�@��86�c��hMW�y�-O��J��d�L+��%�_ސ�n�x>�mjJqǘ/�7��ݮ؏j*Ї��{�'{;X�5���q�m�K놸I���ߺ�2��5<���_�L�k>m�,�m��j��	|2Ρ����\�s�^J�L��0*{�S�ޝ������0����Iá�s��>g�e�����c+������$�[�H��p�h�P8Uh|��M޿�/_�?@��_"�� ����~�ڵ��u���4>��X��)�7��2���Y
>L�u@�^���|ƹis0��81�a�;xM�g���D��oV�@�Z��O�k�dE��Z����%���?�d������0sDG�^]�t�͐h����fɵ� É�A0J��ri{������'����K2��lې��T�=(e� ��o6�Us��[��j\�� �:!Z��T�2���=%�"�ٯ��/L7A Ђ���|���nq�lѐj�v@��Z���Za(��s�RZ�gޤ�R}�A=�M�^�<cd�-��Y�\�7��{{�
;<���������u} ���Kz]7Hl��-U��z1h������&1w�5�*t^R�R��;8�6���8O]$�ʖ���R,�B����э�o��ص�L٫V����o�o����H�V
;�B�D���V��B�#�r�=;��G�C�ٝ���	���L�{7���b3�2����Y~�?ud�H[�Pk��oU����������npU㪔���O�_������Z�\_�Hy/�m�'�S���w[�~��*NMd���f�'}�;`=��i�O��D���3; ��]�>��@�{.br������Dް�*�:��%~C�U�a�U�'h����&}���X0K�b���	/C�a�Z�ԑ����!�B�K����6Y�n�5�7�h��J{k�D��p0e�?���vYA�%���ӎs����+J�4�"�/4��@�2*:��#�6=���I�WI`�}��g3x!�V���Pb(��?��8����42+߃�`MR�� �kNw�,݄��ZHzoÒ��VGy?�ey�7(�=�.r���W�OIe���J㧐�+��{ m�w�v�n��Q�V
�S��*ٖ������^3(���(](�]�;�������3��N\EU)���gW�����g��=DV{*���d����zI�e�6���,�4��e Tֹ��qn���G�˛��*��*�|ͻ�3y�4*;�tq��Z�.�-�Ѝ�r1�z_3��R#bow�e8;�~b�H{}"���zx�}frn��d�9��sϬ��Z�(Vd�B��(��a��*7���El�5��k���#��M�Z�	�G<�kf{&q"��7O�(�WO_���FZr.2�?�$+����yM$5R|�Φ.�:�TP�[Ũ/�F���
��~v�I���
� � &�+_n���:�2�1Z<�*�h�J��c>Dd�~9�~�Hge):޻Ĉ1(,۬�<u�P�D򼏥|��ִ�K���E9I9_�o]���-���c^�<����L%��l}ڀ�\*�;X��<3D�#t�]^C��6E� ݤ�b�ö^P�PE?�D��GZ�b\�^����9��7P�暨K�9������,���.��β��9���̓�z�]�ݽ�m��Uf�Y��4��̞��z�|d��/a���=pgяiKڱ���Iz4��@fJ;cV}�(C�3��P*Wun+��1�xL�L����2.��y�(?��g�HK�~�Y
Fo��� ����J���>2`���_����߀�S�}�J���B�7��Ѓ%�Ui���:L�A͉���=�ߌaW6�8�E�3���&mV_(���
��}bL�`sw��.ם��89G��k��D� ��ð�����;d�9�lo_����l�b6�s��x}�J欠�������� �j��'�Ѩ�������o_6�PA�0�+Ч�!æ��=D�w���'S�;���䜐z��R��	� ��Xt���7�U�L�ޔZP�XS�x�:�D��Io9�뮼��
�^���3Vzi��Mb��@b�e��2�;�Kׂ<�۾^�6wtn=6~!�E�m���Rx��`�l�v��<�@������c�xh����6 �V��8��c ~E����;��7<�]`�;Ys:�_��+.-Rr�������S���#r��R�W��4�����3	MH��=[;}��4#i�,Y _:��7��;�;�Z�U_�^'1�G%��?�Cк�>|�e�Ξ=�n�=��	ZuR!�7�>��h��ϊ� �_��QSW"2��߫E�Ջ������h��X�	ԙ�*@}�
��ߣ���I�&�=W"��s�����VD�B���xҪ]d�5�n�n�<-90�T���$�E�g�@�L6zUۡ���.nrw�jd?���'�~�<����r��Z�n��)i����q��}7�=vˉ�� ����2��(�QK&��t���G��̈́n_G���i ��"�f-!s�o"z�(�f��*�ؗ�L����e����w�h�<{nwݬa��R�B����B�P��zIc�:.�"�U�N�{�j1�:��s��g���)(۩�ȋ}^�+��0�h�e�!�Ȉ]���;�qeJ0t��k g���>"F�1�n8�s>@X-�3�*��?F�^�S���g|y�@�JjT����WZ�4�d ����'�tgy�B�P�F�3�&�����O�|�]|b�
{�^��] ���
��^I?>a�!S+(��ߗ�W�����Ql�:U�1����A{l��/ǿ{,�/ȅ��8s2�6���8<O��&��������Un�W��:%�G���NB	�L�E�j�4`�Yd�C}Rrs�J;��mBB���*еa����_� uE�9Bʭ�m;�Ĩ�*v��%�{���y����q�Y��D~f����}���!O"�O2#@�Ű�7]���P��Lg�:�Ӟ.����-翹O�5�����P��C�����]S5��.O������i<R��'�v���RuD~�2@�h&��+����[6۸����.�	+�BL��{����P�K�4��3�0�o~2Jn�޲nӿ^�^5�;E�㍛��!��z�}��<�z�����E>z�X�3�Rw�[V����P� ł�����/6?�P\�;�}..�HH�,�/&5m;�$X�W�={yib�i��}|�{%veH��]�ݲ2nu�V}ƶC��;�S5j�,2 PƮ
kѸ`ٕ�d@�?{�C��U��n���*��K'�8]/�#�����68�#�����{[9`���뛇D*BF�m*�0#A}��Ȕ�6�|݇��gV�@�����h�U�@Q��U��E��SF�
�}�[�\�����b���H��+k��C�ތ��,�٧A�&M)U�BO%�N���`��y�g���Hϖr�C���/��Z?氪9F�<ԜOr�(�W3�� �M�ǚ\���6��)��N�w_�gv���N4��5��W��_�CE|Z�}�'�U��G���2U�K����qn�����P����!�.�ڊ ��ݮ�J8;��A��5S궻���#,� 㥉���m�9Vk��N�ǹa���}Pdԩ��ln�����aӯ����N��̾8��� ��t�	H��È\�\k>�&���yB�:��ɨ#�}k�z�ǭ\<��w�F}7D�)�0J��Cp��#5'�m�&Q�Sne ��|pP����0Q�#�Wq��Y�֘����v�.@���uYf	��7y�!2^�F��\�XP���i�FhG��݊�YU�����ȭQ�o�)���0��it���o���^7��>�,Y�I�]�����l��+ƺ�^Z��T��;�(�[E�E�E��tEbW�O�;��s��"}���ĸ�Op��~�f�q�X=7It]�:=-`�� �F*�]#�nVǋ��$	`jq9�Ւ�n�c����"9�x���:"��a]�V��HGQЍA��KM5S���Ң�J?�>�;�ۓE˩Hf��v���-3��=rH�f�A��������&U/�o%t�[�&b�O�w�Ȟ����m}��)�sx@��+���:��%���R�AN����"����V`��x�ũ��5QƄwt�L�w�#7����;�5D	���a��S�oՔ��غ$W9b�?�����	�C1X�+M8��8���7k�� �H%��۱��ط�Ϸ�Ռ4
5�3դU`��H�y���wz@�wy�-_�"9,�qg�6�,�c��Y�e�7����r�ߝ~�޾U{d��V��7� 2v�J��ps�� ���_S ex}��4�����Ϫ� �'��ZT�c�#�ݎ�P��6���?��$�؀[��5���E�Lz��3� mv�X���N���r������Փz1V}x�ϗ5�����O�X���I���lJ���g�K���D��m�/�t���²�fr�ŮF�/|}��ȳ�	MB�vU���'�߄���7DZ/��}�B|�2���ŭY�.o>�������'`Z��e�oF�?�VX�k���y�?�4y:K�����q@��ߨ.�}1�v�d��Sn���g����y&I�����e'>���Q�X�R\f�\��pc9w���70��ނ��\G��������y1�Z*�Xv���f#��gv����M�,�Vz�f���8���&�9�4rr������9�vP����Ι������դ�Ql?Y>|��������0L釤I8N=nO;v�<��ư �"SR�8)EY�P1|`Y�ڬ���N����'�aQ���
lI�V��d�E|z"�P��DR����\{]���{C�����	j���;�yt�5�h�v]S���N����{��6����T�fA�v����"�����&|k�9�#[�`8���A?E�$M���<^}]HV�r�i�d�:�����F�K��q��_�_3�9~-��̩��}8�ԺL#�kW��=���[k�_����S���=k�Fc�d6���L��D8 �-��TI%b+�o�?If��#�R���ud��U,6�P���P}fƃ���-@4�GV�S��=�OjHTa��.��&�K��~äp�خ��-����tF�6$V�g!��ݨ�.��H��i���{����m.��j3<��h�/1'쯍�"v���x���7��4�D��^����-2���5�N5�h("-���(�y��%��z3֒r�豩�.�Y}�M� �j>})���qU/\�'<��cx�5�!�4���i�R;V�dTz6��!s�]�������ϼ�p��MפlA��H�����([Y�5M��h��&��9�W�ߦ8�v��%�U��+57�A�p�����pi��t�����ĺ_�t��=�R��@���tAE�r096.]�@+�>ԕ���}���q?iJ^���a�i�[>��LR#����OE9K�쪶��gfå_D0F���,A���[v����2�vZE�C� �9��E���1nC�d�M�+��p5���}I��c	UJy�H�[q���?DMѻ&�^%z�kH�N�=/|�A�W�S:�W���ؗ^T���-)�쪑j	����|w���������/hr*^�dev$&��~U���\$���'�w7�jT���_y����0a�+���3#�Ԁ�?$N�7h'�˲��T� Ҥ~�k�fVl�+!�hm���F����{*�*�����K�S�ڌ����K ���W\�>M��z��!��Q�葝)YO�\�Ϲ��@�@��w����Ǫ��O��J�%��$�5��ׄ�����-�4����[�з��R4Y�&�MDҙS�X���^Fݔ!DN���/�_M_�:�8>?0��K��*bvKLHD�t�F���-���E�?2�{�i�������������S�:��-~�em��Pd�޴�e����nbI~�ͣ��I<�|&��O����_��(�_o�933�����=�bL�ݹ�O�$��s��mnv��2 ���`��O��^�0Lm��_�y���q�Y=e>}ܝ���O���^�&�m�+!�h�Ͽ��o�Gby3�U4Q8�FHU�aq�|ʧ��?=ޜ�?�Ej����ܒur��c~��W-�l��w��PQ��'n[SJ��!���5.�S~j��o=���{�ɷH���y<������ǣd�m,Ϸ�]�����M�����߽0-�(�v�v�%�=mʹ�ȏ��Z[�<h�z?檕M�ѣ��ߴS.̷��1ſ	 k�<���-�����K��~�w���_��{���fkv�B�>V�cd	$�U��}A?�~���>~��B7��|۲���~O��Q?ʢ��hB�V1��2;L�F"��?>�ݛl�����J��\��5���Գ��,��id%=)�X���j��}�s���	� �J�3�W
���%K���e��Ok�O��{'�:�*6��,�f�jP��js�Qo��Z���b��[��(<�t}���s��o����Ío�tzM5��KL����~�����|/��{��7���`o�$1<oc��V<k��K���]���a�JV��G�m�&���@
~q����%F8��ޓ�O�g޲�p�穈]����	�u�=�QĀ#��}�Ҽ�B�#3����u�SX��ep>�d�8�g���]G��.ć?��sj��a}�c��G=i��5jK�a�]9���%:�R5�����r��ؿ��R2�q����Z���ꁓ��9�5�j�}�i��'���+{TA�o�9��!��������᧙$�j����o�f�D֢�nE#����o��/��Ņ�B���3/ǘ����:��C�V���C_W{��K���t���9�u佨\�;J�;��k8823�(ϙ~,��6�n(���U�q,=�3:�C�0�4�I��г7�ƂP^�K���\/\�	p���'�.����PQ�����HQ�ʰhQ�<�q'��xCܵ��݉-u���M���}2�ݼ?L	�M��Q�-3�7sL��G��n��1�JνN�.�{m�!o.�d�3EE5=����r�)x��^�=���;9�7���cuܾͧ7r�_W+X�=Si������|޻!��<nOT�����#%��I9!�ܶ��\���2x�q�K]����r������{t{��.��-����,��ɹ������|��?'�C�[����c�T��D�!w^u�PH��V������Q�\��sי-;�C��� ��),��EG�n�W��گK�ː�;)n}��o^_K7����{5p���7�u��QnN���.�wlv���l�fR�Q�z.��6���/���� �����0;'w%97ћ�q.DĚ��L춾 *�Zvһ�`c����勡|i[�tC�ڄ��陙�E���f��5��Q>֣�'Jj���NT�^����=�iJ��6���V|�Ac��6���g�qҵ���N�Ǔ���$���4%fmY浌��m	��G�gI.�NCE���<7G�$�v�?�\�^��==2B/y���G�>��i�a.#�7ս�
e�yt���?�1���p��k�)��o��g�)���1����{�Nc;NP%�h锷?�d.nb4S�e�����L���-\��M�`s�G���Ӌ����š���ny��ٛ�_qLi�ſ��b�Z>�� ̂�l�|�E�>Ϣ��D���BO��S^>6����I׃���o�<�U.�F�,`B�j����o�u9�����y-���噇<���4��a!����n������k��.��BFeS}�K�~����SC,.Jk���?�s�z�'�ְक़��e�
��SG+�K/FW�d��V�*Ķ��Z�{��䔽�uG��s7��W��D���L*G'7Az�Jn��Z�б���^֮y��=���`^�b�y���i_���E6~�̔=�����m�	�J΍�i݄��9��Y� ��ǎ̯�bN#�P}�:���ot�2m|׻VC���(����=��vn��t��&ԗ���V�7-`����7�������W@E�>�()� Hw�* �H��tw�����t��H��"ݹ�ҹKw�.����{\Ϟ=.wfޙ�yf��{3藄����l�I>���k[i��f;#�H����� �M�
G��!��h�?��j�*](�ۻ����_.�Z��沊4�:��&@����I�f)(�r �����҂U֌�\�]��;��k� �$�l��|�O˖(�^|z��Il$K����1_?�.eXȆI��+RH�Ҙж~�7)�t�6F�`�:�����Q͇���en[ba?�ʡ��>�GW_�����d��/�H�[׋	zN�Ҥ�OC��P�&��'M��\6���B�Bkc�;Kq�,����<�Ϻ���`�w�%�ц�h��Nٟ-1�7��ۍ�cͻ�v~ 9�P��8�i'ñ����̟U��\�"�OJ�r�br�m��ߖG�E�6� ��J��7�.�s��*�"VJ��5����hRf��z�k�������T#�C��s��&�^���?(#/c���1���+��6��!ls���-���]��i��������ܚ��#�;uV��k2��Դ����u(�
�[˵����ǶX��muD���S��rT�5�w�ѩ��L�0�;�y�ʟ\�6d�X���-��"wm�G�1/�g�gZp�d�*a1����t�k�m�K����ɹ����5ҿx%�F�z������y�l�a�8�A�M˿	�#�9Ҋ׿g�E+��ϊ���(슰�.�7�_�.9��������䮳i��?j�Q)��+�����6iu&OP`�F6A��Ɣ[F���O=jϛ�3�;�oz6�?��Ǉ����ga�
�nP���0�y#�sC���ʅ��Ͽ3��|�%�O^��H�K�$���"�d��?��Ѷ1(ߤ	E��|>�����q�卟-}랖���?���D�V1e�˻��d���٘�-eQ��7�)�QT�p�|��節��,�$�:��
�e��盧Y;{y#ǐ]�Q��̼a�]�`cVxZ���X�������Q�f���B������c��Nm��؅����`Q���i.T�iԄ��RD���}���Aر� ����I�tr7��R#y��g4\~�i���D��`H�l�2�Js�T�#c5�W�Oٴ�� .X*��Ao^�M��P���Q�f~ �N��z�� S�v���6��0.��~u*o�Y�?�H���ʪF���=tJ_����_L���v�'4	�-���^]�É�
z�RH�=�;�����e�#�?�l��C�U����n��6�e��	7�'�԰�3���{"m�u���c�j^>Ѵ�=������j�kY�7
�qn{C
�7F�歶ܶ���{l��CyU�@?A跆�
*ie�-���#07�^e���N���<JT!ɘ��`Jȫ"���	��aB2)�!��Q_�qS�_��a����F���ב!bA���qWʷF,��=w��jv����[*�a��g�':���ה�����W,`#�ِz�����A���J��u��dw� ���ꚟ��|?RQ��iop%�X��P'��L�k7STA�S�͵��m�uaWY��ʥ�")u2�ה# �O"3漈��Ǖm( �=��w'�(�A���쐌��D:�?���D�Ġ�� �eEo��Q�x�.�4e�0�DK$$�c�d�5c��f8���(MS��l9��l>H��s9WjB^��A���DA��*i!�v�o��[#V�et��_�:���{հ�~u�#�xy��j+�����󧊐�����q����r.�1kP\8���m�T]\,HM\�ȷ�brE�+&W��3?&��G��Q��7&���˗O't]k��1����,o�*5��P�?��c*��/���WZJ/rlTu����%�r��E�o����Hh����1��?[��j����)��+�� �K��aO<�j�����;���Oi7M�A���h���|��a.�MTh��PjL�q�D|n���%�u�Z�>�����6�v��>2������ířJYt^�x,�(��kF� �S�@6�F��X{	Ɯ�4��3�	��{���8� X�S����2�!X�򊆳����G`*��ZqzO*�v�"��:\}�g ց����ö�p��Q��0�+eU�(B_�N�&4�XU�y���	E�!~0m�v��U��Eq���"�oó�=��W%�a�w���*T�;(Q�1�d邭wG�B/�7������.w9�G��|e�Wk2�*�UƷs�h��y�BA׭7�C{��aI�yQ��e��[ŗ�3�7?�ݟ��npS�8K�nVD����GT�薉W�C���[?��I/9w����Xj��76�PVR�YA*�;H������Mp���9iЮv��z�Q��5/ؙ�Z���L� ���Pk��#� �� [%��d6K�?�]��v�l��7���t� ��߷g���
ǁEѸ´�}1�����(��)5a|�;���8N[q��u�0��S�0R|/{��i�ԃBWH��OҦ:�q��Z1t�i{(�
�զs��~�5=��1�lG�!��-eu�+sb�A@#�k��iL�V��P�Wa������J�k�}�e���6Y'��T\�	&4�������ņ:��agջ�|��� ���v�l���?UU�Hؔ|!�])���l:���M�yIϩ�F�������
!K��{�" �
)E�"�+�I3 �+&f�S.�
�m+��n����CQzC�dc��ݟ�w�f�m���8��,�v�	cӐ^/�NZ�sL(�����~��!�N[��H�llC��ݟ��A*���S�^����3��ʜ���
1k�����~˛H�ˮ��J l�e��l?���x wX)���\��}n�+��x܄/-M��k�o�����U���AB�V���LG5�9άՕ\ <�*����XX+%a�Y��ks��ek�\��G6 :M��!�d��1֗����i{CV9�'p롕}��"�w_�-9K&�]!vj��o3�`��|�yA��ђ�_ '��kL��l�ai�k�����M���x�� ��؜jVc�������I�մ�!�Y��̏X�W_��#��T���W�8#�g��~�-T���;�L��-�[�P{��#]�`#�N��(��S75���a�3��j{�ʝ�V(�lE#Iw�M��RQ��b���5�r��9��ǃ���grM?AR5���R�4߾��=P:Z��f/������~�zM�N�4��N�Z��'��a�>VY�K�7���vUCM���Y�t0A����}�3XPy
���Jy�l;�xAo��w��U�ɓC^�/�q/��3��X��r��ߞ5C�gy
���)��h3�å3UP��׭��!��6G)"6�]�2'�:��j�Fk@��ބ�0�p����#�ڒ�19��V6������Kp��U@v�4o���tP��Y����nlZ�>"��`y�3`[��������Y�0���ͺ�U��6��*=ɉV%�X�3���ݏ�S�ӶLJ�69�Bx��;�����_P�F-�VT��#\�z��W�b��@*x~�`��v'?\�oVc���2��Ό`m���j��t@��>=�Y�p�E�f5W��*3+E`�`8������*�����D�[pt�~P��d����!�Q#�98xQ`�K�>ʼ�����ߒ��݃^Rj�]��^o�����S<=�Czogy&�&��Lp���4nX,3���࠾"T�HѰ��"6���C��o��2�~�Ӄ\;�!r��ԿȌY~�z�BEW��]]E�׾/�]J8�)ֲ�X��sǉk���;�"�.�$�层��1Ȋ��|��d�Sʾ��2�&�V��{E�#_�^�{�B_�S�4����R��i�v�+�4�u�|>%ew��vI�d�~�e
�`���q�!;�g�횼۠����I�/L�+�����|[�*Nnl��O��G��FFVg����fZ��a�������amk�,����0��aJ�bN�� ︾��m��d�I]=��9����}�і<���Q�V������:"��n[SQ���O�7<�E�	kYgbp� Y�v�h���o�@<�+����>���Q5��]_��x�������fW�n�N��~�Wv��¹^6&Yz����~�U�@a��v�igr���~=c�\ o�S�-2갛0i}�6�}���^9��ix?mÒ��F��;ҷ�V/��P�;GA����)
k�ڮ /���?Lc�����ŧWs��z{�����(a�1�t!�Xҧ�����[�H����&�|���F���	�e�<uȳ.�U?��a
|٫�"ET��5l�v�e{���yuѵJ��¾S�vUv��d�%`])9?���`�_��Ī�<�_��Q6a(��Z����kv��Z���Ú� 8Y=w��6+��I�Q[K����.pQ�9j2>wþ4.}�J=��w#K�r3V{� �j�wJ%����JH�AA	�M��P��K��c�+�ZK��c��?+���.[,�n�2.�䩿����a��^���O���4�f�5=ŵ,s��
�~��ߤ�/�'BO	*N�����j�E:�S����P�����31�Y�������C����B�n�Ϊ�������jMӇSA�o��c�$	_���*�:�O_�7"moRl//���=][BW������D���(|��1YՂ��~i�/���|�%��8��91-L��=ۻ�Т���c7��gƬ������1�S�e�r�/P��רo���Uf�����(t�ޭh�C׳�$#�Ѱ�s�Ym���vR����1���Į�#�{����4���&O��V$~� ��Q�躤���[������*U�Mh��b���Ě;�Ov��!?��E��D�$��q�n�7����K���6�@�$Ӂ[A����^����Rjo�7�3;�a$i\�?J���o#ѻY`���';B!��C���� �D� &r�i�mky�M��/qOL�P�B��Q�8j�����X�7��/$rA��;�sƙ��}4_�^HL�"������n�)O>5�9'�?2�=lE�^����e�.��#(�5�����
������d�=ˀ�xnu�	T!foRS\�2�E ���U��op2����%4��O�B�lu���u�QY��]�yyh4� ��y��Vn��!$)�+R��Hа!��J3�������/7�n��P���#���I��U����'3np�e���ee��_3�$�0�YYU9��JCwR�y��⼑�q�l��Aj�h�ġ��k�R�q=͐��( -X�z��$���\/�MT�|�>�����郦s����1h���'�P&����f���ͩ��G�MDH&����'5ݱI���ׂ?_�B��C>�&���܍�%�1v�(l~x��7ғ����ک���{�u���W�l��KH�8��ʈ�e#�ÚL$ݿ-���~z8vp㷝vEY������.��ɕ|2���w< �4��ð���XH���pZZ�8m-I�ņ��_�KK���OU�8��[/�IEɋ�(
4�z~p�3��˼��B<! /�9rN��83^SE����'p��C{��4�����Fn Ȍ6�~�w���s���%Ue����(���U�?+n�~�y7�D�U*B�` �΍f�-R�"(������+����[{m�q&'�w��ZE���'3|U��6H�����9�|RT#��dP�ɖT��6ݧ� y�lGt*S*���4��2�DH}�sחH�
����������Q�j ����d��ggeu2��C�7��Su��>�7��EF*��%/9�.�V�q�NJX1l>>�U�� |E�V���g�Ƌ�/�;�қ0#���ݜƝT�νG۩C"L���8�dv:���R��
����߭X����M�"�Z�Y�>VV	i�]��g�G8�Y��gGF-zu��(�2��x�I����q��.m<����	�b����V��|f��&,��07:������G���0 ̯��OI!�C�6�2��}o������OI~��(�./v&��t���p��9�ý�ܬ�H9;I�Vp��Ċ@UN����(R�L����� Zr=���Rr��^���ǌr�1�h������7�5�;3��3+�d��R��,�7��W��燫��s9 )nW�Vr����^W��`u�
��B�֔/��0��7b3��*�,@t�|���nv}/���ۙ�% �Ʈ
ɓ�&7ަ�㈌E��3�FEW��d������X��*ŏ��}< v]B��L�����m�i>�l[���.�(�#���`$�~�����>��gf��$U�� ^� ��0�z\���)�1�P�<%�'-a����o&Vi�-дI���S5Q��ɛ[�}���GSM41��֟�-h�%X�MD��.IkW�Z�U�ɦ��2>�4.��8M������I1�D �[�H/�fCMJ��O"�<F��+7F��b�0ܺ�G0'��$�$�9*ȉ�U�rہ�d�xe��)�JI{ח�h�,6����L;��d�2= �������;Ԝ�&z�V����m�$���e�Cu8{�Rϻ<�+7'��Lš�8�����nc���������g��b��^Qd�4���V��B����$�@���k��ldȢ���7Կ:�ԦS�pv����r��jh�_O���������aWr��!Es"T��/[S�?Y��(��QF����h�{������:Hm��y%"�_+f믻�}����L>%�3�)�=�Bϲ�=�1v%1���ۑ�i�/wo�#��;�U_yh�|�y�_h�����S� ���J���bp��(ҹ̣�U*������Y�ն��1|������g�G1����/fuHv<�H����(3HI|���ژ�m�����t�cZ��2(c�[��7��cy���R��o	�&��Ƽ!��B���.f��~��
+(ޠ�%N6�@K�z6�y���6m+��"�C�A8�{���%��𳎛b-R�K ��ѻ��*���j�H5�\�4�K`y�X��3<g��!7UD�_n��w���~�vwY��G�	��?�q�ʏ~<�6dŋ��:K+�1����F�Z��ܯ��
��2,z&;'�r�\�EX�4�U�Φ=t�~ػs�n�R�����jI��/�
ԪE��]�~�)��‖�G?LW^z[~��Vu�z�
#v3��d���Z�U[���M��MWa<e3L�p�c��du��&��
����߳����*R�[�4�&�ƨ�����ch���ά�<����M�M. l&��7^�ͤ�ռ�f��CYQ�m�ҷ���%��?�4��~�w�@a�"ax0A� ��XL#����1��:�Tb��WC��g���@�y����I��d]Q!7��S�����jW&cV��?�NJ�ny})���ēP�D���5��M��Wg������ٳO��C�n���m7�B@X|'���}3�QZ�@H��],>�3֖�͝���*�&���������h���d� ��ï���"�G����Ы��v�fw7z���`DZ�WÈ��%:��Ȳ_��c����DQ.����rD���"/���'�0sl2����������ag�ДW��,&�d4���g��Pc�w�K��=�xy:�8̓uZ�&���[*�
����-�H�����՞wGa��'�"ހt�������=��#N�nY��æv�ew�羛Ԉ3An�&;j��G����IC�,��4��"�ע��^�k�@��Kܗ�k��Sl��B��e6�H"~O��2㇖b@l^���c�9+F.��~�MoI��AH��~J��t~<�q���ny�s���m[�X Dl�������]�OCb�Cv��{��{���M&����U�k�2=����k�_�N�cv�ǣr�y�g�Vp�҇,��ry�B��0\�>�[9�~�P���4F7��ɿ�|���M]Z��r�[� ��;�7Ïi�6��ae�=�3�)�ݦ�Ϫ%VK0��XEhK�o���+�2a��=���{ըĲ�z(Rf�Aƒ"HXm�^�w,�L�jA�qg�q}W��O"_��5�~,�@�-I7�i�ԁ��B�I%M�g�\A�k�x��aD�Eȳ��|�~��8I��e}�n�t�hb?k�[��u
���\�-��A$=�eۗf5��=;�Ƌ8�y"Gmj�#$�S�tP{�����]l�<�������Y��':��A��1�O�~^�6c�uu������$`tl �axx��m�Y8�ħ�R�I�vg�Y�k;����P1k��:˴%�"ѳ�?K�������6�~@�R�*0���M������j-ֳ�BV���^|>�V���5|T,�OQ�Q;�t��Z���0��ę]�y;7>e��E�]��C�4tG�
'��I7����Si��Z{��l��\:�o�+�C�v��]��5)����nG&Mo^��;��&'"��_ \��Q�O�Vv"��l��8zx�=�����;cLn�ko�~�!a��A���8��7�@}�g4�\�3�,b�J;��4F��<�<S��{]-!a�>pi=|��|Դ�9F�l�5d=U���!T��������~�N,�m�땦���#  ��
�EB�v(���k���P	Y���Z���ɥ�ȉ��3O�d����������+z�D����s���f=��׮_�}��T�zx3Q1��PV����5S� ���Qh��忭P��O���Y�	�b�eR���v�m��9�w�o/��Zz4孩�'��/��hdB�Q^����D'k�h�m\^`�N�4$ o�����u�\�*L�	����Lq����*��8�M�O�E��ۺ�Q����"��qP�W��Y���3��� �A�Kh��m���G�u�ϵR�GĚ�KU��a��!��W�>��'��K���=�i!%�� ����ъ5g-�`�g���sh��1��D~\�r�-ֽfu^����9�W�L(l5ȯDz�é�I/c�E�JFG̕�> ��hK�vK���m�oۢ��\�59h�^Α�1y���IM̿1���96֫ifv{L���Z�
��\��df��g����v�O&�k��'M���ݶХ@)����S	�8�����Lz�G`͢� ?&���� �* �;NB���b��6�J�+�p��n'+�]�q��)��Y�zL������ U����q�a�5$ !�� Q��GX�u�Nq��|O^�Nn)��T�^�����sX�M��{r�rLW�Ӎ�{F�Q�5j�<�����Ƨ���*��]}�<����j�I]�Ѣ��"Wۺ� @�d=~\��8������yz7��'pjt�FV�\�7<�e���-Qw�F�}��_T=̺ۀ�ҙ�ؓ�]{���?��<O,���Ħ�q��0�k���u�:�d��$ۭ=M1� l.�����d�.\���¡��r-��1�~R����$PȻ�z��(JK���ITx���=���(V�OeX��i�_3�⎛�Y�N��MTZ�-P3xr�R�Gvi*|��M	L[lMva�
&{9х�����rv�mp�U��=k�뻐�=E#����e�,K���ϩ���0n���mQ0�����j�М�:�6�����Κ�!a΍ǚ����P���?2���+x��O��+�d��h|X��f~��J���[��9^����Ӵ,��MdL�� B�0pP�PhԀ�S�d?�廡V�`k�i]��`����0��8�<̎钨>x.�@�@�	�нR[�Y���^/�G"�����;N*K�E��Q�&��( �BwR�h�Ģq�5�M3+ �T/�/�1�|� ��wY7�/���'�|�)O��0d�57�$�|��6��� �Nv1/Q��z{6(�bU�a�t�t��Թ���?7+��V�S:�| z�L���������c��4�5�<bۦS�'�d�͘.X�C�dzQ���]�~��+�,�4#U�WnB���&2�<^�'�\�I��_TJ�Dڈ��el�dϦ������$����$PL0�l��	~�T��/���q)p�ϝTl���積�ڳk���	�p�K��ߑ���{���N�N��)+ǟ<M{�<�jDÓ)��k��aO,��X��nE�O6'�t�X���ң#�/���R�F��8]�)�J��['���X)<
��kv�*�z�II7��w�QhNL�h���>@�J�r���y���ſT���+�n�>G��
���=5��h�c�9���1Pr�m�~.�R�-J#I��!+|{�ߌ�6�:�i�ن�p��5��קW\a>�E�'���Q��eŜ�ڋ����K�Q6�\UJ����v����-d}8I���4����c鬕��S�n�Lc�T#�f+nqt�t0Wn�q߼�i$}Cr�'����m8Rh��c
�
�@"!7Xu*h	�D��{yi�J�N���{�v���&�3��K�V����<0�Y�Lr�F�a�Cq�f$M�ӏ���,��ZV�TU*Ƣ[\.�՚�c��ȧT�*f���\��z��1k��d��
�Jj*_��ԛ�
d�d?<�zTP��̎��ke��K]��U�PhN$Tf�m��(|�Z]���XuYQ5�^/�I�jێ��;�l����G���E풌8��XBJ�����"kEj`q�Lp�ߩ�p���bA~bOk}�%���T�3,�o�Ig���g���g�E�����59\����(�9��x_!��^��[h�j��R)<���e�� ߔ~���p뗏�����߮�4��a�:gDh��t��c�����o!�̷���Yܭ�F.��ʙ�W����o�%6q�?���B���u}-�-���a�vz���2K�
5���S�7l�f}df�ݭ�@#ә[�+l4��X��:�1�:<���0��c�7�8��:�]{���I��/^"���Wn����N�r�'JRïg2��Č�L�N[:����$�,7��-�up��Oo���ش�WN��l
7--�^��26|q��L�V�Jq�X<��5S�x�,����Ƞo��3*f�Ә'����ɭjNX�u#!��Sߣi.X���L��+X�ׅ5��t}�к�nV߫�@թ^3���a���B4���'���D��e���ԇ�b�Z��e7�卹5�� ��25&ǂd�P�u��c�?��>�)ɕ�J��`����Q\>�g�{��4��M���o�/&���,o���	i�����K��a�
��_�4[����ܡ�Y��D��,u�m���v�b�K��+`�tb�8���=f=���H5L����0.�0�Ӥ>��	x��/{�Z��L-��n;?���}�p5R��K4��5��b�D��|Zr�t���d�? {!,y<ĉ]OǣKF׭3�xU�HMg)�u��5�ߌ�ף<�e�W�l��cr���
W��@�V7��1y8�,���y��-�����lb��{H��ߌ��Ū=�ȫ1�Zk�$@[��rȊӦ¢��7�t�P��Z�
��r�@΍A�(|���;��C0�&��z��쨻�U�.��$��W�[?�E���z�� ��?�i�K�3�P�'n�_��� ��y���H��6�>�G�)��l�N��0��lX�Pu�d�-Ȓ����A^|��ۺ-E�� ~���Z����L�0�'�X���і1�H�̤�X˶�w��Fک� ��Y�ib4a�7���-���
��g8Z}~)ѝf��e36ב��'���5� ��D���Q�㌍d�V8`����T�Z[�����O2���輪���FM�M�����"�������_g��w��dN�u��P���5{��;׬�Nlvc��@	?���I���.IҶ��%�ra�S��_�v�R�u?�k����ZD��р6��4�y��/W��B2*<��#UsH�5�����fЧ�Y��LIWp��"H'xv�>_�$�n���,l�&������m��v���j3Z80���f�r�ޤ��B_
,6J
������C�����#d�j������ᓕv�	9M �exY0��͜]ޛ����fm�j�IJ�%c@�ӆ>�j�i�7+�^���sx�^�-�G��(�Nk�k��J����x�maT[2)�/w��[��C/vD���^���T�:|4��x��`7�J ����Ym�jAV����C�Ut�T˭e�47���/���[j�-���]W�I,2T��K��L��B�=w9U�d��������L���Bq-�Zב����;��aSq�/>���J?�p��I��4����B#�Iy�'�;{D&@.�'���I:�����c�r�����mְj���6�ǲ�![n�(T�$�
͢OMS�	+R&��䱶�~���^��[����}-���fV���f/�0�뾥�IQdV��|r!ޜ�x~��gO��q9��+Bg­�\Iu�,'�Gw@
ɸ��J�8m���Y����G��'���}he�C��L�C]�.�+�6�
5��`aOv��N���w�7��i6�5���"�sen2�@8&��+�c�L���WueҸ�����7�e��֎�w`L�ơ�\Ԁ�t1W��}�l�"�v�m�:K�y^��2�y��6I_�J�~`��e�lqO9����|]kƁ���Y��.3f�X�m\J��"�0��,`�#�t�ӝ��^�	��5�B�����j�$T�w�����~F�&|	y_�6nm���.� gRszI�� 
��kf�j�>J����­
Qe�Wxh���o��Э��H�Yn�Ꚛ��|_�:?����t�}���|R�d1%�~{1&yZn�G� ��fm�@�͟��<3�U �{��(���h�,�J��1���f��b���\���.��'�����	���cx쌉��a�B���`>��F��`��@��SV1���rq�h
:����Juj���ܯ�т⎔_��y��@o'�@j�p���S�}�w�� �s�Nj؈sn�cƔ�
�v�g��|5F>b����h�,ZY�5Vl��k��|���|���,-�ļi�w;�q�Qf�#���k>�맏��g�2�R�"�g�) ��ّN�w7�����|���#I�$8^�t7���� x������w�N�t��y^�Ӷx����X����۠f�FH�j+��Mr����ß���C�kQ�T`=�?wO���
���}L9Oe�泸0_0��lu��%�������PI�1�n]��s-[ �i��9\jj��^�1�wr{����dPk�!+D���y�zr���+�O|!��&Lq�s�i>�w$Ԛ\z�GY�J�b��G�V6�P�$"{8�Z�P�j5�8:��f�j-K��\�J5�Y�oh 6�m<�s�-�4�r�gϫlg�mО�ScF���M��P��:_�I���L|�)g��7�hw�fsm�u�����s��) �d���S�a�ޥ\����;��J�����I��x����zS�%Ł��I#��)���y>��N���
�N-і}��?�q`"������L�m��f}��1�� Cr�H��}1����������oI�	�W��W�_��~���K��o�j��P֪�pW������F��\�f�_�B]�ܬ�w�Z�T��w��V�=I�^-I,��T��x#�{�q���,�ۻ���K!���_r�׈��$�'7�@�:������0L�	��j_��������"7�sd�Y�h�9�)�� *L�(�(�ON�GO�o��2D��C��;�}ҋ˭�������`֟7!z֕;�T��$Ǚk��f ��!�� W;�߇�u^{j׻�;�d`:^��$�����;<��q���%��c����3�{
�᪣w�bS3&��y�B��;o��^\��եܠ`�6YB��n�_ݖ�ר�8�C<���<�.���)*���咏E�R�A\��T5�L��S	K︕�]:����n���Yg��_�7�٨�!kH���E���L��v�Gd��)i, ��5��1p�֙�Z�%1We�xJP(�NjJ��{nN�Z��ǥ>8��:bg���`&�I!N��Vؤ���pD�[xf|��p��Օo��i�~�����G[L��U|�3���^�`�f�-Ӓ@���N��<�/-t����X�Fs}�/�::�b�n�}�Խ�>�85��tG�c�4�����|٤[j�s� ��۬U᡾,���������1MoNg��'R��/��j�A��ϙ����e���� �ٓ� �O��ɓ�FԷ6{�A�"G���|�g��;Տ�:]؅��/�2$L]#j���<��_OV��.��{����4Go�"�l�$]°Ļh�t@t�����"x	b�w>-���?�i��j,�c"�L�-���`�}\G������a\m��D={��>v���w�H�cTi\�61���{}�.�VR���2M���u/W��l�wl�芛��>:��6zBީQ��l`&-o�e��:����>Cf�*^���2)�\[b�ˉrg�y�0�&��_n�8�5#{���ݶ6>]D"��&۬?�Ť"���ϩ��n'_���{J�#����D<�D$CKnv�s^7(�Ĭ�z���D�t�eD�4n8sc�u�h\����T��(����4��p��cc����S�o	�87�>��ѿ3�*8��4H�=�
�#��p��(��A��.S��y�$d[P1m~�?;�h��B=/�$�Գ)��PH����dr���M&�ՒT�`IB���?�Ȓ;��g���裞6�(o�M����yK�T����Ek|Z��E��w�II�JL�����%T!�I�}ضLS��6gGs���<s��t�L�x杏��n<�?`[s�5Fo��y������-e!Gy)qk����p�L���iJp�"��h��F���ߪ�Z���k��&�T1�٣���t���0�~赜��ǩ����г�
��{�i9
�-��ܳq}�H5���^Ѿ�E��?����o�k��T/�m��Y�^�M~�����Ǘt4�V���;p������ ��ٿ)�*�aZ�w��`1��f+�,�s��0����X���c���C"i=�6��y��b��f��r��J��{S��o��6j�ㆹ@lR$s��tҿE���M�X�$�gr��o�j���n<ˬ�!�F�}t�K��uJD�5������JO���݊��8�kSϚ���/�u�ql[�84�N�f\�]����z=�y�i6:�/�N	r�)P�*��W�	Վ)��u�ΕrJM�Z��3D9�d��5 Xn��ț�$?���u�(���G���AOك��(�lQ�_�]����z�ޜ!P�oS�g�K�����E��ֶY)o�Z� �Ԙ�'VnbĮW� �M�d�Jؠ�ʾ:FʢȆ�2tggPRiG�k$U59dna�8A�+�7�W�9��|PYe��!(MoJ��z7�-K<�O�A��鸡w" ��)��"���:��Y'|y=�H�I`ȏ�O� ���C��T���!�<
�o�7��)'��/�]�����ܞ��O��(����G��F�
bܽ3h��{	�t����Y� �0C�������{�D@6&G���_NaA��2�:��"�;�/�A^�\��[� ��s�p�_5����؍U���k�.���dg�	��d�Y}N�/�<�m|߆�4�*j��jW�o�K��p����<�����2ߤ��Z����ٛ��4��x.\�k�t��]b�}"IbՌ�M�r���b���Mg�>���\�a�3^�D�/��<��\Es:lNjaK�"�w��hp�A��1*�x��ۥ�ã�ַ��}N�h����5�Mxqξ�;�R9��e�e��d4,���B205D>؜�M�a�ӹ����Uv��5���4pC_��=���;��q�6�=[g̜$\W���� �����
	����u�6+K���H2�l	�23�B]�����|�L#gy�Ʒ�X
��b�er+3�É���H����j�&�(�)�KH�q ��[@�怙ܾt�l=%�lc�c���X_)6�����X�tgD	;�-����kMk� :���BDO����@y�@�	��_�&O���~�7�S�����xC5����¨|�o���
l*�o��w�o�����6mh�_!/3Bq�w_�q�\m�bf�[�l�\�È��=�w�뤌�&�l� �����pw�iՏ
/º��v[} �Ů�8�Q��X8�@8$�h=qw����.Zf7��1��$_�%��$9�N	��j$B�Z6��^�������� Z�l��8�˄깯c���NP���J��_O1Q����k�Ч�L�CW��?Kgr��&Ó��A�l��	����h�u��ɩ�u0 N�\;�~��J����5k�w��EP�� -?T�~�8&��X����w#�6�h��۫���L5�f'%�����7�2BJ����}~�%E��)��_n~�j��Z�$	��Q|����Gq�&���̃����:��zIXO����*��ή���&=��Bf;���37І3���P֛_ :6�;ᬇI��5v�|Z���ЭM ���^��G�4ۙ�M,���}�<ϴQW�C��H� =z�7���ؿ��r�y���F�F�^�z���J)p�%	�ME^��{�ay�������Eq�'du�D�ڙ����j���!�釲�F�� 4}����wni~n�l�٭�%�oO�Q/:Suyb�:���_ǘ���	0�>��wY,tYU��0�GQd�0�g�����
�&����J�EABT�$%�A����Α�AE@I���k���" Lr��n��������\�5�s�s�s?�s?��<ȣ�);@ůӯ4I�R����k��=��{����J�H5�՗(�<M�q�w8e=��^��~h3d��Q4��'Ȏ�/��0���~��{a����l��� �����I����������q�~qj�((�B�N���)eP՘s/���l�6��)ы�3�nt��T���T����t7��A9kgz�9�ګǟN�v����GsxE���kmЙ�!h�s�q�PsC�ܡM�D��feF؉��l}�5�X,��5+��x׃I��Z�Y�J>qbKv�C����T���K�X3���ː�3�1��'�Z�[�;�{en�ݫ����9~�5E�ij��M�t!.D
��i�tJ�|v�j�ż@�!��Z5G�1�,ļ�� ���{K/Y�����y9�ߚ��ܧ~k�Na��u�
����IA�O���tjLR}jV-4e���}�$%��t�^sXSq��4(������)���bq뒑��~�S6s�M�K��u#\�*�-����I�ⴱh5���P�d���܄�|���A+������R�ue�#����:l�r���J�UO|P����t;^��/n���x�c0���Z5q�ո]6��gI4d������9A��1n�߸�?Nţߩi��� l^0���+�A\aB�LCp�5���M�uE�7]�?�Q?|��g�ib��K�ި��h���^e�*ذ:�R��dC4�ks����
��sWy'�����k*O����3ˋ{b�V�9?��k��y��R��ˊ"_F������e��F������ȢY��Q�W[h_����ox���KTZ�-� �ma��[��ߜ����iT��:9m����I(���D)�y��p�'�1�	c����][�|�S��}����ϟ�F��<�T޳��4��G\�;� �4+�3��TСP���tU�|R2����������iF�&�4k8�_rͰ}�T��n��0l����O�Mo8��҄Y����%�^��aX��a���W��BE;���.��a�ְ4�[��ȆF�XX�m���K��e�8����������Y�\/v�(m�kd��#�~%�']P���m_��GtS=�:�qP��x�
譟հ�(i��m�1W�}�Ѭg@Ȫ�{pO!�=�L8��,�N� �2I�#W�ܚ�I	��`C��� O|!y����G�i��t�XHL��.f	A>}����{"Zw$��O�j�����;�D||���؏�!s�L7�,C�L�6�P�
���_�������gse3�@`?�i�>q{ǹ�S���L�h�Q
��� �km�QM�V��AsZ�)ҍx6_��x�/�Ș�G��Z �!h;�2�q~6����~CQ�O��$�16�?�[?�F��@߰�N�@q�|ȴ�a���@���F�*U�FU[��%݄ "j��*Qp���mΣru��
�l����Y��}�旾��
~����N�8Z| ��X���GN\�����L�!��=1�n}�y��A�X��CIS�"vcJ[���T]�R:����O$��U�7[EeX�s�( 6�ӅH����g0���"L�g�����ѳ��pjn|���8S���}��N�\F�V�,~~"v65*�^غ�u,��>tKo4[�RA�eB�C�N��JJ�?�0��(E�D�E�s��6�\��|M:!8�v��g�H7�τf��PD���L���y'hF{nm�<�b��7���M�F*�CO-dP;F�h4��'�R�¶Kv�1��������
��^/�K{��~dkb�6�0���X2�����P��<�O�@�`��U ��8��J5�,Vy6�������X�mܔ}GT��D��5i������@VlQH�H�n&�������)�?��c?�V=m��}�ɾ8��A�Y��I<�io������Q���|��8ä��{?�:u�0h��_%V�)����?:��ج׭�>��9l�BG_����V��]�p�C,m<6�r
�sz���i����`�O[�����c��/���H=88�f}O���

歚���;��	bn�QD�5��%�l��_N�����`�C��l�ƒ��e��?S�6wGr�	�hF�����k�C6A�x�h<�xv6~8ee��d����2져����w���+���鎖��ke^Oye�BQh���M�J���ky/�K�͍kS斉%G�ڊ�N�dp��F�����m?� �}f�[`{��Q�Q��2���!|O���hRc/v���ܹXS�&�'���~��^�[Ŝ����~&gg0�n\���Ay؅	 ��H���'cD��^������>Q�
�?e��M�Vg�4��]� X���xTj��9Y��`JDө��l��q�<R��'y��G�	%R��T�?.���]ށ'~oB7���_X��'�ŝ��~�	�p�����L����=N���0q��TUUGY�^�
}hr��Y��Jb�s-5btlynܵ.�YW��%E���&�:�������`85/9�`!�g�;�^]�2�!k4Y��-��PN`��e�rk�s�L+}Ҭ���]sJEwaV�����l `��G������������q.��4�3�Q?���>�6��l��di��\Ɲ�Df��F{��:�b��yu��܂N)o�a�g�m������7��5o�����jy{�� v{[ޣ?�~�z���ǘ2�e�?������PZj���N6!�S�H������[�N��V�|�'�8u����_D=���7�r<��M���儎EX�_��� ����ω<m�m3ˎ���L� ����d��N��'�d�`c�=1��L7 <=��(U$����h��_��jB�C.Z�Zu*��<�pT4Q�:�hB	eS�0E���E�#afIA$5;	Al�hS=����A�@_���X9�<ĄY�[�h�(B��Ukܻ~}e��B?�VNJN�9A��
+�mLtN��Ʀ8�xƧb��a>��S����2SPWu��U&i�4!�_YE��#�J�J������g�aN��]��^�le	�!�1.����][������P�k�C��L�@��������rӘUy&����<Ys���P��B�XZB|��7mxa-����:�#��o���O�@�������`ޖv��C�E̰>��΢�=����'oO:�,iu>0!H�-ּ��\xDo�'��`�:���Y�`7����Vs�Rޒm�G���D�+����摄������s��򓤺��a��Z�qN��{�R���l��nR?��0S�j�k��tz�gT�J��BH�'���oǧ����4{��U&�70E�ƫYv��Tf��a�h��~w���'Ɠ��T9T{��&OM��3�bi�[=�w���Y�.�\����� �u�ynZ7Ρ���1Er��&3B�/ڿk9�%e�G�!M�'7����#��<Ծ3za���ة�� !�ka���ʓ��##�i���{���-�����4���L�㔛����;��cv߹Slэ&r � �o@�B7J����vyG���S���k��7w<W8�<������/<�cai�|&����9�ɝ@�N� �p�]�)������zݽ�E����)����8Ό�h��v�R���Z0�p�v�;�V3�,��y�R��1���[�߿����p�j���Cb\�C�΋mt�!q���
��N�Z�^����녒� 0a�U�G&��?�'@Na��}Ί��^�uܤo����_ܸ1;Y鋓�fX�����s>n�����X�Fc��m�7�t�R���R�4�rw5��C��ř�Kz�^�!�Ĺ݄�H��G�]5b�%[��1��g�?�pl,>)&6�ߢWC4�Kؿ3��+�EnG�{��N}�����o���k�����8Ojt^i۬	?\�H�|�-̍@M���u^���k�j;��j��P�q�h�A0���|S*m��p;��uC�$��3gS ��e�Y+-Q`��C%&=�X��x�
4�+n�`�ώ7������&BE���T����&� ���'��#e$Wz���0�V��J�FI�(�Ѳ��/��Z��D�u���_^��;<�e-��*_he)�^�YE��S��^U�����ʈR�&��vxӣ�Ns<Ȯ��+���n���JT���y6���k��<N݆�=fK_���N�#���Us���r7��@#���ɥԝJ�_�N���~	xQ`�
���ˍ�oY�R��Qp�q��~v���Mf���Ѧr�>Bd�zCt�Y��Bݦg�~�0��~��R]6�E��,uX�M�b���aG�jΉ�p㗼��o���[�u~�%:�
�Y�%4~���sLt��C��Fݣ�fC M�<����ӣpǶ@ў&W�?��^ۚ�rJ������}�61t��4��{�&��XKvm�����
����F�%5�[m�~�M6���AN/�Ƴ�8\��&u���^o�\��;c���5���D
۞���k�8����f��3�=VK/|F��EX7T	����U;��|1�b>޸�i��yk{@��6�(>7q^@�.S.8�������!���~���I��^tn<���{�p����w	$���e��2�Z��D��!I���3^�F�2��3��@:C����u#��˞[��C�0��$�_UA1�i�_ZbD�AUǧs���KM3�������j�}]�ܖ���=�憩{E���?���7�����_i?��Q��ӉM����{V�q@���C�mo/���/'�D��˸ ��$Z�?����'/�3�"�`��e��J����=^����?3|jD~A&�����<�d	�y�ƻkO_n^�)���g�e�=N
!`%���k� �a�醲{QY���� �� �����ѩ�,��W!�cm������#Q�NJ��Y���O7�l��m����l������c�gk7O|l��n�ے(���~M`����A�������W��G	��]~#I�r\B�ˬ�NH�qω��5�Կ)8N�T�[C	��+����H_���M�W��Uf�Ӯ�^ؚ��\lE<m���'dGܹ��v��w�w��<� '�#���bƗ��ѠNx}ه��R�=K��jD[tnz�o�Mt!l��%m(KC�b�JH��Jl�҆6/N�EF�&�����Dݞ�[�u��s�1rV�x���̿y�sݥc��� 30�Lm*�{��2�h]]��.�$�)uS>k��y��١�(��`K'���H���}�?���z�[?�m�o������ZT�<��8Ȕ�a%�5"I���O'�c=_:��U�|A��:B۰ǂo��JV��U��ޅ8'-W��|��+�m.���Vege2Uo��X��*�v	������7�|�v19NMSX�}�ST/Y.����9��<�hIY�^W ����.���t�S"S)�b��jq&l�#b3��woHl��z�	%e����{պ�lD �K�����?�`�i���&Kg�8�Ha��*r�%7��F~��N
�m(�����Mǆ���߽2駟;���[�o`�-��hM��ש�a�Afv/[Ak`/$_I����ۅ�o�s�w,���Sl��@��?[�;�8�@l���8D��z ބ�i�q#����F�w6�[ҺF�Y�,�Q�������:&�;Uc���|�@�7��R�{o{���@�G�O�wV/y*1���[N���3[�L8�sc;��D=s�z�+1���]�;��9�2�,D #R���G=+�.C����B��~B�GY0=P,lbj�[(�oeB��6�yؾ�4mrЁ���5S�]JJ�����MV�V�a��A�b���,����1!��j��m��$�%�����s>^.�V��KJmv�&����N/>��4���Mt���Ȟ�|�K��������ty1�4��Z��GA����֗�wq�O�|w��x޽'w^�x�w����s5�t�����m˛p�5ѣ*����~*��2G��<̧�������hKy���|��<�Y�K�X��dS�a�z�X�N1��Zyp�ԒЀ���
�9�k�����&�ּ�?���3�����ŕ�z��M��H��C�o��➮Ϊ3SP�㴊��_��J�W�f���DQs����F���1Ð��;�Oɺn��#�U~g絭�=m�y.�W���袤c&_v`SFS1�d��gjw�D�H2�"��i�AbFh
(�sn�t�9r�FQ�x"/�1�
⨽/s�5����<
Y� �ذ����R��8����'��5e�qX���d�����T@~[�pi{���)���Y0MoJ�,�9��bB���v���8Z�=#,��A��H �n��6Z�BM]�<�r"�K�z�>�"��ӹ�^g,ؑ�7�6~BBI3<���G{=��ۛ��X������/@����X�RjF�6�r�����C���V���R�g;q�օ1����aR�dԇR'u���G�D��p5���|�V=�O��lސM�U谐���f�0� 43мU��We�^]9��m�����L/�Wﾑ�w��&`�����6���I�Zw�������D󖰒��D1[�~y�N�Z�N�w�g�IVi�O��D����J+�/��,7_��x�2��}�o꺥�|�_H(�1_58)�*3Ū^H'��6�?�+�Ϡy�8�ã���:�jn���v����V���3��}X��ՈT�$2�0��?,�����iw����
��pBN٩Q��=bi��X�6�ґ�'w�EFa�3�ub�V�JJ�������_S�Q8���x��4�*V{ �����`�F����i9�y�����2
����'g��U���T�&6?"�;->G���Cr%��)C����TPj&j�*[%�b�\��[�|y�#IC8�LK�Aރì��j�Mo�&�8�� K΂W�HYc�ü�J�M�8�ݓO�"p�n���r�v~A�'�/����tK����["`�G�	�6Rr�-h�:|@r���!��R˸�G!����g��@��h���mB��ĒҤ2(�H'�dl�R20F�^OCi����u�c�5E�a�&=�<�Kwft.�"�z��>�9L�Y@-�(1���G�����HPXص�v �*�O0�tӛh(��n�R����H�E������e,�DjG�5���ɧ�*d�#�i�_%�5$�o�2����I(�����A˦GkMOL_6�
%���K�7M+?A�<բ{⊟)!"5qIC���p���ZuR�^�<ԄrϦ��n��L�~��%��d��(������&%G�P�_�:�~���aؠ;��kI%#zx0�ˣ�����2����\��1�F*z�^C�n��X�DTU��td���*P��Q#�_�9�(ri�����l�z¤�]W�#���4Y>B��x�T�����s�W��b���y���EV$�}`�Xz��-M'xE8W!�3�5䮔��y�T�=�y����x�	b;jݥh��AtOJ�bƻt�'z�|�A)X9=�� }�3N-�"B2�/�u��J5��`���q��(�v�4��"����枱6w@>�0��@�X}���E�W�ϭ����*�R��t�X���N�\�;�
�Iz�=[�L׺��X���U�:Hbjۜ�l�"�l�?"���o/@g��Ss�3��*d�,症�Eۂ�D��sg��U ƚ4ȡ/+:�,μ�ݦ� -bT�O}N�u�xU\�X�M�d�M�GU-�j��w�_:�|��"�>��L��$V�31l=����,�fb�ߡ�*����� ��M�}��x������~�{b�f�c�~�����f����҂X��Q]o��
)��	��Y{��3�M�jY4|]QwO�{��R���8�̲tV�����zh�;��v�1��]��V܊��0�����?��-׉����#>]�_l<z�"�0}���h'�9�n��ϐ�#1	ɞ+��<��V4N⽍a���UQ�tG�(���H�הZ�6��+���yy(s�@�J����SgޫN\�.��*<�T 5�|&h���G�cJ��-��k[O>"�jݏ��z�y�kS��U����!;��O;1�!�o,��.�wY�Qu1Op���Pֿ|y|��ݘ��^���j��s��g(Q�z�2�������;a�LH�E��=[�5�x�4y	uJ0OT}�b�p���gM3�6�vU�.��q^�w1;pnKײ����V�Q�:����& lރo \Z���C��������p���ZuP�8�D�7�
o`�]PE��ٝf�s�n���v�+N�!6�)�Ey�6�9ž�[�Tu(e﬎�Q0/�-r��2�����]}fn�!�5��� ˟/�x/�������?k��"yH�^���uZ*P6�����Q-Opm��xZ��A^rF��U'��� ڮ3zK��/ͬȝk]*�g�D3
���\��Vtھ��Ɲ$�"5D�Z_DH��I���HH�~.mr;��ߛ�V��P�����3�n��j��$KN\��}{ f^ 
Ǯ>y����p#U1���0� ��t��L��N�*��_���מ2���뵻�S��v]��QC�"�\G9̞���V���,����k7 \�8��H��A��Tj�<��xL��X�έK�y%�t�)?/Ya�d'y�xX�B�ާ �CѴ�+�T��R�2����T�����"���p�eA/Y<#t�����!ٴJ���d�r7�_��k�
�P ���]*XlS����3b38)���p�B�J�5ĢR�a�+�;,�n�X'=����7<���z��PGI��9��_l�Z�p�z�XL	TTn2���uQ}���Z$\�Uw�C��a��PXwT���q�V;��͛��	bQ¹�$q�VHpV��~�K�c�喅;�wὪ�x+#�y������w��z�r�qC�I��n�~��ۺF�Aޢ}��g�q,�F�nIy��\�� �_�|�sn4�R���S��Nq1�ub��1ǽ�s+�W&y�Ǭ#��ɣ�v�'��-)Q,R�L�����Ǧ�_xfv�� a�Y9�������۾'�R���`�/�%��b{�"�#�v��m(�^��$�6fa�������x�-0��F��G��/�c�ʪJ9�1�P�8��$>(��[v�B�Zi��c}^��z�X�Z~X�J���J䍞�=���<ݞ8�:����g����y�ɜS�bõ���%ou��*�p���r�jy�#�XQ�{1�գ��J�������nCz+�de��қR��lx}�a�X9�yu��9J�m�i�d��}��y�1�g� ��b�e.�` �l�y��S/��pPy�g�h�n��՗�skL����R��GZ��	�9J���N<����}������f������N�"�D�6���/h}��
��
)ٴxZ�W�w_Y�:�ĚdE�.���~^$�|ʰ�������ݞ_Փ��.8�gѳ�Yi/�E�W��`��E2lS�a�$�[�w�[-{�����6Jm��ᇳa#�
����ڳ����Kߠ�X�R��l����e�ɣ9d!g�����a��cǐ��"CL{&����e� b&�@�*�������B���q���ɾ��P�.𚊑v��РQ�+�$��T�Ğ��O�����.OܨD��M���s����|)������@ō�@֡�b(=�*=���8�\�Vq=�0l5�s�9�}��K͎T�
ѵ�§уD�:I*�K�.�jJ5sЅ��'%�|�a�,u�{mM��C�����[8Z��2KZ]7@�@`����v��;j��\aq+�IEO8�^��K]��Smឈ���O�&s�vru�e�������sEd�使��	?�R^]=���c/�O�fř��`�*EA:\V_���^�6��5)&o����Y�*ϋ4�[S����fI�L�_��8���$چ��m���d�:-	;y9�L��J�Q�OR���y$ߞ���U��~W{lpT�f}�\tyB��k(�z\��S ���w&^˷N�ک�-oz��$J?+��ۇN��H�%K�:I��1�W/��4���NOg܅U[�o����E���t���.v+�>�6�����*����V�P8�$��և33�itH:<���8Ή��YB- ��i��.rr��R�+��WkE��r�VZ?�c+�	^s���p�͜g�hk2��AڟnvuM�C5^7���.$�4_�B��k��$���`b����*-n���?W�Oݥ�wr�{��u�w��;�m\ҝɜq	��z�w.ʹܘ_�;L�>��`����{�&���aK�B�ӛmeK����I]e��Ip��aE��n��˚���\�]T���]��������S�@s�B�#�R�{���oh�Se�2uۀ'U�+1����s�rf	����A�8K�|(�"��ñ:��c�'6i�� �Y�c$1�<�IѾ���A˄�uR���w���]���l��1�[�9R')t���$h[D~��+W���W��0ʰ\�@6�cVw���6��a��x�zi���<�.�ˆ",��.��V�,�H��� ��9��!j�ލ�?_\�#�7e�b�i��Q��$�R��U��2HS!{+�
�L��[I��{8�@�\�?���_�x�����O6<����Ry�kY����9�S��ÛϜ
�ֶ�ȫ����N��ep���S�������eG�v�!Sj�a��=���Q��D]~(����ҽ�}��-T(��E�9�ѰdSP����X�7�ҏar_ku�k0��O߲�&-�.�)s|r�kp��,9��A�=���ӥ����rK�[ޠ*N�l���|�Pm���C����})
�YG��c��]T	OHS��6ڜ�n���d�ޞ��3%T'_�i�|��2���1�.�mF��d"K��h"�����L���yM�R
k�+8���s��sf��HI�Y�|�t������֜"4
sƺZIz�MR��߱N�����~�H�[^:�;?����>u#r�2�Cs�����4�DÄkuir7��!m£���ѹ�:�L�K�{b��0�Ș�߶��*�ؗ|ھ�&�-���S���W�I�Ê��'�v�w|S�"�MD&�����c�*�>O� ���%b���2�
Y��V��Ƅ}�4����yֵ(����.�����ko��g<D$
�z�SV�h[��x;�<�"V>�ȧk
�p�W�N}ڀcT��&l������7_m�ª����.o���d��B]���\o�*ſ+E��a*���D��P�ž@1�F�(&M!5́rk�_��ћ�	�0{�1.�L,�?�R)�[��^�% ���)Nx��Y�p��p�\���x�*t�ħx|�Kǯ�?"�~EG�ljO����j=*���;X�|�_3J$J��佔�	�Z�,��h%���+��Y�]��.Z��uA�I��˂���6Ź�k��8@%ZG��M�C�C�70*m�ح�`�b��ש�k@�L+���Z��A0s?X�?F%'�b�/yM��'���3Ƽ�Pgp|�c�-�f��b������X��N=mw|�BVծU�GH�1>����GY��!�?��%�������������H�hHn\iY\D���<�_X^�[?���l}��b<�?�ͿBՑօkl�`+k˻���٥��-�!4p����,.\+}kغ�����ϸ�)�z�Q�+�2��送�{~�?�I�D�mn�wV��If����݆8r�+��7c�B�B�dp %(Ͷ*�3��`Г>.�A$=�Kx�إb�Я�aG]V.�cSwVU��X����4�qFT& +��'9� ��/�.t��%B�����;�|�V�3Y\f|�y����'M��7M��(�}���Ol�e��effa�~��}Q>_�������l齃U㭯E/��a�#����������۩0˞�յ��r%�\jO�� K�l�J����M�Â���I�hvD�PHVoZ�� �
#�qym�%�3����A뗬�3�u--�R �8���,�ߚ���A7,b�pa��As�O4�C�	f������(\��k���-�2�?g-�:s�JHIy�c#�=��XL�ed��q��p�K��q�<�vՆ��O�W�����L�U(Ye�9A��
�]����e`�\c�Lfk��&��/�7C�b���Ў���ݯ*�~�w��ե��Nr.�sYcqZZ
wc#aU�7�����S�ږ��{#|��,̊���䕉Dĉ���K��O�n)��/}*��IL��+�c�ǔ�~<�3���>e�-�ǈ�z�|?	�y��*���н}u�)H�4�(�z򈂁�����{�'
߁������e�����a֏g��������Z� �;��vĨ���*�^T��������!�?�Ζ:)����>��������<���h�<�I���$� �|�t��̪���>Y�~��]��u�ŃiZ��H���������>��,�N��F�=�G*l��1t4�����5���nW-#q��~uYlv��9���J����|N���Ҝ�['�d�퍶v��g��Z9��΍��s�FHV��B�T.t��ΐm˔.�4SJ;�r��g�K{v���]�ۥ�}�I����U�mS�W��ߞ���9d�ث��a<����>zy'K�g2�X����]����q�U�}B���2	S!�)�#ϵ�A��v�8i5K�%�m}zu�	�s֢�q���qI�Ԍ��B�?�i���'�;�t�~[�OLstYzUfK��V�a|�B���In�؈��A4�����[�?�<��,}��d�s�H-�)��'�!�@	���럚\LF6�F9�=�h9���5��V���$(���J��k�2X�����v�6Kxt�D4�<��n}�O怳����&Y��>W�T�L[Ssdb"��ނ%%���.���~�X�����v�ڈ"���#�IEcr����9<��i�v'��D�%�ջ��y��b�ㅏ�>*`*{��Ϊ�t��5�,v�+dWe��^��U4��G��.]����J�A��0�;C͕���������L���Z�';�W6��Y{�o��U�[u�k�$:L��O�})n@v��?�=*�;ݗbYY㦸!-�Ӕ����!����*���7�̑��p�X�*�6��T�u�7{�}�9���Zǯ���������[��݅P؈��B	.�D�ΐ������9���d4
�N� ��G�v�c�����`�+K|g�@!�>��*[R�0M�zDI�7|�K��t��RJ��$z�K������~c���K��A�ܩf&���K�Sa����u�'�3ś��K�W�|����d�AY۱�RJ���(uC+ nA��������\g��k����/y����OgP|W6{���_�M�ۈ)w�x��&8)�L2�DX;��#j��O6���Z��/� ��2N8��*?��\����$�PJ�k��̢$��a��+��)	�k�U�����q+rv����驏��Z��uk�i0��u��pRT1G5�xI7�*��Q�_�'S]�#ʿ+^|L%���l]�����e�?y�C��ӽ���5Uꪴ+���K3|��#J����=!�����H.eb�k`6/`�M5&m"`pF�����,G�ɕ�Wk��3B9��sɖV���1�>w~�jVD5�) g�Ř����B��!�q	������l�o ��^������M�Ð�4nE/DoZ9�Ĵt~��ۥI�-J���k~�����N�{���ى_�[�ro��G_����b�{�������L�j(A�4�nr\�.�=࢓�ž{��.d�_�tkbFΤ�B���N�Ї��,+��M���+J�5���x��AƊU�B���w�o�9�>C�Ml�>M�(��|��+<:�ùP�7��ٸ��YBe�+D�?������sʾf��M�!�Vc�z�#m�B�h *ע��ɳ���?��ϖ�Ò¥[:��a;��a5ҖCL_�S�~�_�=�#�Ǐ-XN�W���Q��.\�;�����m��]�����oKw=v��N�=�e�MU���z2����ݺ����\����Ý���d�fL���d675��Լ���fV���DL��2�\/�:�%�=i�����=1��4�3F-�j�7�L�L�`:w��}�L~y����ɺ�nr����t[�_� -�l�	�u~���sgi��h�#���5#h�ٲ�u�H��=H�:�o��j���djW�S�^�Қt*yQ��#O�|
�x��ED>|G�A�&����T�I����W0hu�q����7Ơs�9�*�`}b�IM��4���T��-~��|di*��E}��=�\����&�n[�ʛ�\$�oH��Em��f����C=��#Ak!R���Op83�
��x�d=��4��F0�ǻ:�*q��B���o]՝.��%��e_�٭8�����<gw6��>#<8a�>1-/��Y�
�g�
hl��<D�hE:+ �]�Z,<�64z'��"�#A���ݝ��h�c�cH/F��R���<�.�j@h5o�]��*E�I'���.L��?g �16߽�f�����P�\�:�cZ�;�®˒�?=���;�
Rï<ʁ���ϸ��������@����Ē���mb}&������Og���V��ua��	ZL������G��3������xu�e��c��j��6ҁ�!�o�UF���5�Cb������wm�Nܮ�D[KHܡ���
����	�p]�@�2F	�m%�	k�~]�H/�_莗wm�45h�H�ni�f䢊����sQ�3$��\��G6`<�ˁD�����dm�.�����m���2�k��&��6��A��L�.��r�@	M�B�b �<��}R�.���N�;�A�&�_�����V/�L����dI��PU/0��o/��1�7��Nc�m��.�U!	j�=U��H�`'y��r	B�Gh}�ڪ�K\�!j�� $IuC����j���I����dߓJ7t���6	���Z}
�u�5fb�F<㪸�]��k�����XG��w�#F�깚�
M���N����ͨ��A��Ir�6��H�0j�S�;E���!�y�g��:��YY�O��E{es�0�6�j�����̝��[�O����I/n kU��M-w�#ϼ�J�� .+n��?Ҭ����Sy��:
���}�Ժ9���$���?Sx*���~���q%��,W+8$��i��?v�Z�v�k9�Xs�4���}�(�=`����R&�1QN�;��GZ�4x�iA��8�%����O�7��`1�0��t������V5��7�4�P@��l?Ǒ��@�_F��L�+t�t��.�Y��ΛzD�B����i�?�7�ÊJ3܊��K�h���vF�̙&0��d1; �(PV��O�~�kW��Ax_Ѽ��E�����Ȑ���=V
^����+_flO����r�^3�q���Q��]V��n|Vk*m�񲻨BoD����M�ݯ��Ռe��hhh��TEz���N�;�<&�-��Ҟ�����3m�)�
S���D���Y����I.B ۗ���62��4�~�*t��^�i�?�'k�z[y�b�:Ǔ�~F�竡�ݜ~�6Ƽ�pŭ�{NuDn�&gJ���,���|�`ei]xx�a�u��Jd�#�K���G>�و�QRY[�헜�����@���~_z�5��?+l��&��J� 9�1u�	p	B�J��PY����?�S��"�p㭢��l���%��S�AR�;�fw��O6�)W5��ui�O�(�Kp�*����W�׽a�j_}�D|����qv�1	�to*;�1���x��}�ҪY酯�D�D��'����	fUy^�OcD�P\���;��Q@b%�5\���W�:��dR,p�GZ� �x��)�yUr�]7���+���#q���x�[Щ����B2�m�*Hg�֪�l�I�����t��o���cX�Ũ�}.�y<���im{pc�vգ��7�)�:kU�Qث7ɣ����|%;�ؗqK��Omq�
����jZ��#���f��(�8�l}��	��v�2�H�\�=\���ϔ�K=��Ej��W��>��@�*c��"�H��4�XrPJkn���<��-P�N1{ª����N�ۏy�q������Zi���2qtI��}3*rdc��/IɿK����m+o�V����/
����=�%�b��y&��vu�H���Ck�/�	��8���y�e��$H�`!�LK�����W_����NO|�ʴDV�q�&To�!Y��������C&��JN��-��".��Lh���YQ��%��o�!����x�8�V���<4�d�#9Z1+�������Ur�=w�s1�z�un����WG��n�NL�f���;��f�;(I��K9���U�z%m��8���
z5EMc��p�t.sd~�R->1�sGJxOIpo�qn�?2�~���N��/���l�i��l��@}+� y�^BmM�h�z�������H�6�����F�f\�kM1)l�$��G��O\�(�SǶG�K��<�]Y��(��6@br��$�B�����$��.h��ߌC��z4�Ŷn�������1�i���o�m��̪�����5ްo���'�����!"|��8���5`��r��!g�dېdc� ��T����ո(��ϻ�t4���q�Z`�Ы��o�dy�Cא_��L���x�c	���~�T�uX���>�r��4��E@Zb@Z>8t7���I)i���Ai�������~�0p��{]�1��콟��u�{���d�����L���7�����PY�o���S)�;�`Q9�09x&��Y����%�p�ay��Ur?��,͜�3��~Pu&Ǧm�=Q�\po1��5f�I�7��~���ޥ��+gqrݚ���{�%_@�6�n��̪�ܡ�V+AZ+o����X�$\��j����V,/�$��2 &Y���~�保Oy=�h���ߐ5��>�(� �q�Gq�M,,�a�i��{����kZ���H�0�Oee~��r���Im�Ɗ���bl���Y���bB���wU�6��T/�é<*+y�)�H͞����t����3�F�-�?����a�'�2�*��rS��6e���)Q�[��FH�5�~�]B����j�[�u,R����'�2��5�9����y$��ϝ�
]rq�˓SṂ�9 ��~�O�$�������Q�0 ��~�c����A���ΙYY�q#�>��-q�^���:��n��{?̴��6�����60����Sp�������D}I_�>�k8C?^]w���--Tu[t�(�5�˷C3�>��\��@lё�8�$]�縧Ɯ ����@�緩��Y�㒀�r��^�����f��,�w�"m��`ך�gC��C4s��� }��w�u�Ǥ�H��3�<8$"SX���ɑ�yΨ��L�/5CU&Rp�V�q��>�g/*;���}b����=C~��|$��������"��yͻ6�_�q�pok��a��|_��dW�9����>�j~dX�_]H�]����C�v?��z� /�M������ �,J��|����y��HJ���G=�,�`�r����`x�Ȣ�=��Q/v�D:-�����ыgv��/�Y�yg�Jw+����e�������eF�6�bO���m����"�k�]cGݏ|�oҗ���:~U��1�4Q2�6��<�z��>z� �\}{��>�?�/��8��9��{��1�Pp�9h�W�uQ�'���J�{��K5a8���&��Q"Zs��*MTs�Y��9Ւ9:�/�j�٫;���Z�0���	ͩ��@��ُ5�>Kd�3ZG��5���OW�����3Ym�g.�ۖ36`���2-ȏ�l���.j�t������MƓO�'%0���@��zf���Z!�"v��&�0���6�� V�v�mW����^κ�����h�	�������]+�_ӽj���mYAO���nw��M�rF��4�ء���6�Ú��.&[���'P�tnQ=K#�u�S$�Ǵ�a����w|2���N�Z��_�Ӏ@M���`����qn��
�����}y�;sή�F s�l����WSy� �%�m�
�ͼV��I�`x���k�7�[6٢����D=��c�h%.F08�_�H��u�J)/��R�I�'ڝ|�3��Y�\X%��_��d5lp�۸�|c.�z�\|�6u�x���TNjw�l�޾����v�M�	x�|3���dz��I�q쏧�&��Í�B7"��ji
R;�g�
KL%m�U�����a�ө�Ɩ�����)��2ߢ�a�1r�OA���[��65�g��I�zYuK��/`y�0,a��ZO�Eh�H�4��&��`��"�p����oj/&�Voy�1���|���k��;��+�#�Y��6�]?̈rF���㶵.g.�J�sij���[^�k*�0�ӐV=e/�N&W:2�d��(�~���qu��X�XprV$h/�%�s��!�\}nXU�5o����X"/x��`�x_���Ǆ&�_V���I� A֢֮2�ѫ��.�2Qm7��р\b�0"Y��D��N���{��5#��t��N�b�!ѿP�"���r&�H_��~ȧ|�GP9�,��O��o�&�?�Nkz4�U���oVZ��*)T���{�m�T�ٟ,Ud}o1�k_ ��E~��t%{��1�W����5.�����5ܓA���O�u�Ň�[5�Ø���-�Z�Dy����GA���s#�D���#!%���}Z`��[���STs���3�]AX�M]"�=�"�*y���A��	r�'!*���x����6ɬ����ٽ�~Aĸ#xr�d�u��5 ���i[�������!�t�E�%�!�n������������\,�-P���<_�
?[`3d�r�J��2bm$ 2\�r#�:���$ǂ�e9ʉ�+��@�m���Խ�ؑoG4>+�f�05��xˎ���o���{0\s��\��[U�x�*��i�b�D�Z4t�i	<��KLٶ't��zY%"4Qs�z���Q�k
_��n����]�����P;Ə���$���ik���-���2'S�-���!��kG�m+���9px
њ��%�(I�6���[���	.��k��sfzJ|U�a'�4i���Qa PV��	:�4�A�Ƭ�l
�y6��8��1���F�R"����e���Q�5�"RoR	-�g�ʤwdf|�I9`Z��eԳ=�@�Hc�Y��_�U����(m�5$�I��Z~����\}�y+�����Ȕ�o���,mL+$�0�a�R?�\��zhTِ��n�R��p��0�͙�M��$�S��.tJ��A���d�1S��O��;�}��s���軐��"B!m�
l����gR���Q���^g����ϔ�3=��sy�k�#�y �r�]��w/8�������	�2�l>l0fi�#4�~yN���7f9�QҨ���A��f��`e�	�ԛ��p�삢�\F�=� j�"ݟ�_��WG��>g�T���#M���|�^�Msᙒo�$.��c�������j���O�g-<^�j"��S���~�G��B𱯣G�א��N�G!����\;����>��7�ג�;ݸW,�%�>a�*���b͠�vfȼ����ݶ*��-V�/x���]�a�'h��f�M�d�6b�RA�3��az<�r3'��\7�7q1��ѽ�ԡ��.����5uٻ`�	���*yc�芚�2�)�%�G 
ٶ��5+�"��a�޺6���{�Ý�#�#DQ�98�E�%���%���C��*v�3�"��:"�T�j��eG���) 3}]�c�Z�M�������%���Xa���0�G'-Ӟ���8Ѩ��8:!�ν�eF��f�}%ߜ���QA������}A*�8*̂��;�*�h9�5� �
*�bv� �Ɣ������79���F#����Mw������g-Ж��]c���7' �x�l��D������j��'/�N�Zv�a�K���A�Ҙ���>$Ӽ�����w	�54�e���%�'�I�\y���)�Rq�ಣ&H?+>d�%�h����(�u���VV�8>9hF�f��DAEncv?�@g�]��I���غĤ�ʨjTfG4��hf�w(����wC$��CÂ=�5)dY;{�q�U�Wg>6��Y%zc�]���5)�BP�"@tߜzْ�yFig���Р��O.�d�"�h��ؒ �> �i�
LչMs�Y�(���|.�Uw�����ϵ@F\�w����-��$5�=.\4./C��ҳ���7�V�d'!�[�yV��2�H�L��"C3���Ȏ��j��9��&���I��#� �qAe�ַv:�6&vL�YH|æb)A�La�KX�^v�����i�6�)�ތ��5�o����]����^��AUlF4Ź�O���+wփ�h��?����h���C3��֞���d�j���˽����f��TKO''ƵQ�М�Ώ��ϙ�<EFC�`��|X�����2��}�]A���2�6�����ތ�Z�#�ӑA��~c|�O�"�x��pK7a��*��3Ws��N�.��@��4��4p򩋩����<q��k�����"�_tW�0��t>t˖�����FQ���·�6̙����M��d����~���:�K� �W+�tr���Y�����5U�|��N��
��`�����'�'W��:� H%ٛ�ڰ�τ�Q�������>7f4��'���_���$Ŷ�&5��a��@S�����s��`�\�+����A,��^��L�c�
F������T�S˛�:{8��׷�^��^�3`�`��B;��8iQ�Nt��x�P�<m����vaQvb�@�ug�:�|d�>&����Q�A�� }7�-�J8C�:��5�+�����yC�%��;A�X�e����͊L�I�ݐ@�#�J+�
1x�S˛��`�\�@q�J�p���Il*$��ypV���	����S�yv1�b��a��s���gi�+*���1��Ig�����u��@P�������o�J�/���[�t�p;oK��1�|'Ųa�������>��2�+S5�{DK=��J_��k*��mqfg�ֈ���X'N��&�d'��S2����/Yq�s=�3�S^�;-!ݓ7鬠of� �D�/�j���J�9rf�}O�:�T۔��	g�3�O���T7��V�b�.�1�$�-Zg|ܝ���CM�x�u�B�$VW}��3��oLF[hzR��UVk~�Ѹ�I^�ɜs,��B���8�8��������D�Yx�1����SK�G���T���k�T=4���s�ܣ.�#�aZs�̆B�,�{�*�E��&=:T'��#�Y�7j���U]����zO��XUH���C���'�����QSǲ�A�Ep!�ْ�J��W1�Suʍ���X�Ɣ\�ap��ze8�Pt2n$
��4!��X�Z��H��޸�>s�������U<�-����$NNS�+!�G������2����"���w�<zQg8t��{�;(�b�=WDf��U8d�ꐖ�kd�����؃������p�]M��J�V�E ������Ȳ�<���'>�zXT�.�����HCu�xw1��fd��$�l9]ubU߀ut��Y9��w��V��SXXM7���oD�DU-�Z���"�s��[��� �(.�Z	/�7r5U��k^�9��H���Y��c��a�������ND:}X�>�ցw >�+�����p��ⶅ���@�a1Ɩ� 6+��׌� ��5�i[��a���&Ph���t��zh߂��E��D���xz|�g�tTq�/��������s̚QR�P��ԅ}G�#��АA�T��p$i�p^>��WM7G�=l�.�-kN�lq�z;G7i-~�m��~k~>���!I=�ku�eg�	yb������|>��l������5��	��&�ɱ̱��oO���Aό38k��g�$9��n��P3v�����l��s�mQ����ګA�`���۩7� �N��̶x�:s�쐵~���ޜ0f��_b9�9�K� �
�a\��V��#��)� ۂO�R�\�A�1��T���i�{~,�v:;��#U�O�_������-�~}WQ.�&G����O�m��D�I-��I�Zsmv�-�����Ί���{��!.�yx�\
��i�[Eo/l�/]�.6���G��?�A�s}�ڥ5̽�]�T<t��h��7�0d�f�*ɰ4hµ�fҗ��ԡع��S�d-d
V��Uἂ���o�a=�RF#�P���L�<Kn�`�V���~��.eΓ��u��۲H$�~�)&7�x}��:/�>0J7��uaB� ���S��4 �|VFDjp`�D��e��0]e8*�������1�{d�����H�\��ͭ긁{~J�������lP�0e�,����D�Kd�"�-ʃ���:7g��X_7y<�1��3��SD[2��"�|�7$�o���܉0^��ڼ�s��={�L�@���7r�j�έ������U���9�����} i�Ah�&+l5���G��p�@wg�f�Il�Њ�ڢ��+E�9EoS�ݪT�K
ª?�MvQ7'�}��@y���Ug2��6^�A�8�����rP��k��饓g['�����"ֵ��Qg�r���]c6���a��.k�|�x��U�#>U�Ǜgoc�_79Q��}}�ˋ����yNr�!m�2��TNjց|W4��ޢcr��
� <"<[��.�Ng'��o��I'|*�����O$���|K\���NQ\jԥվ�#;Ra���[r���y���m#vK��d���9��']�_%<:�&m�s�>h$¯���>�.W�*+dEںy�r���*,�Ճ��hL]M
�GL�<Ts�<�_2�̊����Φ�cl��y��k�#g����V%'Dc�Q�^n{��$r�K#�`Ҽ�[�'V��	v�J���������.2?�G m�W�k���w:ZH�G����]�����(�+\��Yf�x��p>��X|�8]�ap�5? ���)Mv(�`:t�����nB�j���\�֒�[�w9�M��N�q�,j���eE��F!A Ryt��8�e���?��{L�Ԗ��=��Ƨ.g\6F]挓a�c�r	#�QT�pXP�.�QT��f��A���G>WMW��G&�&�kSr�"��J_L�����@�84��S��"�)b�0��y��{O�([ޡj.y����_��`��9s��S�D���I۔�Ծ�r.f��l_�xWA�g�R.
�۹��,�)@�@�U#<���N,��U9�zzl�"MnϥuQQ�Q�L����{�w�}�>�A��l*�rW�>��e/H�z_7�0�"aL�؟�<��������c`pe��b(j�����h�"��3̜u��V������٭�t(L"���e���p_NR���Y�y����� l�Cm����=_����m�0�]=�9�w4�d5`��z${�w��r�|����>��=M=E�WHQ��ɵ3���k�b���*�>�!h�E��s����CT�U�����A`�w3��L��X굜i���A:Yd'M*��"����dU��*/�j��}��Y�XLV0,�i/�����$[��݋��#���׾5v�L�w��~U����띢^���V� ���FV�:^��D4���P���mR&a�I���y��1�r���K�~�l��.<�25*���7��3�r��8����)�dq�XN�(Ԟk>R��M.ڳ�MM`c�o͂�F��	��u9�z����*�#jv{)C�]0n���"�����P���ݩl���EG�ݏ;U�i�3b,j�	v$���D�Pu��n1ŠK�2rn��ҵ��-�ˍ\�E0�B��p�B4�5���p��W^ѝ
t�7u#HT
۵L-U[^=K��Θ&HH^�B�z	H��y�|����I+�vj`+���=D�_���u�w&z���|g�0�}� t�|cl�kocӎX�����B�n����G8�D1�DD-���n���D�g?��6/&���E��np7�]�OK�~7���ɎH��&�uJ�i��,��GJ\,�MT�\��M�֋+��r��4N�m�Sv��'93���>�O��kqKZD��_��:"Sp倾D���Z�o�SOS��σURϣPU�P�zg����Յ}��$q��R?d8�;K\�#�?��	dF�`��Q��Q�i�������P^q��' �H���� �����z�:#�~��mw���v��EM�#5�{�[�d1%�b��?h7|�q� \`��R�d|�?�+7��۫5�G�����'��ݓ��O��>��]˻�����X��,=�Z���8��ˋ^�����).�Μ1p���l$v5�H�TQspY�����q��.�@g����QB|9S�m���"�����Z'��暟J+�1�-�Ը7jq���]�t*N���_]�:m(���J^��s��@;��q����#Zm����KZp�6h���s�4�~\>l�ށ��A	�ϻ��0X���IhB�����g�������w����0F�7:-ܝB�h��h�*�6ǉ�vW5ꔊ�/�F�d��I�C^�~�b9�G��%�E���p]�&��Eg����t��Cԛ��vʢNsNЩ&s3�峒� ��� �h�;F�sx\��Eƹ�	3�o�	�u>H��k8�	��{C�ms��9�rB6���M���/��G�W"��$6�V��~��kSѱ'K�o�:6Uc��dy���c�����VH������gI��N!�Y;W�=4+���r�Mp"܈��"���@?�=�����Fxt�?*����S��9 �t���U��n漓#j\�q���f��,�þ3�v��mx�'���P���rv��I��O�*H<"G	vY9b~~4�ymt�C��9�rz���a�Кm���5My�� ��_?�U5����1 �bd+�����D�LOq���� �Bv�4|kI���Z\S���j\��W�D��^����x�r����߱J�_��0.�A��f�إ�C��|�ڀ���W���V�Q�&}g��z�ј��m�-��Ҥ}��oj\�n^F���c��Z.o��[!q�l.�����()<R��[С��ۨ�keU~N��nT�8��αR�����?�na�O/7%�I��\u�PK����W���$��ޗ�_�dMX3Z�t۴I��񻄣���i[�|;����(8���q��a ���f��UKq�Ĕ_�eL{Š׮x��ob�Qq�n,������{�E	
���+�[���`}�+�^���e�#�����2��Ze�D/W!j��K�uA��1�q&����"��vt��Fx��Y�"tj	9�ף�I/����	qf|�|Ĺ]�����l4�ȫj����_A�'zT��`��w.~k����y6��d/�[rv=� ���Um�E0q�x���O�^�˟�_�m�/&� �%��ca>� �񨽲U��\s�ҥ�(�&}�i�0�yI�?]�A�"��q��b��ȳٞ�f�Ffۤ(H�K*N2��,���/N]$�oh%�.>�ݬXLS�J���
�-fZ]U�]�(�ڭ�����5="�X�xΪ�{��g?]nTg�J$\׾.��'��A#|��i��O�![Qշ�	ַPV����j��.B����>�k�:a�̳xC���wK������>�pĘ�%:�a\K�	MY��"���k�[G3dY�:;G&�韖U!`�\iv��O�""��6Y�n��h��1O��A�\.t����P[���P����6R�u]X���W�o�<�HȓJ�ʄ�,��)5����ڪ/M�GK��S�Ӈ�3����t�i\�nݕO�襉���x�i���S�J��K;Z�w���>�.TIܦd�>K�DK)������wG�<ђ@\W��L_hRt�3(��N��3L��z���s���$'�?
�m}�`����N��=�?h����� �����c4nK*���\F�J����^k{�c߼[����P� h1�_������}V�"����^��0�[r��n�%�g���)�o_c�v�{�ȇ����K���S�u^br�{.�ʷ�10����~�+���˭���8�;K�?��=�m��I�H��ß`>J�̼�Sy��>��JoVԶU�?(���B�Ol�� ��v�p5�@Q
:��Z.��,��zow�����XkE�T���	���\뎯�Di\�w*�|�v�=�.���Ĺ�J��~�A�Ït5l���3-�����8�����`�Xi�t
*K�y����).q���Ϊ������f�ɭ"4�'<�
�1���u1R,'Su��X�{ɋ��_�܄��R+r��5��=�ey���ݘ��Dh2zHuӏj�$t��`��[�?�%�K%�j�B]�;^�%��|�[��S�SD_Y��Tږ�+�~)�Qo�1��r�F;��2�9��i?��MO{)�=ޠ.p"�P�M�C|U1ss��íT4�+���6��O��"�)�z�jW�q]��Zi��4;��a��w?
N��V�$�.
�~���o�y&DJ珏n��Fx�M��gc�3��Go?�8����e���\�����Â����˸�����1�M<�l��D'?�4�F*\rT�W0��x��U�B2��6��{w� �����J�~�L7���WR��GL�(O��\��6.8�i*���x�#�]ß�#� ŵй2s�(ƞ��)�W��w�Hj�M��ӗYA�O��F
�φ]l+�>�ryZ\��je]��(�ku��O���*y��ٸ���g�ۮed*$�kR%r���U{�'T��*,�*P	y.���M�y_~%������Y�ɩ42/a��5�W"�����].����$�����E��ZL��^�8l��X戴�� �0o���,��� �T�TՁT��Ʀ�����;gM��I��Q�E�<�uH�]�!��R�ǤSZPf�yv��E�0sɺ�a"�دpt_{Ɩ�rm��6�KVh���u%}ݕEz(��Q
���/|=ƭݪ�B�+O[D-�n��>��6�N��k�o�z{z�Ϗ"�\�_&�L��Ų��g�2��F��}����B���V�2�j�ו'�ڌT�l�U���x����O���*h�r[-Y�l]�~���ɾ=+Q�&<�����i���X~�4� ��i�I'G�M"�m�g�
���0��?�ZZj���^����}|�R��Mc��j�����M�%i������nE+��w�F_$� =��[�\��E)����p�71d����u��?g���i=FY��{cW�[��oFdd�>�.�}/���(�����[y�mÃ��]�$��99Tޣd�+��w��/�7ͅ��<6QKfT^������I��#ȅ��GIl'��^�-�o����C�ru&vN�"CRٱQ��C�����QbM�-Ȳ�<�-^-��׾z��JӉ聢���cq~�~[jƴ=g�QA����D8�'���ٔ��5Q���5��N	)����8�1:L�P�]/xu������Z ���ѿ�_e�m�!<#C(`0��Y�����V#GYt{U�+�+�{\��ێX��(���u��*7~�.D���UX��-\0�]Û'~���k�e@ߛd�rf�/�5�a�"��Y��&xR6:1����&{��X.U��⩐�੏�b��7ow���"y��ʝ���ˮ�D�!�&����=g������d��������kcty>Y�Z�A����ȔT�_rA�%���{�2���B)epk_J��O��qɆ������oW6 �Iq|��t碗�3Hv'���{�z��D���������!�uY5�%�33��o��<8�v��kݵ����i�;̢@r�g[`����x=,S2���Z���nE4�V���:_��G�����BՆ�m/b�F�bJ�R<�כ�P/�υ�&�\#VE9���+�ZE8Ɠ�i]zw2�$9՗4���Xf-��$��~\�^R���4�&�N>47m���D����/6:�_̈"T(��XA:P\T�SeO����%�q���^�-����uo����or�`M��'J���#�%?6�~dS#�cW�}}��ަ��qF�H����!�Πּ`�
s�L�Ujy=�s��F�)�Aru@)��&34�����wOH
�k�AOA�Ӗ��n��4J��Gm4�Š�b��H�����QJ�0�S�*q�ޛ��������Oū�58}�|%����W��~�l�G~�VX��
UᣙOb���ǚ�):�!��y�p���"z�%�V�������Y7e�e�L��adGxB�O����u�M��� ���A֐�q�$����хA	��țj��x�J֣ʊզ94���!y�%��$�G��[�i�(J���i�3�u�]�.�t|DU���c^�Lë��DW��q5Bg�2�挢��j+V����ꋻ39��Rϸ��w��׌y�œ�'�en����Yd�PlV�v�3�5oi����,�MJ���;��0�.�}1��L�4ں��E2I)z<����_�G�Ob��@۷�.��IV�����nsJ��_��)��{�K~О�+j�Ľ������F�8t_aa,0�4���b�lñ^�l/�v�X\Į��Ԛ����Q��U5�x��7�{�59�_�{7�b��CFV�
�8��LX0�*�O��u:)5ꉠц�U��B"oݫ�z��Bo�$MX����zn��u���f]�'3�s��;}��H@���F������ڕ|�&Hp�$j����\:�����@b>{����eBטˤ62�2�
ʎ+�F,`�V���N���k��D�6 �gXY�U�O����ٚcO���H���>�i���g�t������u�l��#�*Ņ�e�B�����FS���%�A�;��u���@�ll��c�Z��3'���8BD!�Ǩȓ[ꃋD@��pW@� D�pwd7��>�`�wp+M����E���vj��>��Z�����30j=u�գM�a{<�ҟ�9R{����K���~�"<b/9ޯ�\%�%'(x���_P���t��b�"��l�0^��z�D�6�z��F��[�m�f7����zdN��J�:�5#���p��9ҥV� �*K�U@�ظ�HQ�1cO7�N��ƛ4�c�HA�l��ۏ����F�.N��ץ��i�?�ɋ���,�M���}�b�XU�D�y�{�7"2D��� ��ᮝ����@j-[5]{�ą��k�GM����Ή��'�6<��~m>$%�~�)IM���%�@
�#�.>1�.o�ˇH��)C�����u������S�+�R�k3!�Q7�4���?���v�M���� ͱ�W��Zi�Zy�#G$̹���_دӕ�7�0����w�<B*s�
r4 �ۼ\qq�/���,:|�oӍ\���)�,�~n-�ܟQ{�;G�Z�����y��&帉����Gq�W!�}{�|�zӛ7�d)i�w�9�~��1|��/��3g�)�!k���C�N�|'|�&��ͅ(3햄M�l�B:l��؄�xѠ�\��$A���<��%|P{�[��4��!Kc�wz�X��P�������Bi��nз�2]������o�~6'��nX��Wܝ��ř^>�X7��9��!�w��+�i����xi�7 -���6�1|>� Y���!F��݂��p�T���f!�*�2�j!��2 ��k�R���������ȧym�o^9���ۇ1��
��5��v��#9�o.�wE�i�-1t�eM�����DC��� �IMKS���Ǒ�/5�ب��"�q����M����:�F޺���E��F�f�v�*d�a:yZ �,���';;�>�2Qg2e�T}U�[BB���Y7$���צ���޴��u�� ҙ���ѵ��a�d#�MY��n�&V4]�z�j{�+,��pOr�R]d�9�3�
��WnX��؇�"�)�>�6�je���Z`1�@�*H�5��w������m��E"���u�,bj8�����`�P�p��Y��VQ��?7z��hs���p>�Ǧ~���y�E�vW����B�&lXY|���}���c�5�{P��OO� Cvrz5�������/#s5n��Z��Y�����F����-��0�]p�8���������
�U�.5��A�Y� �9�����w?O��(��`�����%��l��r�l��s�8�R�-��<��PT���fc�6�^>��[/��چk�҃�v�`q�|���o/�����k֥�U���O,sBg�+�B�1f8��v^ze�<>�z�����H�8�O���K��q��X��gQL}k��	����9�O<K�x�u�K �:�[�I*�y8��0֨=DX4���K��{���?iK#�Si4��I�@)�]mU��q-���]����$Jp��׃�s�4�'�����RI�ᯑ��W�Sj1��ۺ�xDX`�O4m�ˀ4{>x;]'�ZJ �>���������"��۝�7dɡ���F�!��`�pN�V��E͉�����H�[����%�#8���.��^픾3�-�
Y�7�A��`�Ѕ��Y3cGc�ϧ���u�4x���3�U3��� ��l�(v��5��: �v��J�����ׅ����4�Sm&F}z@�7�|���M���[뀜����p]���Y�W�E��T@j^D/�A#yvX�������]�F�&��*�->�@ޯ���Z�d�>%�C��A������%K���T�1y����eg �KW�2?���|[c=��YJp�B n�k�^�<_�bY�b�]Z����Rz~:0X�r����I0N1/|�5s��\�;�T��+ ���',�mw��_��T)�
{.Vd.���#����G�7��'��U4�2}F����nyH� �D��t�O�Ij��k���7�	��|tT�C/����G������QJ3�g��{��]@>�^� �$�O��	o;��<�0R�q��'L���gj�U��K�n�5��ܐ�ى�G�1h����3���S����j~���_\|�qm�
JQrXJ�m?�Y~휤uԍ��ֈ�w<�N����q��vɦ J�cjQ�o�ciң�w�~[y�]���}G����r�v��
�/r���n�t� ,)˓aʝ�2Ѿ�~��!�=��J��`M�O���xlQ�*@�����"+���K�^6��ٓ��i	.��m��մ�tMz[�߇�Pa��m&�e�}���}�"'_k�����T�L!����`����]� A�����%��Z�<>K�O9��.r�t�j1�+쎎6�,���|gԴalU�(�'ٌ�p��`�k;W6ӽ�C��q ����N�A2*��(�:[���t~��Nq��Q�ӧy��O������~^�[�v|�@��$n��N�Xd�vvW�d\9f/&�N��M/�Y+,��px�a�q���8'��-I��~#����`�7�����_S�=�,c��]T�W+���jޜj�o�a�B�k|6�k��]ڕ����Zބ�P�����:K�p�L(:�r��4,����C��:�2nZ��П���q�c�r�ƽӒ8~�ߔ��|���0�s��u���T&�'@�W�k��_l~�)3��p�O`�� �����ZA�� ��%Q~N���z�܏�b*���q� ?%�#H�ߟ�ؕV	߆�F;�%��!R[/t�i��T��^�;B��X<�Wm?	)�<I�@Ew0�w�>�1�o��0bs=�ޚ+�k���������a����!��8�ud��q[���v��Y����Z"�r��Y:�
��~��͏���2�@p���ߟN��:�'�W`)�Q�.y���{�=Y�p��o^�:�]1����ӂf"
R��6�6��.f��v��G[�0Q{�N'fr"R,-��s���IN�n��+{s]�	7�q����\Q��4�g4���Q��äX�����;f��搩��Nd��ك��Ҕ~��f�+'�	�����f:[O�)I^��=�>^�':ې7;�li��n��25d�X��h�^ɀc��7�yUe ��sU�>��������b��=�Z�D{W$4FT/n���t���ţ��c��v���|5���S��L_�x��5v�������|�%�HTr� 񌫎�s�,O�Y;��R4Ua��S�p4���_���øx&����N��45���b���Ig܂��� {���������4��#��w�,����Dz��r �9���C��ƽ��]:�g�Z5���6B���6���s��G�����X*�&� 3�;��W��Iv?�sط-��x����v��ה6J�I D�s���|W�~x`�	J���݌��i�-���V<Ałb�[�Z�ۿ�r;vk�@���(���҈�H��?��q5���/�e���SX�s,SQ���V�mI���H5�pE��;Ir�����yP0}�c,�64]��35x�H�F� )McS�*E�ʙ�	�C�+�j�+�˙!��f��0�?��>�#��s˘T��������,�ي�@h�W�V��y�U��M��g�iw�^��t�-T��oP`#u��46��g;��a�c:��Y�����#�-����;��k�����F�����3=cd�uŤ�N�nr��H��ߪY���΀�,ȅ)�X��D%Y%g�� N>�5�,�T���d�X�$FQ��%1�H��,l��SP>S���l��W�����VK�D�5�٦`��j�|��	������D��R�k��M�6)i���ρ�)bp�$�g<�"�k�S���=�ԅ��Y�&;z7���䤶$������",��1�1׃���%F����0�?�,���ˇ);h�|�e��Η�v�qU�Br8C��u5`8�1284s��w'R�5|�������X�U�hXL���0��T�R̊iQݏo�Jm�9
�"����v���|�n�"Hi�h���"��� ���m����3���%�V#�4��j�-���f<���-c O7`m���@^6��}�,Qx����36oq���,'mO#_�MZO)���;�.�Ef��t�8x�sj�#y=V�e�uFl��=�i���K4b�)&LG���S�=G�5R���zd����L��� XW�A�ً��ta�]<��;cNXSH;��3���p�O�Uf�ޘzu�-N���H�G:���H���'�<��J�L?�*�l@���|mtIWk�5}+���s3�]I�a��]B3�%�}��S�0���_R^���-1���
��O�|'&} �7�Q�g�37��oY�?y��2�7�L��A˹4І��^?�m�%TxDׂ���sFZO}K��W��ə��m� ���:Y	7��;F�岭��p{�lC���RN������@BV�eU��@*�W�r�D��
�zJ�?za�xD]�*�^������8��:�)����/�]�P��FnQX���G���`�|�oo�i\���U��� 	v�~kW��U|������](S}��y�%�=�R�s*Y�t]����Rl*�<��˘����k�k4@�Ԋ��9��	!H�]��>��Y舵��Ѕ�݁$M��� -�n�x���Ύ�c�ʺ��۬�������(?�� Z�,���UMj����A�.��'�8"��(���sК�V���f��y�X��Nc���mZ*�>}k�
�`m�iD��q�g�����S2f��tlj�X���v����T�'Ɇ�Pȟ6��Z�?�l}PS��^DTD��tA�tE��NDJ�K�E�
H	���"B�Az	������w����?����}w�}��}ߜ�2���~�n̗y�܄��O�������Nc��y�966�W
�k3#��.2��>]y��^�<r8 ��܆��(A�p���S�����;�g�4m��a%1���W����C��UX��+�rA���F7v��a�t��Ԋ y�oϮj�8�\s��΅4_a���/��d�vlVy��Z+����Ƈ�f7e�6N���U7�d���-U���R��cE-�!�q���B�z��ix�xP'�ဎp�}�&W;�8ɌD߶���dz=�ݮ[�4?V�F�RѬ�3�_�=�'Q���n1�I���^��8Z�D���m?9f+���<r���븮����U;��\�](�q����@T�����DH
Si���>W���.�S������|�y�5Y���9W���U��I��j����nO���6("L�z��������Y�㍘Q,�(`�-�#`64�+=��q
�m�zW"y�<DOW�uy�簡qǵ��W/vTVm6�{�R��J�u+=���J���[H���%�خ��?�~Mʋ�ݧar���B�Q]�zqwn�/t`����s��/�u�v��p�|J(�*z3U�*e�`b��(ҏ:�s�XW�^r'��l��֕p�l���i{��aj_>@�P��^F{�;$���ԔH�۞ސ�q�.�^���=����V�F���,Дc}/�c�=��դv�-y����]���׶_�ԗA| &J�w_�q��$4,<Rvd�Vep�:%*��t?\3���e�e��n���ݟ,�Xm�3�Y�>���3!0�:�(Aן�m���+�;4�S�a9��ܟ9k�U�7���,w�KJRe2�
�������͌�������Ɏ���Vm�W�M*�ҳ7�����ë7 뵴	Ѻ�p1�o����R17=��]�� �}�T����[�����/C�D���oc{h#'�,��y��⼖�q�V�4��["jR�����fG�����~c���{�l\�x��}Z��E<)˰�ofcV���7yKd�w@$��:F��)�SO��})��q�85�Th������v�r�N���5����GVW͝�L����`��1m�z��ѻ�����I=���������ɠg��7t����(��
\���� H�n-a�����1y��в��H>˥ؑ�)�+5�5P����`�}�]Z�	�[{q�+��z E{���xu�FAMt�i7�6�]�c����a��T�e�<��򣛣��y����qT�����Jfh@� x��<گE�D�M�6#Tt��E�����ͽ;��=rmr���O���|W�V��n��G��{:㇝��e�^�ʥKݾ�^�a{��W�drv��#�6ܿS�����1��u\��ӯ��P�e
t�$ ڞ�"hQN}Sq��ր�<^;�V�/g��ukP3���2��e���`R���8��U�]UX��W��qxM�`0�P���a`�T��T���z���Fs���JVQ��� �Q��G�f/�o��G��ɚ �)���'��_^k��V�f�cB"�a�B���;�0���t3� �p��yM���j�cv�R���>�s������t�׶�Ӕ�'��I�1O�n���3a)ޝj�����<�UK숎��ƭ�ژ��*_+�X4��$�S\5��n~�����]{��p�&�"K�K��NGm���+��I�M���"���F�j� eX���c�'�,�:5/��_V�U'U�߄��j�x �+r�2���P��0y:K�J���h�<��F��.��Z]q%�
\;;n��N/��Q+��鱠��}� ɬ9f�i���C���0���q��j��|NV�	�@�ߋ:�����χ�;P*�)H�f�l�S;TB-�\�׼�mTN-�����pB �������� ѭ��7����h��C��5�KI[AW��_Q�+��n���9j�5l������4���?��Ν������U�]��P��b7��ӟ���j�.�S�6˺��o�k�%�A�|�f@(|E%]�	�=M�~@�Dň����N���z�8�TU�k�b����w=�5ɺ:�P�1���!"��c�TD(��o3� /=^���l����ء���S��~��Tw�ӰU=�.!����5�LY����w����畩\�m�a���Mۼ�[
Ҟy��C�69�36�	A�oҭл���,�讐�N��w�k��J��9�������U?�zJ��Q��q7uw�A�
goWn���ׂ��p��ݦ��������(�Z;to�;a�ʩKV��B���l�҇��WQ������.u���W��1�����������CJݓ�n�uk8 �v&��~��^�	�����B��d�յ>����'���F�U|GQ�k)�9�0D��Ap�aJ*���0�d�+�L�p���9�L�Nr��@��#U�����J��Ϯ��O�Z�9��_ i� �ú���@��+�� ��w�&������Ε��oNV���tu��MN&����֐&Zg?ŏ�����n��z=sv�n[��w�l��U�?	�[�*���$��̑�Z�Tj��3"�X��O���	�5^����S!�O,O�R�]�!�rJ ��8�e�8�����O�}�w���$��=9_;�L��AE��uc�]����`��a�dI�H�;��Qz�W�j�Ӆ�d��
�X�r�}���CQ��Zr?}k�G�*����,?_�8!9�~u\���=�{��b�#¼p6LJ�n�~�t�Ȝ�UJ���JgU�H����e|���.>���T;�6�+���ά5�MQˮ�:����k��3j��B4����Ͻ�M^�~%�X��XJ�27�*�!�s�r|S��uՋl��[�y:\�{ZJV	ykq�2�1K����Ra?�hH91%Nư�g4U�ŷ�]u5�Q�~��>�����?[�a�ۦ^��k�dhs�p����ۢ�-��M
���7��C_A�Mℷ~�g-D)D[V^(b�'d��C?ܠ����˸:}�_�k��`K�;��X�+"�>������{����t�]��u�28YŪ�;��٤@��K�]�ߐi|�}v�g��{-NR�\b�,6�Z�$y2�EZ�8$Y�Z�و�N��4V�PL��*��WhBY�W���G�$��1z�G�8M!쩾��-�a5br�7�S�]Yg��A�+B'^�6�걗$:Yn�+�ӻ�$��pn� ��K�A3����繍���T��|\��fG,vB�g�HѭE1�	��N��1 :�}���c�����_o�Z�j��~� 7"o9�:�`���y���	|���_�n$�n3��}>8	�v�^�L�X�:�/��O��v�nmG��;�� V,l/�]��h�d�e���)�5!�>���J��g���9�D�������!�b�K�5��;���8�{�����c߇$�˵��.����0 �abq��s���b�m�����\�HЂrcv�V�n�H9D.�a�i���{<v�Uډ�56�E�މ�)c������uj�-B+��!��������&r�8��Y�&�~o�M>}�I�#JX<�%ɏ�?�F�ʍ�c:���������� v"C��T�M'�-�>a���v����*��&���!:�GM�ySܟ$w/q��p�6`u�0����$�ڼ�y|x��B"���E(�1rg���Kn���� lv%z��(b$�+�gz�������*��EI͋�g�	�zȼ��ެq�	�v��$��j���_�]*ڽ�ˈ]�*xU���Zs�!�y����:�x7I��oǠ��F�#`�R#�*��8dT{�B�9p�nLĦOҽC��f^P��C�D����Ta�n�w���wS��]zq�>g�qM?�nU�Lb��$]\�,�P+7p-r�*mc�V�qr�Jf�.���y�b�?Cud�����w�Z�s��;5�V���:���7�n��,j�c�w�e���[_�ؘ�"�*/��2��}��O�_��ue���tp�+O_pǿO1�A8B�$8��k���|�3n�B^Y��w{���J	)��o��.V��(HC'r��~�y�GS���Kߝy�&��7R����=�T �Q-�.uҩh�!�x�k������5.�Y�b �c����C��9�j^ɧG�~i��S��'y<M�9���"/>�"Z�zL�A��~=L�}!�WzHǁ�ς�~�� �OP5���<[����k���^�i����T-z�U )޹�����g�蔗��[�&��MOc)�mp����c�Ivi�cC�ڍT���'T<wܫ^�	SQ@S���P��`g�r�� �8H,���U��J�E�v�!#�������	۔T�P��+�*���(�_���kk��f��UB���hzW:�S�`M����V���@[�Ȳ��	@���x鈦����G"x=�l�q����%�8�"���c6�|��Z9-o���ڡ{OMZO��4	�L���	�Ƚ���ƵԶw`ѿb�w��
�@�W;K����%;�_��� �k�QNA���[R ^�J�哧zj�nA�~��������+\�a���WQk����xꌅ3)8}R�ILs���|ڡx����+�U��<9�#�lS	���Π��'�Q����x
����3~�x���Y9'�&U��A�>�N���VC�65�$�ֹ���%C��g}\�Ml��?8�TX'�f��|A�<��?O��G���;z����4C�SV>$�޴�Z��4�]���}�؛G����D	�BA�� R�a��ܓsA���NKWЄ���2mH�V���_g��um���Ĳ��Ϟ��1~o	�@�
|�N��F���P%��#l��q���	��X���ߊ�&Nk�����������)�SS`�"�'�Y^8�Ϟ���5y�������g4.�����o@����r����Q�f�\���'S�Y�YT��7�>���S�������'�`�o�I���NK��)U�s��;�y�`�@�����[��^����������Q��j�R���vI�]�<8�W��W�ݧ�_���=�,\c�1�q��:}�v���sCB�p�v�]H͡���ہWw��&9�{�i�k��¤f?�	oL��^u�»Q�n W�E2��u�����\�S����>�:����|-��]Xm�H�-�*�!줌AbS	/)?�������\�!�(}fI�(u�_.ڬv~��R)j�H��Y�d_�f�q�(<L��{�y���*V^@��,�'���e�2ﺠf�h�N���{3tk�pf�%� ����=�_�v|�S��˹	'��o7�?��/K���N�@{[Wm�}z�3��=�ҿ>���CH���M�N$�ΩY���W�J2(ϓف�MN�[o4�������iX�uqs&5_�B9��-5��'o��#���M���~]��ﰓ?������P�4 ���$���ө�Z��F�LI۠��E�PX������.��Zo��q�0��ζ,�e�^����Ճ3��>��Kq�?��/J]����;�nI��"Q���?����T�������W�@C8f�=*#������a��� !4��c�N8oE��I�x����9 Šwɰz��\!�U}���8ɄYy�����.){�yej�a�i�L�4�]�a�=�2��0���P�}y�v2FK�u���[,{9���̈́ەo� ��G�nƓ*U�ï����.SD�k�a����z�]�D�Y�X��87E7�g�R[�K�H�(u��r�]*��='JO�����mI�m+5�W4c-��h�F�9e��d^Aѣ�2�x�5��܌�e�/V!�0w�Ot�>����G�t�=�4|�N�֤b�� �����{�x�<1�=��Y_1:������u�G�f�`3Ъ!2H���I�&�� 1��֐�ת��h�z�R-�6���|p]��HV&��{��W����.���L���v�A����V��5g������bZ�M|oh��A}&Ng`T
J��Z���&���[��Pi�>�px?ql�@*b�]5�;y�M�T�-����~}�8Ģ��ȡ�ϝ������h���vL~���8$����
�]��IN��@ߍ��

I@���^]����MDef�';m/N4a��WB��QE�ZW�� f�����QT1B��Ewx��:㥛xk~�B=�eݷm�D�RP��E<:J�د��Q�ӽy�yw�Bp	�������vX렽;a�k��g/f꽲�|	��C�g\"�$�_ت��>Ceg��P��ɠ
w��;$�����>n� 9v����v�"q�EM���Z1�J�6������{�K�
,*!;a��:���2Ŋ]��tۡVb�,�
:�K��+4�52v�аqO��ۘC�Q{�ۼ�x�ٞn3�"��䬨h逥oo��g�3�W9��lhvL�}�3ҵƏ��I$;O#]�IF}u��ޥv%�p��(�u�ߑ>}��,҄���s�*���U�M⵹��{_��h�Sз�׺u�IV�E�Ďz�}'�<�,n��^7��Q-�&�`�qߪ���KKȟm�x�[,�"��`�����9���
[��n��嵁g�.�|���]�ߐgށ�N�����L��zj�����P����ӧ���E��L&!C�"G�XS�����&t�=����)|e	����w��
�{�_��r��+/�����\��nS�,k�O�4�u��]<�E4�cE%�a�%��P�66�C��Sh��[:��Dv!V��*c���1}I\������D٫ �c�����=@�������px|�d���sʞ�@c���u�s��&�~�4�.r�I��˱�%;uf����ϽǤ�2?D}�'�=�Ƶ���q"e"�~�����d�Y=��T�y�h�
�(�i?��[bq���>������3X(�vN�AV*���t�߇�x��(�u��_�ɣ��.�0=�W��Gbo*���\M�zK�����T�u�ׯ�d�u���ZW�.��Ѷ�SX��g��Yf+��t��r��f���u���{b$����A��m��&�A����s�tr85?����74�g͊�ji��#��Ch�V4�8��	�E�z��η�uT�4�m�g��rY�����4���~���`��A�;;��
�f��TuH"�#���F�@g��=��p�$e~��)!�����+il*6ʀ{����ʯl��i*�<5'$}_�?�&���F<�΢�]��h ��~�ʔG��%Y��#��I��+�R�ޚ�y��y��g�&�L�g�_O��I������'�֔1R��L���~��N�Μ{_:B4��-[����"'��U��.����6fx٢����܍&��5���rBw���ۮd�5��L�6�{wU{��ֵ�iP^~��9��{��V�G����u�ʿ�-��2<\��k]�Ї���Els|N��g=:Uڪ��k�b�r)�D�TP���5Ie�1���b[�<|3(\���.R�$�	<f����䒛7.��\}�;S:���fzgס�BZK�jd�w1�09��i7b�0���'����EN�g#D�ɋ�WQ�Q,s��*�+�����@��<�ȫ�;3}���|�h��
�[��$�x-pn<ԡ�Br�5�&8?%��>��5E���mb�|3�"�T�/_׶�|��~]��yҩr�UYB��_M�f b̰u�hQ��=�J�G�hر���ڻ�	�Ľ�:C��������J���3࿟�><�	p�:�NN>��T�dq[�!:a{W�I2u%�Z��{��8�c��VC����j����W�b�����Y�o������Ѐ�K�fU5Fʠ�&��~��G�-ƘD�f�+���\V1�-S�Y����GZ��Tc�L�Z񘯌Ij�W����r��컴��x��|jJrD7�H�P"���0d{�t��	���뿮��<6>:#�!hcg:�lӴ"!�l���`�׍/N�$�� A���w��J~d%1�<����-1V܅`�B�>�ȫ��2�7)���-����S���3m�ZlDu��fώ)����+]�_�筽�粁���⭛��K�TSy܇5�g��`�[��Un��� ��nV�ϪD6�tf���c�@�k�- b�^���{��հlY?�A��,�epw�s���WQ���}�=;5B�헛n���5<_�b�2V{�M�`ab�Ķ5̔ͼ�(��ҒY�b��6�W���t�	�!8��a��]�d��Y?$X�Ě��o~�a�eiu�����M�� ��QQ��W�o�z���t�:�^��H���s�j��ڰ�r��‪¬���ɃgyKNQZK�f��t���3�����훠f�r-�8�߼_<^�޶���֭ͪ �X��)�����ՙ���4�+�	K�����Cfݢl=瞦���:�	��=\X�E;���]c]���c�Q�|��Wηnj��7�)j�I
s)�xZ�c*.�Ӹ+g�
��&g��I��]�������
��QO������ʃ�O�:b��� ��b?fMN���9���QW;�����\KJ��Jc��L�~"�JY����ʗ�U,�k7�kϒ���xLc�B\�}�`Ӷ�a��:ɾ;���G
^�M���yl)<��Ĕ��;�ڀOŦL.9�t�M�m�/���]��.�,�0�V�^�GR|��C5V�D�
�-���P"8�S
r��{��\�D����w�/��\�2"e�v	(��h��YÂ���@��n��xB�Y"Ni� LuO߳a�-��Ѓ���ΊQf�*o7P��=��E, ���;,T25��H1�������o�І۵
r/�_��?����-Pj�ŏ�zݛ�zN��韜�˻��+&qה�C+��0\IF�T����@�0?Y�E�w�������x���]��)9~��kD%�=������㥛/�"�a�.Ԥ�REE�E�	3��tQ�|@4�@ൕj�/.���l$����b7�CV��U�}�&n}ٻ�Y�?�Də���N栾y�E�v 6鼤�3��t+]��[]c� ���-���݈�I����2:[HGK�_����f�1��:�r<�1�jӭ��2�� �g*�3/>��}Ě���"����P��M���<�@��?^6J���Qr6J��6��h�mP�؝�0vE�ɚ"�������F>XUR�jh�����%�Ϥ��]��n��,R�43�����@%C�Dz]!$ R���H�g�����TJ�ՃMd�כm[9{��*�5d�@ng�}��Ȓ�ƙ��wfX4��o��<�h;����/U^'���o>�GC	��b��ސ퐢�e�m�BO��,�\YTa�ߧ��� ���s`�����1��t��Կ�h�}eY�Q�} J��f����a��+�n,SVz�����	�A����ns)���5��X�x)A��4	���ɲ�Sқ����:���T�q�q�����X�l�'�cL�Q��~�cުɐub:�:�YD���@�	�M>����y{}�L��h��!��Z��Ħ&e�7�����u���{�П� �V�zO{Y?2GD�^�j��P���/��L�Lл1���(�Kv��+=�)su'�in抆O��&�e����
h�Ŗ_����/9[�y8L��.�Cv��Z��6�R�ݑ��fr��%F],In��Rg�<���C�l
�рK^��=�Wc}H�r`�A[+5���ҿ�猴&ƺ=�Iq�]����<9�Ѫ�b���J�-�I560�a�LP������mC���l�y�[��tJ� �Tb�	r��ܳt�
��@��y@�C��	2[�.�W5��.��uW�L�E�ǐ���1w=f��5ݧp��<�v����<�e�YeY��]7��p�G�~O�<��aiLQ�&.wx��Y�Bx 1���a���ߠ�����$��w).�E���n��5�'��Ѥ��Ay���m{�U5\R�Y���������� P����26R'B��g1�5ٚ�3h#2T��j�Y�.��>>QI6+�
%��E��P����T�\
L��i�2�p	9�������O���*�F%4�	�:�)��w�vo�~�Z�V|�{K�Z2J���K�߄��h\��Eb��_�+�S��Z��%�G�k�aa�iiMCOO�5��Mk�F�Sҿ˕taK��i�;�q�����$��dq[(����/fL���Ո�p]iϒ�ՠ��]��R
��#��OA=G��N!���%��>I�y����{�H�Qu�f�6��H���	[�a9�8&=8�?O*D���d���C��J@�rHSy����Z�X��Ե9��|9�%"�d�ޯ�!�L�'�qg���V���Rԥs�a)xyd��U�O��b���~Ȍ��4"I>| 4�dof՚��e����wl�Cß�d�K�_��M��^:9��t3μ��"���f�˭�>���MF�ɒL�w�$�9wt_�f��(�m x���J@r����>h�"��V���E-5�����B��Me�����4< ���F�%J�+�+��o��M�˗I��5f1R�/ ���c�:��@	h����r�K����
��Z����`=�YkT��pޱ9 A�!�@�:��_�x�4��f��؁P ��VRB��T�ҿ.�#y�ɔu�?&�J7ui�'Kϼ�T�z�P�O��ڮ�@|�Q`�Z9k�@�᧝Ǚ2x�6Wvͭ����
,˖mf� �a.�r���{�M�f�&1�����;w%Ō\�х�2�w�XI�Y�Ѡ�g#Wz@��ҍ�w��c�7�@d�.�����Ql�C�z�s�pH�k���2W�'���R��\��h�/��<?H�S���Y:[DU�Ī?-����|�?}愦,j偅�Lƚ<��C�-
dQw�-z�Ai��Z[ĘǨ#��څ>����u���M���*�@���[��֏r�~�~������F4�_�QBgR�e�a���_b��Wa��A��U���]�׎6Z��-D�C�4��B�؁��~�����t�s�BKZ@X��ݪ	a}�(ҫ��,��G��3��NOᏣXF���F2��Z����}�b��I�\��C���I�'���A��+&����K��2�����u w�k77��yC��!sjvO�1�H#0E�q�k��s�隴����kr�4e�+�5#9�骬L|t���F�g�%���	�Ǥ��uv�v���8��I7�r�8��w[\�K�:�,w}����X��5�/;���H���q5���{BC{�"����{��T��g��,�q�J�fl��r(������j^�3��_�自��y+f9�.����,З,�[�u:1K~7zA�sw��-�tyqDCٮ��,����7~��XC��߮���]��+��X��R��ڜ�H��{ct��}X�c�ʍ�k����;��'3	��ip� ē�Ղՙ��w����}��b�*������
#"����Lʰ;�*Y:�f�, WiU"�%�e!��ym')�g���h�p�~�.�iq���?����#󘶥z�e�Wԡ��@KL��\��%Ft|��f5l0#��f"PZ�6iz�u�bXA����f�P� "^��	B<��=�e�1#d����1�+�e@e�gi_Ŝ�7K����K��r���H�u�M�����Ӝ����0�;"d4+�����|6��p���j\���s�o�ݗF��u�)�l&G���e7���G�N|,ss��x[��2@�%��±Bv7���ᓤ��B��"�''wÌ�N"mg�]Z$�`}���K�R�.�;jY���FmK�x��Y_��R�� isBs3o��=1�%���:~�Q)g\����_so�O@�F���6�gLp�-f�l7ǧ����^����m"�hW���H�_��D���zx���QhW��8������1��0 P\�qA��#r�^����N�Q~fhe7�.M�y�z����0Gu����A������7��D�y4��R�=S�O�wh�2�~���W"�S$�G�AҜg
�-�:�y�[I���޻V}�'S�Ҙ-s�^��VX`��!�2��������YW1y*�k��k*|h�5�?&J(��tp��)�U�ߡ/�|�d�42��V�9���?>��]��*t0�S@]'f��4�>	�	A�G[�Y�$��sp�<t}�7�'�-6eq[�,�0z�Q5֠�.�;g_����J����4-oI�h��!�G�}���a����`N�X�������gPb�m8#�L��̧��?R�f����p��U�z�i��FO]0��BΙ�тТ�2����7I/�5��%}A�y��`G�����]w����Ɓ?��\�_��Tʾ��v�u����n��B7�	6�2P�-=xq����u���z��0�G�<�������~ѐ,s2��^�Ru��=����nK�k����N��gn���*ع����@�b�.���������DJ���K��vwK=W�(��i������Mo-�(��:��|�#�t�~u'�Sj���e��|��kCd���I&�l�ݢ^��<��z�X!���n ����Ud'�q,��ʩ�K����;Ȱ����5q�M�<2�5#���q������@�)ya~g������/}�� ��o����f5��[z�
�'���ϼ���f�[?���������o�c����K?�XX��j��4���y^}�(���;�@!���R��ތͥk��H�|�q[�|V����PYG�j�P��{/}�:�dJܾ��,pu��2����)&Θ$쩅��5r�V���j��ߠ�O�X�pB��7���%`W�p�����OC���5��gU�k�.�Sl��J���i�6��eY#�d�קI��������Ė�F���i�����,�����jr�I��i��M_KxF��{�^LįeoQ��*ݹ�l��,����
�����(�K�A���h<h���|�sj2�T����J-�Ƚ2�	������K��]���� *�:��߸ֳ1/� cU�����:���G��������Ew��Y3Z�����,��2����VVC'�t����IKĴ/ꍋˢR�C�u��2�71�l�׃ĪR�qf����G���͙�O���=(�ͼ�>@���w-��"�c�u�4x��t$��0S���uod�Bk��C��#�oAr׽A�*����3n70�e�˂�5�&)��fXc?� ~u�iܙ�SZV���oz�N����q�߂���h����W;ӑ����,�+�i5�K�"F>��x��n��R2��_(6?��E$�t�$�?s;�P��-Q"��
��*�Z�#����h�@^1��9ܧP�f61��&�~��o�}�·y�h<���)�J ��|�
��<��=Id���T�� �k�C�<yq����V_R`'=Vz#Ѡ�Jby���k��ýy��J7���CO�%\26^║I&N��;���v�8B�?�jY�9a~����F:���Bx:_����}�fĸd�ȟ&�c��wĵ\ț��s�k��`
T�e�ｓ���g7����͝
���u�N7q!�1���t��f���6�y�-z�2�N`Nk�, #����yJZ���d���W�2�&�@�:�hi���ᑭ��&3��7'K�����'�G�3aA?p@��q����i�:7�'�ȴ@��q�,6\ �m��-��:�E5����u�z�Ie�ڢTd(���;t���o}O���g��s�<��[�����ok�Ɍ��M�ʳ� 4GA4���E�Uە��ߟL�R(�됭���fL������z��N|T�{0b.�'����C����ү�q�E�}�cS���6�I�<��6��.�"*��r�x�\��/HL������0���������e�Dޅ@�&bl?Q �D�������@��O�L�g�Y��K�z}�+�.c2K�4��F1y��/�+!����o�D
�X�!�P��z�bJiO�!�&��&g����T������̟�&��-�q�h�	ݠ����j�ĉGK���ף�A�t�ϔ�^����;=�]
/w@��}���Օ��޵����P7��5�8�˅$g�N�h�p�G�.D��	������D�P�>��i��b�긭��L�2��;�J�b����P����?F7ìS=�٣�W�Tp�I�z��ړ��4zv�-���21(��~�Y�p`���4{
�V �V�<�����aV�?�y6�P�*�"$|�sE�m�2��0�78�7ų���_��#`��Jή�,�-(����=3Y�䥲Y��j��O�M�R(��"���/�c�坺8eE@L��Uڿ:�'CU�x��չJ��y<�Ǹ~f�8�ul�Lvx��E@�����'��O�l�_�����8�;�=8A$4|n<���"�@�;��|��3/R@��Bw��3Ě����L�6x �$�]�����X��}g������»�8���㙩鷯��+N5�:�Np��	�;t%�-�/?H7��i�W��Z��H�����c�c��#�)�Ⱥ���a�+�E�����p��@���Z�����(���t�N�n>��Y��S7�4u�`�TV�7��� ���_$�՟��fL�*|�"��ֿ�Җ�Z�T�������?Ś�f����i��(��PU5'A:#����'t�7����;�L髱�M�2�uJU��ܝq8� ���U�͚��q�E^��Jէ� �/�����C�,�2�;�0��X��Z�,&Y�6�� ������4����9`ҹ&���=���v��'���|	������f�]�xg�6d}&������]�s���l6�ڪ�G=�|C�¹����ڬh��f7Jh�PO�9�ػ��L�KXR5����G/<�>�94����{+�.V�8��V����߯���{q=����Zueoo�$�v�h]����b���	E��]MЎ0��3~��\���������7��<��}�����FG��2��F�j{����T�}�fJ��c��籲���rSօ�4�F[�]� ��:^X�Ӓ7և֎���ʵ�w���b��r%�^Vk�[t�O��F�{|��'��6j���u���y矿Rg�	�I�3��`��~���5u(P���.���;������?�?x>����:mc=R�Q�e@��mpġ
e����f�'�hRn�<[%�FQx`U�ɩV��R�뽗�&O�%�4�[g;��^���)d��3F����*�+���,9���v����	���G���Y]0g�j���8�d~����F����������Ҋh�>��}��f[g���<J��0u=���O�|g�F�������w��̺��q�G튄�e�|c[�Yx���e���� ��3r����L���#�Þ@��ЅZ�?�U熫��Pi7Y���i�i
� O8QMF/��[����=�w4rX��~�A�J	}6h�gk񣡍����#]G���������G��I��� �y�W��]�u)��&)��;���Be�h�$QǠ���h2ߖL��*��/����L�p�Ef��(��Q�,�r�Y\�^�q�]]!R�w5��F��$�=�n�d�����&@��	m����#g��t�+�^�?5�#�[�3������=�6�s��L@��eq}0��RQ�5������@$I��S�����C�PB�.���E��ė2�q�������6���E}�NE���Y
!HO�n�$N{X��`z��^=X�tR֘f�Sҿ�b�|aB�L"�W.Cd��SQ���ӛ��
��՚6������1�DE5��9�@ZtrY#v�f7e�Y���xN�ݗ�¶�rW$��8�r������Ӻ���.�T��XuU�"��9�ww��S��P���~�T�� ��g�'��ӯ�M��C)�2�G�S�u��1]��TB*+h�4��X21�S���=�Fޗ�ٯ&����(���� �J�7^�>r�*�;ڹ�u��k�n8+���fg�p�ya��� ��]�����:2�
%�=גW̶��i�~��K���h��h���kM������^���e� ��)��/����[���T
Q}fa�zKeC����i���ɧۃG7Ÿ�
��W��?�곣�i~H��υ@��-!a����v�ĦN뽂�S�v� ���&�Mq�� mUV��?�UX��g����?�`����l̋��!�w���2�A�^��h�/�,��P��Y�#�]�k�7 �����7�{�l��শ�3 T�x%p�3	0���2�����gE�����nE�"���G�%�M%:o��:��D��v�Jvߺ^��m�X�o$��2��H�
\�\�2�-a�O�09��)�}�Lp�4��M+�iB��-dt�G=��z��+��0��7���5	�A�:���ve.�UҸ����a��}�N������o�m�:��7Φ���}���~��ȨQ,/��&=z��������s��V-V���O��'D��q�c����ɳ� q}�d��U��p2�+�_8���{��`�^s̺�dm{ܶ%ڡ4������WW�E	��g������M���6ㅨ�Bu��Ҕzn�{�q�U'�f|�F��J����ǘ)�+d~�=m��#�� Z"�T2�"�'�ׯ�`<5ItRj�R�G�}�'�s��O]cs_P�0���rq���~��EZ���J���'����-ښ����r!�V
�8~��)F!�J�6Ʃ�� ���M���zo��lx�U� ��x3ӵ{������U'������گfk�Z_�oՍ	��h�;#�c�K��f��Q�PM�����RI��F@�EJ�D�ADJ��K@I	�n-��%'Lr�Fm���������Y=�9�u���z��;v;�����ϕL+ߋM��f$�}������+�=��l9t*����w��F�ɼT�l6V7����^7�(U7��s�/���+6�ӷ���a%�нf*���ȯ�??�]����|��s=��u2����)�	�Z�"j�:ju�f�
�g
@��Mnt'2zg�6�x�M�KN�p?4��n�e��:�b9E���E��_����gk��hK��'�u_��%���T�War���IfB�}b'"p=B��sv��+������N�|欈����>=��|m��"��Z��a?��ud�ǐs]�������.��S`>��`�[ �o��zS �I�w�R84t��*����5�U��k�,�2�B�p���]\�ㆸ��a/��|�Af1[�*��d.�$�]C��5� ��Ŧ�@P���l|�qڣ{��]i��-�kd�r:��V��mLʄ��L��-�$����3�/�Aŋ���f��$��B_��W���1�"�Y1.d�VeS��,�2p��S�����{�Z�A�m?{��Ѹ�>40[m��s&�"3����M�ϒ=[Gy��3�����v�O�R��>WVp�dW�:���**�{tSV��XMm-yF����c��%�"�`��4�J�S$U*.��1�7)�(�*��Cn,P�ao2�	�1�ު�����T�N����Ą��0^b��������rT\�Z]o��b�v�ZqIT�,����?�:�,��h��o�Cyv�M�
]��jQ1m4�ƜH�x�'�	�]F݋���K�T�Fӓ9F�f�$����Tb�*|f�d(�Њ>�3���#�B�,T����dO���w�'X�\�p�������q"7R O8�0k',Jg��玃���]���T�7}Ҽu�rl�c&���:U0P��ܦ0�aR�D�ξ�n��C_M�A%Cw�����V$������_�#�}�T\
R9�1��^tD��m��m�����=��vC�~W3�<~��M68�~�p���4���]��zoZ�$��~��v�D��&>`Uu@�^ �R���'�J�'jv4=<���Vc�r>��/PB*4�-E��Z�Q�]��w�k#ʢ�Z��c>��H�ң�-W��*�0�=w�������s�4֎��F���y/M�5���P巓�V�ڶ��i��=���&o��jR�L̀����`!�_�֌�RM��QO��Ö�[V&;�653
�������驘3M*���ԍ���O,���G#�/��
�ØK�fየBz�/t��ն�x�&2��9��Re�h��+b�L�h��>&M A�#K����n��\I�y>��e�*��b"-v�!��'�`����I�5�o���v�ME�rQɕ*�õ9p�����]�|��!�_����|E��{���Q���i#�H]p����L� {�ʺ*m6��CXᗍ�u����H�!A霮���~��&]�.���da(�\�4.H�m�' �����-���٣�)m R_-��R�H�l�ܳ>!��:r�n�yē��8���jb:�o�����������(؜�w1x}��s�5w���O~Ձ;E�LӮ�A�	vӖe�#\���\b�g�����Z�B�BH==�z�Ms��޵��>���	��}�l���ʲ�'#+/dv�`�fgG?��~��\�F�.5��J�3|*1���t����	d:;)�+.�mMm�;�/K����=���{v��*3sT�CsQB-�w���q�g���2Iz�%z���j�f��Y1�u/�� ��$��.�_��86�X�{��.�fΕ3;�֦��	`[s�̋�Vx?�)t{����8�����Z��ڃ�h��~�:92���@���@�����շڪ�Wm��6�g�%2-o�iN�[emr8s�EZ��[��z�|'�0�]�jk�\AZ��6K_�]���Pl	6���R��R}[d-��<��2V}���ųF츠S*��]jw����[wO�8��7�A����&�f�x����OO�3�#t�&��~�S�^s;���Ҫz||t������Y����
�e*����6t[�J�����,$�Z�L����m}�bl�Ja�`+��e��c�+�Y#/i�Ϩ���Ȯ����,H���76I�����zZ�|/��ǋ�_z��uB���_�"�wH�~6�ӱ�����C��uD� ���w�篚�y�'`�/K�����UHr�l�%�]����ICC�]7�S|��`|������Z�5�������G�ϳ)5S^K���tQ�����%PO����'��V��ԭ<5M���c��Ϝ��ɫw���B�o6C\�%jqȚ��}r�BLYE��չ�PF�� �ƲM�r�~�u/����x�3��P��f3��������@[���B�,�"�=y�/��	(��7�i����� ��1v��d ������%y��9Tc�?�o��\ʀ���x��z-&���,:�t<U���t��g��� E,�	�V�!+Qѳ!��S�H��|� Y�ݏF�2���y����=O�u�������u�'g��Ik���B��'��'��4���O�Ȯ��&��"����ֺ%\�2(��G`���nQ'9w����O����C�N���.�Ϯl]�0���&Q��kwl�ޝ�VT�%�˺�!'Q
h=�T��f�#}4�t���G�u+7x���P6�
�&#eZL�=-��|t����r��!J�rm`%<�{�!�Z3yalA(-V�t��c�#*�|�Gx:����zi:e���a^���Rgw��)U|�8HX�"֞{������
 "h���������=��R�RV�����#�M#Z��ڧ���^XP-�U�(��dΊ!�p������=��^{�3��.��77oq� 
���[�m��c��8��:�#�L2~��\��:��%\��>-��1���Y��p�Iq���Dt�FYU�~W�!�c@�)h�2þ���R8(ڜo�i�Y���\��fǸ�w��d�=��`�<M%~j��(�|��9��YT�Q�<)9^�����:l�������>��ܸÿZK1�/�MD�n����-�<�FC5]��u�g��-pz��ѩ�@����F��{��-p0�����E���5&�n`<>�[r-�/��&���ı*f}/��%X����q�<4��EŶ����,����,	^-���� 4�k�*��ة)���1�~�a���5�M-9���r�(�������q�҂�ը�S��z?i���������JS�?��~��4�iӊ��s��<(ziB�n_��p4ޅ y�Ϥ<W�L�wm��O�I��bҾDXOM�Bі)�7ώ1�77N��BC�ը����;q��QU�u/���]cOW6�,a���߉W/�����K0d(��hb�(}pw��Ëc��
��x��O~���R��ݹNR~�pM��Qw�OA�_Ofb҅��^��0��1�%�!���K�����L;��8����D9�-@!{oꉻ���̤r�p�%��m�)��-�um��:���U�C��;�QsW�I^5�P�������x	�D�����Oo��y�[y��|M`7{ZX�aǝJ��'ys�逸�ycCO5%�
�'gk��U�F�[#�tx���i�5C��������z�#jcׂ'�u�G��B�޿Q�H&�����蝖Hp��s��w�Ns
<W�,��%���d��ޣ�GEw��ڮ���%EY�Z|��C�^���Z����@�J�_b�KtEE��It��7Wx]iZzu"=�-�v~����u�ZQ�����J��u@7;bر�e-H�m�����'w:�%�B�G`ka�Q�sH�Y�W���?a�A��^��٫t�/��"�c!�qT���o�����ы�*�*v��(�T·����ד�&M�+�چt?ר�+膒4��*����&95�
�;YvV���L���Ƅ
�1�|���{��\/I0����s��yވ�i
|O�v&.Е�*�ܛ4)�'w?�h��y��8}��x{�OS�y�N�K�O**���d]��w���&�>�]-�Ж��a�B!��uk]'�\8=gC�<�5�yN	{/���&J��ʵ�
�U�΃� G�Y\�Ш�'�G�=�1�}lbn$�_�Y�0��H����w	�Ou�X�+�@�(�ԃP�ݭ	��e|Ry[��j)<�Y��g�敩ԵN��">0d����3�d��t >)�g�����R���>�^N��b���׬S�M��@����*>Td'86�s��j�t�%n���xN��k����}�:N���*���Q0��Z��
��Y��������#���ʢ7�?��6��I�M���0�?)��߬FߵPy�F*>��w��7�ğ�%��T�3ߍ��0����k�w�u� ��8Qkc��GX�uB2F�Q���W�(h���zx�{���C�;�4ծ	�H�o�eʞ�y���㷍y]{{�  �)���h�a���뗾�	[S�+!�6��(�@$���W�L&�i�b[�NlYkǇ ߍ�Z�K�����'?H�k{���0�:Y������6T{������N, ��M�4�^T�=ky��̌���}��[� S�;�h���]N�Hhm>���O��o�������ڬ�F�p��!�s�a�=�|�5u��Wt]@���}���� ��\��v��|��5��T��^
�9��qMu�
3˼��vt�uOmϊ��VV����9���e����d5߹
~�"N�e�s�P������S1��V�i�bO�k��>�������3\T��_�]T|�*v9�Uz*���b`�G'�{�}�<
��q�L���ڧ_e2	��WK�]S30����Se�٭5���VՠB�����A����+���4�"�U�.��P��3��T��0�a�NP@��U�7?W�K�On�>�ͮ�k1� ���1�Ą�h�4 i�m�W+�тR��T8�;,�D��
7�ޞ��0�(p�3�F�Mr�ך��'��|!V�(dVm1�ǫ1��g\�${gLP'<j���Z�Fg8��*�� �2]]N��lI��AMA��lL;?��*���a*��F�8o���[�~���JVV0�A�=�9Z}3�(0�'$J���Z�(���&vЭ��X0� k�5<OMxo����{�:�T�����^���/�*�A����j��s���eb�s�g���ُ0�������;i�]-:˳�w���>����G�~s����nW�"Y�Ī�w)K��[�j��QQ�5�H����Q� 2�谌�hzWb&�&��	�bQ4%R�s���v��*��f�ѩ����B�>;��<E ��YF��c��FN��ҧ�n��b��ʡ�st����h�HI�n'����$�3���pP@4L8��H���M����mO������2[��G<�oTw����;�ٝerU%\|:v�פ�j?>�,A2�M#�d#�6�؛K4��d Y,H\�&���\؋�FV�>�!'�ɏby���c�3=��lI�5_������#��.QB�<��0D�}t[�*�2e����;n�w�B��^u�=�����jF���|��K)W�d��.!���F�F��*J�l���x�ͫʲ�Gy��ɤ艆[��h�澦B{����M".I�󗼻�F �����'0>u-_���#����HE��UA�*},Y6�z��n��,�&���%{�*\���.�+�3�3j��M�ޙH��~皬�mf>9�6������/��9��K�3�\��@!�����FU�k���U|�u���2�|\�+���Lˀ�۠�fٸ�C��=
�\}f2G�{��P���X�rX�6�p1�L�+\I&WIf:*���Yu,��Q1�N{(�rE�)"#��e��~L�t���_�3���� ���}���e�gD���W�̽�Z)��#��o��݀(��ߡ&*�2�[h�1D8�w먀���?2MÊ�\��	��\��z�jI��؋X�Z]�XWU��ۂ��b6v�y������	B����w�4&�،��H�O�x��Q�,�z��_�����"���~�Uy��v�Bx�k�9�(�٧�.��9qP�+=�˧&�;<��|m9՘�]����K��ei)����GE��u���t���^�v9�Sƃ��+R�{��e��%,|BIk�4n��(�x�m8A�,-9�7:�&:.�@�L��09��F��[�U�>�9�wE{��I]�}okzll�H�R�)��]_waok
�AX#����R#����u�ɩ����o��n}�h�}�����~�D��:s����BK�s.���73��yF3��� :I� ��+���SJ�F�
�e-f��?�A�H�[J��������U����̋g�ʪCWK��D�f�:�d���"��h�G��/.3�]���y��8}�%+sko>�n;�u�Q��W@�&z�yU��1�zq��蜽�*���d���cJ�+�I�wi�#Ъ�^�i�_�ҵ+
�U?ƾNF�� i Ni�i���y�g�k�Ӵ�賜���-�M������d�����1,�0�[A�H��5����I���)�O �9ǲ�Yet��	4�������)rX�IJ*�f����U�o¯��;��C�h�P�Qm���|�p���L]D�>�D��K����躌L��k����&Z����<�xW�*�
r~��^X�7Q��c���g&c�H�c��]�D�x�~F�b5m��U�j�O�x�=����h�ucK�����pK���?iį�� wc_,x�[ܭ�F�����H^!�}k������M��� �]�a�4�jd�����GQ�*(m�{Cο�V��;;[±句��e�������f��黡j�/{? /��6 ��L��P(��1�Yڣc�@��U�¿jܭE������˖k���aY\^dO�R���5�x��n�4I��Sft�`5:��N�ت�&O�O���F�6^p�˴袆�����v?����G��+_BB�;;�_�)Z�8�,�����ؖ��-���4<��[����v����У�k�%����@�[6-�a��:H��c�ʻd0���o.e���0�������� �c��	PF���m����2�Wp,��h�1�`l��e�}t��O��,�G���1܆�/�~4��w���^2	w�[�G/v�����N��q��Y�y�;����uY��f�&�Y���q�w�w:V+[�}7KI���D��U9Se�Ԉ���<�l���;�>׺N+ P=K/{$��_�>�`�ƻ�Fk��:Z�&��X�@��(Z��62�mk�-dp%��#����7�p��8��?�ub�:��f��a�dW�>b+�C��o &ź��.#7 �ۂBU�
��c��`���޷��v�lɧ2�1F0Oߟ��i�W�ޠZ����1�|��F�m�~�|�����b����*��0��kIum�n�����]�:�$yeXqe;U��X���9|��V���.�}6����i~�ż�d�z�=�����*{s�0�(*�l�f�hsU\7$%�Tqz��Z�݉��H��C�4�������Q�{gv�]v.k��hu9U,�zq��YF@p�wqE
���@�e��N�3+ڜ�o8Ֆrgg87�����cMP�Q1@C�,��砷
_��JK�r;��,mB�7�T
���9�Zx]czTF��8j$=*'$��}�nU<� ��?'��TT���a���N��f@ӯ�`�G����zي[�|��ixԪ�$h��/Ο���m/�_hVy��x�O�#on�����@L��s�rk�[��q��Co+�a��%L�p-Mn*��l�T��F?2��z�������*�!I��|��SΑ;��Ԃ�Ȥ%��_d���J��[ܾsl��yު7j���������c�SX�T�_�K��m5>�k�SWdk1DGrӼwrp�+)��tI���l����O ��ϲ+~ �0�,�����$B~��]�p9� �+2�t	~᪨�dG�g�=�I��
���~x蚮/��LR�δ^i����I��k�]�Q9#m��坝RPWX@t��r���'��G��P8���c�Np��Ih��C}>SE~��.h�=i#������X��Ee�qK���<ꓙ���	
��559��l�k�w賲�0F}j��Y���3��8��q|]Cd�.z���.ZBr��sh�h��>�|E��wc���c���Ӻ���đ�?���i�V3������Oe���.��]h�]��}�W��Ö�x�Fe)���<Q��C�%ĳ|�d�jg&o^'�������~�-ջt,�R��`�V')]�tI+�Y�XU�!���,����L �����>&Ԑs�MD�;�F��ta����I�2��R�H�V��71/�D�l������=m�vy�
�t�vm�t�[�\���8�|�&������k>�i��F9cS3AA.>�C�N��k�)��O�N��Q��˃�7[� ���⼸r��jy��;7@�n���ۮ��&�V	�U*���lI�²�\΢��j{�k�d�Y�G�l���E����-"dn�eԱ�9��`E w��L�5��B�ٳ۝"����e�@۝�GI�ְ�4�*�;���n��0�0O	�%z�>��&�����B�۪��買��q��U����N�10 ���~t�K"�*dBK�;N���
��PN\h-͆lf�q�\����_ˠ�:ʜ�M$Ĉ���'���W��0I��q�T�&<P�&'5��Ej��$2��ͮ��]�t��)R��Y����-?�tUH|�E�@���x�=
�V��KV8F��ɽ��88�Mw�?/���o�Z���u�G�!k�{�C�ϸ%��Q�D�_^�L����BͿ�j6��d�I,J*�ӻ�R/K�UT_8^�=L�c�6�mli����XF����,*�%�i��$��Q8Ϛv�Y�|͔k�vy�~^u��'n�2ޚY�kUW���~���\`�RDK�U�$�v���_�揷�W�:!@�~�%*�V��eX���"^��0��Qw[�F5�	���,�7.��l�E�M�.�+쟞uY����@�Ϭ�΂��fS.c2��fRϩ�7C��3���&�u�����w���Fɷ��p�<�\��ŏ;l�C��f/�8��̠0�q��ty�9������_G�.��g�ݵ{�L��So���i��mE�Xr=�*�a_��ą�LN���|{�~���Ryh�����G ���,��g�����0�����ߍ��C��9OE�X�6����Ҫ��{�4.� O9�輸���ywPz��>��T���'��ڟ�z7\�!�Le���mƨ��H�e���u�:������/Pa%�u��Q��S�9�[��6�آD��s���m%UgZ�ܖ0���\���و\U���V�ΝJ������:�E/�-������N���앎q"�[]��2?bBG�J���L�t����"eo�����eeL��=	Z�w~ilIQT���y��E�rݪ	����W������pY8��r�����ۤ&T~�r3jѝK6+Z#u^�cз�Y���n��S�E�����p��*eq�K੯��TK���m
,[����l>��S#��� o1-
�
�^���+���{�M�˯jȴu�L��=�<Z��.t)�@���A��LeX�a~!�36�@�Ġ�0s]E<��QNK�
G�'��k ��* \�hU{+�?�a��fD���$Wl��ɩ��|�Y������d���J:(Xs���J�������fY�ۯ���*ig�$-B��g( ��E�+C�>���C���~)(����~���&.���  ��n�B��7Q��L鵫/�~����'ϊ��L�	<�`"�6E�'����g=��ey�.���
{� ��> ��|o8��Qc�/�ǯW�LtpNsb�Kx��EnA�X��	���aӅ��Օ���1��A��î�T�ޮ�EE:_�/�ªo����Y�|�ݛ�A�6a�<�y��o{��Zv+	H�S:��/�l��'��w/H������>f���G�ή�w��(�������$�VW ��6�JP��ou��-Pg�u�����������髶::�|����̼(��-d�Ɍ�"��(�0����`� ��F��XWcYD*(�d��ˬ=�s�K������tI�jή�����ƭz��"��纕�	�
�.3���X8@�����GEB�{+�K�*B�gu��Z�=���r6�땔gi����5n>�:��o�v�=v��?����L֥uh��������¯��C��m��s����G����������3����U�dGGF�-��96�)V�Ϡ��^���>���� ��K�l� P�+#�p���B��U��W�1�FK]��gJ���L�-��Lv�� ][�,v����۫Q��A?�y�_	��;�X4��Dk��Z��	�U��V���m�to�D/^��p=>͐�zpT���4������.@mu��@dY�}�T���P1�eif���q��'�s�z�ò�Ĳx[(?��KP��maæ��Z��߂����  pdw�2@~-���Ӏ�b3/�qR����c�����{�o��i����to����	j�Z�l´K"a�/���%��c�mg�XhvO,��$�<����q`|������UU��n���LV�$0.����s����jk���N�_Yz�`��F��D,G������R݋Ak��;��d>�g����s�Pl�Ztz�au�Ir�NU���+���3���+��5��KO�����?�԰�͟P�a7�90ժ�h*P>�/�H�7�2��.��>���I�z���h����Tyr�|�z7Kk�NyYPP���r]��o,�T�a�,\�2yC�q?�����s���n�%�� V��nr�"��r��$�
�d�*k��jȖe�D1s�P��.t�����B ݐӍ˒b*���$����0�0�Pq�(_�uF�6 P@�J���f�ƫ�7^��΋�$��l�Ͻ�o�K�~��`��bO�3;,�T��GS���)Jl���m.&K�)F�8Ja'=�a�1���L�Qڥƙ���:�:��ABJd��I\g�0pUǷ�D���/�� �p_�&�f�(�]�\�>�l�4e��j`��,b�	0�!\6�PZ�����|���|��yP�kf�S�#gߓ!v3c�g��gB�c3�uWx�����.#�7��3@Hq��u  h���v�z�w;�?�ΒM�_���0_�90���k����ȯ�!�� �I1B<�[�h�ii��	�ޜ�u;a��u4%P��1���]��RA�.�J��=:�̒��={7��D��ڍ"�������G�l�ښ�0���Y�%u�m����e��3; ��eD?6[���!�����\/��ǐWcݎ�:�Mج����x[T�-w�뺵5N��(�o w�i��U׎z`F�^Pu)������C�Q}���ϟ��g�/��������R�!](�xc'��l�4����9F��m��Ը�ce���zF�֙�N�ʂ?���fA�H�����i�3U�n�3H�Dl��ɖv�ZjW��Ed`���VuLN�Ć����m$e��J��e�B �(�ޣ>t?\��Ĥk�?�T� �B�F�'{XC���&l ��W��.��+�3��N��a���`��$%��O�&����+�a�;H��2��3ɅF� "" `rL�Q�G�\`$�^��M�� ���6/��.#�T,U$O1���7V-�1��,<�^�rci�����Zb�<��@�����)�P[r�fo|A�u1!��O��2�.��Q���z�$�q��Rn� ��0��y�>��M�A3�m��
^�/B/�
��מ�Il1H2�Q����WU_MuZ������� �Lz(�mk@��}�S�Dt�v	5�^�Ӧ���g�oݻ<xqU�P$z���c/g��Ő&f����������j� @�[M�Rꐎ��X7�V����z����c�AVҪͰ�x�� Y��m[�JC���]1C�R��c�g$β> v������ϡ� �[�OKYېGo}�]��҉z<��Ж�=i�t�����0���ݰ�+���P�B���a)&���S�j�<*�)
�2�~�d�� k ���Jt���!��l��r����B��Qlg�!Ǔ���W��LM�[_��G���m�r�l���Z3�W  O��}�'�F������f+���ο*�l�����Xϭ�����im#���8P�g�K����,���Gzip��0�����ą�_��u܇l��B��_�T����&�]�֜U<+
��sh��Ϡ��;`A�_��J[�xV��lLh�,u}Wb
^�閳#l&�O9�ŷ˙N��iƲڔ]�Xy�x�mLر�o����Oː3]��na�����e�g�N��Y�G�AT��V�\�]և$��j}59>Ζ4��;�^�n~q���,\I��F!�2KS��ݟx�Dm�X怿}h7=	��
�����1�/^�!t�D�z�A����a�}�=7솋d�1'�+k1�������1���On<���0�Lt��`�^��|�q��<H�њ�!� �j�%e�� ��'^���b�Ѯ�rїJ�!~+��;�|�1�-8q4xNW��;�X�v�)���n1���ԦH�u��P���:����_�f�#dqڍI�L�p�W�A$ȜƦ�t�Gk������I�+��c��Т��6�u#���	Խ�5+�H��K�`j"H��W�%s���L�<������6*��I3�}K�ی�h.]z"�F���$`��:QJ相v�Y��� r���(�<��K��7�}]�$�������/�uVVFd���-N�XlWT�;c:^�K��!�r�[k��۟�M�6�L��(��FGU���4i����P@�Ķ��.,i�ۣ��e��3����^�����l���J�h�Nx���4?Y0D�\����%�G4���T���_�h6
0�ô��g����@��٭n�L֪_t���U5�0U��3"�6�*�,�����0�y`�w�/w����їAfG�Qcڍ6YnC����6 y1�Dz �HW�u�5�N��Z��J/�@�}�^t�'�٫�M�4� �j~�o*�v�Q'�A	��ZH�`KE�I	�Y���d
O�*�DE��mĄ�D�s��˾
I�8���Z_���yi�W>2w��7�D?�^�Xoo�2���}��[p'�,`.���۟�^��c]D%6�Ƌ�;���	o�\c-�Ͽtf	��sY��]<�~Y��J��,��<s��]�2�g/���ᕜ��\:fA�J[����iܿ����2�N���/[7-�47�gl������z}��|ɪ�z���o�K`���h��р��"�Z��4/Μ\�;����7pUXɄ
g#v�y��?�P��i���v�M��jѻc�"Dd�n�:��~�8�t�����v���8�yS���ߎ��J��V+���6�큗�q+����$�X !?O��(_��]�_�>%_�ޫ^:�A���I���Y����JM�R��w�
7Z�k	�F���v��n��{h��f�Ws#����T��F0ID]Q~Ƥڗ���a���5;$���FƬE��
�i�e�q;�-m�4o����W'��5�?���H��`�+oe�篧9<󞾹�*�3ǦF9�2K��މ���N�Y?��mD�*˽!z����:&N�f+�#%� ���yNL�$|P���dTS~Ǽ�: ���
RX����ҕ(���9ۃX!;WCdvk��V������]���'��.��;�kO�_�/IcI���L�<�/X��dt�%6򥬭�j[vo�=��a�&�R�Z����R3��x0r7P
9�W�猷���Kek^��i'>�	���$U���w��rF�h �\0��X6�d| �Z ����ha����=)@�"�JY��k/��? �9-mlU}e�f�����ɂ`�E�����e.�hF�zDB0�SGyH�32?����1\I��0���m@���׋���~� ����?�>$�������GmQ��=�
N�Q^������7���~�:�9gR���w��x�Mo��r���@��
r��a5�ٹ���o��X�n��q�K}�.3���γ��&)���M��nfYl�*��2�-�u-�Q;�(�Aj�P�2�?��W�Xe��Ac4�AF/QT;�BAɬ>�`Xsͤ�,mo�����l�� �x���ŗ�~�|�ܬ�J��DyT�=ZT��M`4�T��jv��[l���Bss�);&�,�I��zK��Z3���h��>��TqΔ1pG|��� �nmt7u�k��t��osG�T���5@��7���Mn�I�Y�!��ǝ��N�_z��(���T�M����0!�z�hy�C��
���"�Q˛y%u��:���Qƞ�"��S�h����o�}���E�mlz2�`�ٸ���:���l�*4�m�V:!��ٵ1*���odnF���Ղ�e�jҨm�ҚZ�����2�����V}s�n��l�(4���[���-��aB�i��V�%qg��;��~N[2L����}��<���QF�t�^E��L��6�a;���ɛ+�O��@KЖ�1�����~�H� y��&���'����"ǍSƬ�u��2���2C'�L��<:����mI��v�9���h�3MZ ����.Dj�^f�+Ե5���o�N�G�ofj�H�d��&�!�D������Fq�Xi�fX��,�r���8���+��-\ �ܴh���[�]{��G����plA w����C@�����>�e��c9���]�v[�1uB�B����cA'i���
J�
�It��r�a\r�:�:b� ���9�\X��ͬ������D����Xf2����QK�RA�책���� ���C��Ԩ�4��V��!q�U�[x-W0���ߙ�~B���nYc\�=��������a��{��ſr�1����RO�����#}�� �1\!���%���D\\9�*w�����������:��d��l[S����~�ڹ@��q����?��κ�Q�T�9�M�XOͰd�_�J�;���D����:Nن~�Gr�<����������7��g
�o�&�l���Z�`�h���j�!���;ů2t������"^� ����
��%+��%3`���蹯����}8�O�z��M?R���8���Y�{/�KZ���W�9W�5BA \��w��w�
�待;�gY��y?N(XB>\a-�W@n������v�1	M�HXV��&�?������a 51��<�6��`�l��f�$Y�*4���v$� Q"]�Ԍ�r����
�t䣞�{�����&��.�g8g�$W�4w�N/�p����ёE���<����23��~��9�2�S?�F/*�)�4���ot�A��f\�_y�`��8�ꭣ����l�gǨ�7�v���P�}x��c�t��+���y[ҰP;��U�?C��>��}��F��̆yh5�m��߽�
��iC��/7jK
�'_�T,��"��Yy����UN�����P��{�7�s±W�A%S���Hr3[�4�X:K��He�4ҪA�]ʙ*��$8�8F:$��u���ewш/~��|����3z֡h����%�%� S^S���R��������S���vZg)�_��E�DSX ���Lc�T�taV�Z�|C_����b��j�ÕC�=��Aj�]|�H���|Kk:�b�]n�(���X��а<�6?J���G�NEVM�On�^%A��b�굜�.˓ ��e	Axi�D���0�r`|#Zj;���p}�Q=FO���-�F�����YE��.�>-j�{�9y��9&\MYD��>p[��$oь*�yk������Ĭ�b�V ���xP�ة=�ך�	�]r3�oZ'#Q�M����cN���s�
x�C9�-o�.K��B�{�ڡ�b��1?I��N��!5]�鮭UTm��K��i�FS�<��J2���T�;m�q#���;���O��E������.���BGՉ���c�$�����4Q���Ԅ�@��Ոx�aZ��]Z���a#���N�Ͳ{	�{�)��QQ�5`Vޘ��6��ҡ��M�2���\�"3���E5�ut���r]X�n���(����_fU˝w�D~{=�mtL]��g
��D�d��$��&�ڭ!㺆S,￑�r=�=�]t�e�E���l�<�z�nJ1&z�˦��g=#>�>�9p�LU�m3$���m��ʴ�➭A���"$boȠs�����n$���������y���ݹ�V"@����̶����}�ױz���$VL��t��h��f���C���5���e�=�ߞ�[�r�Z%A1*�5��r�kgMcC��dm_�,�oe3�o���������{�p���oX
N5!� F�ED7z/ѻQ3jBD0��މ^� L�:D����:�39ϓs�/��ʇmf��^{��~��޹�o^��,�r���P�������=�9%��ؖ�ł�2v�J���g�`�{�oJy��Dj˼}9��t~ӳhXm֒���/���L�����ؔ<l\��I
ܒCL9Bxu�m��ſ�젛X�@��;	s���?Xs�$�id`��^��lWT�t��
ț�k�F*emS�y#Q�=[\�D+엷����|kH��M�W�ژjY��=bX9�	-3�vƌG
nw�唰��<��Xt<Ɯ�2����lt�mQ�5�C��>O���:�pǾa��^��u�6�r@�Y�iIG��F�0Ӧ�'�nE����:��R��/!�Y�Hv���2J�e���^!m�&��s�e�S�Gx�6]C�Xv+*�|)����i��~��{}�p����uļ���`3��I��cX);@�Sd�,��y���#2��e9ƁQ�%����Y[a���H�ZW�*����|��6'�
&%�b,h��I���G,م�=�~��	T���bNg�xV3J&�[bP��\?��ʓ�Ny��x�9nDg'xB��L3�� �-V b���C}a�c��*&;�G0DY0���P^���9��H1oN4m�z�X#�"�uځcl�53R�V�0�۩��[g�5�}N\����(�h��r+��}��'��K�h;�ԡ76��?���_Z#U,`q����=#�ӟN�*k�_����Uۇ7���<��٬��>��[50:� ��sm�䀘t�7"����V�����A�Z������P��{��"5rM0��H�y����^��$(C�5Ë5�:�g�����lFB��䒐��!@�����W)Jŏ�}�瓓��?�����yf:>3��M<�2N��$P��Tl�P�Q���)>)V����A.J`Mur/���1�:˶��|g��!.��꼜?5�������y-�U�=�{-�2�R�U��l���q63Z4���]���x%q������h	��m��r�˖�����R��,��`������ۓ�j�����Hno.�k����f-��̑{.U�e"�3kN���&��e ��W��V�a�1�g���5b- P��K+܄K�P2C4�������,S*��Ag[�Kp�6�IL��s�SMZ�K��q�3��f��&Z�����nr-���|�	�9�L��=�į���]省��m��I�ǲݡ��7�B�j�0��d���cng/��$�z���\U%H�.���_����&��*d�h����Β���hN{�f�\�컩[���u���ER���^�i�^�����UFy���,�)�Z�#d��/n���($�L>�|�UN���%���"�7����Bm0�A(&PmU�뾐�=���=�7��y�Y9��{�]�E��;�u\�� i�b��(_���"��<� |8���47^`qU����r�+�TX��v,8��EP�����3;%����f����i�A��ds^�3��t���u%#�.m(���q�f3��Q�>���GB��e]�u�q�z~�vq;�������IU?�*�p#����D�2��� �l���b�
�j/��w�����7P_瞰{���촩kX߄�{�-���< A��1��BK& &7a����M'��˗�z��$*J��.m9�؇DR�0��r�׾���-���)��ۜ��ɽ���~�j�@a9G������yv�E�f���Z����ȣ#;�:��Ģ��Ҡ�&�ӻk�subك��H�#�S���V�QBD�y�@���'���R�U��$�T��0�{��Q#�"�7�oIu������߂��k�/�*�̡k_c��S��]��D��a\Yq��1Ȏu;���er�͇��8�u���� ���a��Z	���M��/���tuD~�]��s�/^V���/�+=e���i� ?���}Α���`]����0"]#!�/t�.����/���_S������GI7K��=�)��P�'�K]�Lۻ���:�
�W���?S H�DȪ듃����_Y]��y���'�Ϛk���/�D{��~5�V�!7MT�����5�� �����ӌ׍���$c��e��>���m�����b�+�夽���en����!�~�I��P�'u�:-�����R3`n���A�j�d��S-��M_�����ny��%r�f�E���oԱ��o�r��;Ɓ�E4�$Ww=6ⅵ�9���gj=M-�R�B�6}�<��,�;�%Z&��z\�?41�ֱ�,%�s�E��`�|�Uj����9K*��%�.�� ���"�Ei�}�R���i]?u�ܛ�ԥ/j�=L!f��{V#���aO8ԧ��)���!��|��W�~�X�_Iru��~~W�KH2��	8�u�
��6�۱�jM��W~�0�X??�\�)�Y�r�Ɓ��l�T^}_=q.\���Bu�>�X�v���U�����v�ߎ�������tt<��c�}u��,�~�����Ӎ73"����ҩ�3;_E���Rb��j��C���>�G艳���B�(o?C�	s��aU~b���m�����������o�w}�;y<���uX�l5b��1��r��u�ϩ�
�@�L1
�	O�>v�i�S;�>7��ouo�qU�^B����!Ӕ��i�[��_/+��U[�Y[��5���A.�u����xL�}�_|��	�u?���E��Zu'k���K0���LK%�����Q��wNy��ٟ5�֋�<�O
v�8*8;��˜؈�
B�=}e$~a���fD f�|ۃ�]�8��E��|�,d��6�g���6�|���Q�ĉ;Y)>�f�*V���>|��PKQ��l:\Q��h�m�~ډ���4oG����ߟ�tֱl<~��Re��W���'�nؐ���Hs�f��қ�,8��H*)`��}�1�/���,��V�_}��V����3orKeL���E�G��	H�P>�_>M؍%���-Q7��^a��5X��qe���+� �2��nܝ �LD�\����粃����iP�[/�����f��(%�|d�pkIq���OcR�>DI���Jc)8nF��'EE��*e��J4ˁC3�L�s��5ę|-�l}�)�}��*��5bGf��$�P�LF��Uc����>�-��[��k�'��
����"3���ny�y�GI2�NQ;�>����S���NJO�������e��6x��[H�����<��6��x��g�i�|�M��!��}g2)���S�	�t� ����ٶ�>j�s�pp�y���������1EuuL�c�Ոx��Ϧ��D��y�'��b�x�_hb�[�I��HW)oe&�e^�4��E��������L��R'�^�Xy�e��њkVB���m�4�����7G�)���n=�|��=s&oR���ӊAU}��*s�ˏ����ó�;�>�C�+��<=��@p%���a����%��z;�Nʮx�@�,��J%~�wUJ��e�rX[����Cz3u�S���)dށw�DA�o<�.2��9;
�o�|+2�yk��kg:&�4�CO�s,%dEi�4Ŏm�o�}x35`�-@z�<Mq�}��*�7%}ߜ��I��ID�����R"���)���>_�%�]ޣ[��eA������U�l��,�3D����.���-���)Ju�R�N���d������w��C������32�O�B�������TL��}�b-��m�)�^ �#�e�R��'b�b݃nSH�}҄cXq��B2�kޤO�U]gyv}+��?J���T)v������Gw���˝�ߕ%b{X�;���:N�E}q�E�:B-����Ŷ�D~��S�ri�Ɖ�Q�2�����,Gui��3͈	��d�����=l��b:�L3H�������R%�%�Qޮ�� �sd���Ϣ�g2s1�P�k�Q��Y���e�]U_N��煈v]�)�[���E�4�E _Ԫ�\rC�4�D���0��E����얳g���FS�b�p2s�	�8��T��2��Y~j��WT�<��+�Ի��0x}�{��ӈ[�z��l0��ϩk�c����2�E��7�A��IUV7q�L��U�y��)D��u�m�����p�@Q�z�pm����먬��5�x?��L�s�di�"�)���2� ��0���s	/����9���q�M�N,�������jq���ݒ~ݤ�8�@*L�I'���S��t�{I�YM2eofe���5O��u�E���g���U#Mh� >S�\x��*d�]ZZ*���pSI̵᭠�?Ne�Ӟ%�d������c��%��
!ܜU�����*~D�[�s �ɝ2�k*���]�� ,�CFm�'�~��u�[MD0��Ƀ[��������Dȼx�j��
�B�0 d^U�|�)]V��bw�A�l�O2*1�I�^X�`_����%ހǢ�f���杸)�,��d[H$��;>�o��K:})c�#E{s�q7�<nTW�u�FVʚ'���_73$5�S�D���6�Vnu��Z�AZ�q�DM��#����̽��S�B���Ȯ�*��9֮2����x�D�
8!<F�sn�e���q�ݜն�qNK��l��+���p���lTUV��C��W0s�i�k�ĭ|�p`�d���X�?8HjA� �8�L�r~c�~7q����kb�;���߂�`�������hқ�Kl����f�l�2}��z����q�����-P�i��D2���x��(�T�XԨ�(�$���/d�jԘO�>?}��'�P����C�W���GbՃ��LϬYգ#)ހ}z�ŭ"﷋���S�azt�bV7���WQ4t����7Ԍ�*�!L'W	�3���q����bIT2W�R0��d���~���/�į��jvY��O������Y&�����z��/�lgs>BK��U'nR��཮.��_�>3N�+�o��<O�A�Y���tX�"V�o��m�ٍ�@��<b�*��PJ/�3_q��̋X�};��`"k����Y���Z�g����㵥�T�_���9�����Mҥ��4�A���Cɸs�ri�UFV�?����+8r$'U
�7�m����GF�Z�\��~��HhQ��3��_�RT�;e�+{fU�%�ӉAw�S���v�sGd�TV�G��[�M"	r_/�ݑ�<<=꟔v�n�i5ҧc���M;L����8]��Y�sbf64L�mh��x���@m�h�/`o��<�0��Q�i�����+��sSu`�l1�U��I����0�O���a�!���||a�`���TP�,R�j�jϸD#kH��e��K]D�g��'�w:tQ�˜\Y��̫%tFɰ�e&���J��<����	�ei	� �]e��!�!��xL�HpM���P' �Ⱦe�N�}�0��8ei0�.lbˑ�M�G(F�sy�P~��=-��M
�<�8����(���/#��:dfl��i+|a� ����ʋ��pxz<���ҕ2�J��^6�����s���0@%5���؀Oeɍї3�0��b������8��Z�0��� C���7u�M������|9�c)���ga��R�Ż��1�v��O �z�-�{�W''����˞B�:0x�&�Q��Bӆ��!�2�&�t{�7"�M��j�C�W���_���S��Rڂ��qkѾ���p`�cnH*�.�R�!���]"���v��8Dw�wn��Z�(��Щ�'��:�-	�3�Jm~�:����4�l:��e��X�]�1u��tD}��?E��I�X )`5�D��u��(�nX��ݰL�3՞�������D' �����JPr>����	���N�-#�԰}7vMy��I?�^F�#q��������#K�m��g;�B��&���G��	��סq"�Р��&�aMlQQ�	�_�j���e��]E��I�xq �d�L঻�Wn�-�����4EKFk��|�Nk��Jb�P\����0N�ю,@$m��ǡ=���-��f����M�Oq��\'�V�6xf��ᔋ��~jm�!��Αv��*A�T \��k$�tj����O��ƔŢ��L3�{o��!�Y�n�PPΌOW�U�>��:f�!E��a��2�(z95�<ŽV��@����{s�	�8b�2���;+��:�׶�0�ߴH�>�i����w.*;�!$gSd=�ә�ڍ{ʵKlm+�G��FI]���c�
��~����$]P�{�Ub)�ڈ��g�z��Β���*�95����qT�n0S���Ǯ�j]���UP26��?�Nl��	ʑ�/�oYʯJ[S�:Z*9:��?�J�*��NjK�/,��!���5H;��y?��lb^���hf�<<go�)�]�����5�]�k�0��-	�"7���V'Q
�/8"`>��R�7��
���Ą����B[��z�%�a�H��>�p�/
nH8����7!�-��&4�7L-�M�w[l���U$���(x�%Qj=V#!�Kp4��h{����h���`�ӕw/�X��4f:�@��u-�B�nEPՊMu��f�DV�7���9���uJ�{����,����'�IFG2�J׫����.��{EKvD���NF�]Q�ۯf������Ӛ|��*šAW��ݤ�ܤw�HS2�нj�dq�6_���E�ju	�s-8 ���0-98��3_�p�W,�up�2��;>݁:o�婒9MН�.�T�W��ދ�Xb�^���Mm�ud˄4��*�8��~��_�2�|`C�;�v�}^����n��*Ç�Q3<�=�:˥?��L@���>r�R��+���$[9-���r� l�1 �V�x��CeӅ%!� ^�!���9��o\Y+q���J:3��K��7]<.���3[�ZaL��$�V��|��B�MI H�!7���u�+׿�էF�h����+�d�ݪ��CGt'�}Z���KdV����X�E;u@Me�� `n��3HS��?�[�~ڬ��n�e��������_�)dD3A�
߮�s�C��\o�oTx�,(��ZʅoQ�8q�EIs[������>̫Q�����?^�K55�l'E�B�1�+�c�� A�mIX6�䬱���Xs-��Bl����� �d�jURXa��)y"��}.{nع�j�ڡdR���(l���x�VīH����%��4��T�p�^����=N.2�h+}��>h���&7�� CV���y���q~�����#Jk��t�C9�F�,���68�� p�\�����3^*�Z(/�L> ��╧�R�]%��m����n�L8oއ�K�U�13u�Îͯ]��ĽS�7���Fs�t�;��1U(=�Wi�W5Rg˷�n�8��熰f�8��Z�h�*��JN������6L���E_�7{�B�Hɨ;H�Sv�Tg��,x�&_�h(-zde�k�/W��PՖ�������\��2��`Qx�^5�� ��� �"����Tw�)ą�暓�\Z�,~��:��9xb�~#���ٌ磐�}����4��mɯ=��4�����TR{�c�ʱ��\�ڐ����������Q�O������jxVf�%`���i��X_�3��]j��������l�כ3(��]��"��! 9=vI3>�%���E�ӄ1����H+��$����B���H�Ś�M�0�z竾nɫ�3p��^}����ƺ�ҷ�vi�m}�NW��������U�i�L�=M�fw8�gd�,b�h`�A�=PR��z��xR�'�:���IB��r~���e��ݩ�$f��@[3��]$���I��L;�&r!�f�L��}51����V�̿��A������tU|gq���+�w�H�g�I��"���Y����tz��=̥��3��L~���r�qE�qQ2:IP��h)5�0_6���T@���<��˫��/�\Һ�96F�I��:�r��I�94�Vg'�c��!�����$D�ʙ��:_���0���Ȓv&�ElZ]o�5Nε��4��R�M6���T�Q:�9�%]��{x:�O%��o^-�aп�hB�DUn}�|3��Q�����ˇa#S������C�`��V�V�Ѕl{��~5�K�~�(��'��o�-A�Nj���������i�z�8��u�i�h������ҜV�~����r�T�����5���u�����&�ӯ���7�z6��g�������i�#�Ȣ�n���ܪ}RD�9�
y8v��K��\���p���nK+hJ��F;��G����^�T��"��ƌZ�B�Y��J�g �Ի�G���d7:)���ejw����N����ư�?*UY����j-vdg�+Ґ�-]e�6G������s�Tl�L�w5�Kg�a�,��94*�q�Dnמz)���ƲJ�@4a�ˎ.�͞�îFԌ��zd=wg/���/���t.)	���ޮ��/�󏒲U;S(�M=�Ҳ�:�9�̌����-�OT_;T~sb�����8(�,KL=���� Mm>n �g*�."`�J��o7�	B��Z[����z`��>�F��o���3�������v�q}����?��S�)h�����_��R���h=�5H�G�8��`�ZI����J�(�:iC�/�uz��ğJ���f� 1��V�Ieǁ�[$�Z�����̥%�)�"CY�-����Ϡ*��.�����Q~h�����WK(����'{�9w�&^D�l�`��_m>��I#��ՠ����v��M�+�q�ؖ�C��/P.m�ө�noУ7�-]~��	�R�M�q>��9w>k��O�B(jnN4�ZS%��G	F�Y<Ե�����^�f�1���&k���7pY�~k$�8�_]�?L����~o�)h�I��}�w��Nb�0�r(���2����P�T�ϒ2�X��.�6��CM��'��@Zp���O"�&�c��Z�5��+i����W��:��1�_�����m&ٶRG�2���P�:=[>h�P4���_3rdY(O��
G��PH��c`�R�LDt`_�uK�g�d�}}���L}B2�fV�e�Ō:�{+�5e#J�t���ɳ��m�n�<F��J��#�c�M����>Uk���������1U�$���%��<=�*�j<���U1��d3y�#�l�D<b�S[n=�%��̘SG�a8�rw�뿁� �Т�dŅ��Z�{�}2�E4=�"u�n����n��s�ڊc��}wr�+��֏�^��8B*�%��k�ވ�5/���A����n�x�-q�4�Ҧ,(p��x��	�N�}���ң�6��?�wC}5x����pq#,L��}�⷏_^���/;�6�6ݽ�I<Kuj��ǒ��LD���@���.~
�_J7��֥�H����c�S�|���~�BR�}��l���%���Y*3q���\�~>&%�V�b^S�?{�t��M��۟~����_o��֫u��t��Aü9�E��k$����Y|o�A��� p���[��F��M?l%ھ�ȵaSQ�!��\v��F��eݝ�
�b�"���]�R�t=y?Q���Z��5���%�e���i�_T'����A˼�����B�i:G��fQ	�L��5*!�=I��H���혐��9�ЭT��wS�^q�����?R�i �4���q�Ԡ^l!�s�\�4&�^�^E6�S�n�d8II�z,RH��Q��̴�wb6��+����PY��J���1�7Pj��	�7���Cz錛��K��/�V����[yg����ݑY���!���K�%mɫ�P���&Â#��7iX0�,��d��^m��,���˺�������qQ��U48��8ujhg�̄������_����Jd���12R���R�i "Sz�|�K��r!���	��ǃ(�a�I^��3)��4��R���јnG�(�iA�f�;H��E��u'Ȇ7�MI�4ZoK���r�0t��!i�ޔ��� �襆	�&)̞q�1��e�k�Mq@/����ݒ	�O���]�>D�4_�bS,�3�T@w3�pMϺ���X�t}QI�PT+٭+�ǯXRl1�΅O���l��G�#ې�AI�.�ǣ����.�����_��VV]�P\�i�$|\쿣(����Fؾ���/�,�XIe��d��h
a�0";�$$#nr�8u6��
T��^��^@Yax�q-5�WɹOnX�_��ҁZ��TXܡDn���ߐ��
tl�I
/�ᦕ�.iC|5�ʗ�b��l���&�5��~�כNj���������F���lp˔E�Ű0�p��n��QU��@^Y�U�z������7�>��?2��H��~{�J���ӫ�����r���|̓��ʗhL��Ť�A����*�-y�"*Q�.��|kP}�����iX���������W��-v��A���+?��K�Ӂ�E�&]qt�MBh�J�\ #(3�Wpe_k:ҏz��2e+��5�:�0&�)�>syN�i3�'���j��-
c��d����~�V��St�r��%g'&8�ށFk����t>�����hl�$�U����l9	��*Q�44��a����<#a���!/V?̿q��%[y6�0����`�G�r���rDҾ!�V�2����]);���?Ζ�1���� ǳ�*�J��/�6a��2i1���nʑ��Z��hU��DS�Z����G�ǯO:��q[|�9y�&e�/Ȏ���+���Q�O-J�������B8�ί+�0��]�zQ'ʁD���V�R�4)@��Ebօ��e�]�|�5�Fԭ���T@O�*��0�v�U��ޣ��	�g�i��TL��-(�W%F.V�Ĉ������[R�T?
��0Mg��E")�ƿ��Sa�2���\͂j����١�+Ղrp�|��Xז�f~�K�����(����V��w7b�=[s�(���[�)��Mο��|���lm�L[Hd`&�y������6N��q�����ͨ=��~<����-�^�	N����I��54�^Q-p���eQ����<�J��mL�Ȩ��6Oޘ�O�JZv�b��	ف �d��܂Lu�����xe	U
l����[��4W%r̵�H����n@�a�U��W�'3�/�+�m�X��*��}�m |V�� H21���Z�I�!����-c�ĥ��<�
�82��=Gr8�_��čb��,����or�~���ю0��=����+�>�Ҁ��n�����n����0�����vg�k7�0�i����Kɑ�<��~�(��/��خ���ctY �Pݺu��R����P�1i����n����*Gڨf�U3�7/��4cl����3{J�19�b�uq
0?ċV��6���	�����O��8�)KYt�pu���Е~���h�+�r}i�M�c�3������T_�^i����2ؘ����X~~{��p��ٗNE�W���k���Z�Ǵlt�Z���V�F���_��l}�{2Ԑ^�&�q?s��co���XTJ+���ȗ�J���s#]��S���b@4zT#��Bj���5\㗂ܺF�>9�H%���r{�M�����QG�Y�U�O�nqs�-��)�O�sl~������:�T\H�����y�H�(ҳ8�q��f2�S��H���3�3� ʫ���O�mJp��'h�:�t�xv.�nʿ��E9*o�}J<���\ϋ�������#���TE���q~r���Y*��T2�Yc�X �=&`qh%���p�g|0x�i�~qA�.�zh���o���Wu��4��1����5Wx�=��@
v���DobS��-!�]�+�8x8Xۥ�	�Xu;<z����:�E����̌��0��Q�fwץ�T+�)���}���x6���#���[�����:�b�揑��tY���q�%��-���87B�E���L��h�D�����n
X�]�0շwL��˙�o��B6q�!�a�z����՞��9�Uh�C��+��z�����ЩP�=����f�%Fp����$���R������7����+E�n��f{OJ��vsW�-4�n�N�}|Q/&ӾI������u�k���k:�=��#8��X���>rh�^���rY�F��f�J�1��?F:e�r׼ji�.餩]�|��jDL�Ejw���W���˂�um�$�2�M��0(���������΀N�R7Oʠ�f��/��.��6W�n����Cy�BNEcj�Z�p	���P� ���?�c-T�]B.����YZy2�3D�6͸��ò4Z#}W�?�]H���A���sy������c���RA9FM���LG�?��n��\���x-�U��0���.���ދMOj�R�9DV^��Qۭ*�vgH�u�oBR�8o�
g�ST�����>�Ȩ;识�U����V���X�����?�� ����4����hpq.��ʓ�Hv�ݖr�������AgȾm�؊Nђ��u�'���T����3R˔��)&���	��:=gB�\'�c���S;�\�:�HQ�R�����*�-�xVO���B]����{�������u-�A�d	֦ɱ6�S�ň͢8�?�%*6O-C�@%Y0rX9]�_�Ԏ��؆Ù}����`�%��>�u�@:gI����3�OϞ��t��������zXA^��`'u}�u�w�?���ʃ����ϳ���..
��A��#��9��e��L�?��橁����M����,��M����y��Yh��&�v}]�Sk9�TK�^��x�*�:�+\>�rH��wR�?�k�n���*��B�9��l�='*��`�|;\�f�~�~@��k�x�#O�V�Hw�����n�Q��0Ƒ���!�g'P,�kU�fC\�L�T�N�(cž��n|_�c	���۟��,��e�S�:�6�6��9�����1�[�G��ٶ��p($�7�v�N�K�gbn��=Y��	�� &�p�eAb�7fEB��_��gvSd�U���>��V�b/��z�!�ĳӍ�M,�1Q63�ς���w�������!̾b��)D��眭���`�Wn[r~���	��caXP��VU��HG���Ŀ/����QX�f>��V]J�{ �\	e%O�RPs0�385�/%�F��?A�L�G�;v�pH��b��Pu�`���3g���i.���!���g<¢��]/�ӹ-ef�~�Sܠ�Y:��d'�z��9[�<���ݴ�b|:�	:8(���sQ�^|cE�K����~)���T_�;|?W�^u��Y�r>�tX��kF}�5S�9z����R7V^��x��Oڔ�h/�]�!��񨷱���Q��ѹLڹG-�e��T��S�x3����;�b�P�Q:].%����9}
�*R-I�ç~&wx.�f���}d��H6B�X��{[��A�g����)�� ��?ul�kCY��7��J���*�E�?~�)�i<�]���N�o���E��Xr�o7z�&Dk:
N��I�6�T�HCb�7L\P��K��g���E���_)H�ٓ_���e��'�f����Ik��S�_����WT�;�et;�Ӯ���� �-��k�4]�_ �zF
ζ�������p��]`5�_�0�i�)"t�H�|1gy8�7U*�6�Y�?� �?��,���0��,�)	���k��1�g�88� h��g�v�U<�-�E���۞C	�ӓ^�~����<#���u��-5,��j�JW�>@���7�GF�Q�R�����j��Ժ�m��d�g�����Mx@�p�4.�z�D�S!��_C2G��a��żv�ִ��/�"Q��b�������a�e���ӟ�i�B�zцg/<Պ_�~�X�[�	*�@O��Շ����^�!��х��N,��I��-�>�+%���W	���?��Xp�7�r�6U�P�Q�5>@�Չ�Hx��W����}�܊
���T<Y|���s/��Z;�"6�D���99rԌ�}X_��]�N_�b����d�bR%�{9��x��Gj�H�F~���=lRH��{�УQ�Tv	s�S�b��M�ӟ�Ir�˰E��O�6�&+)��q�^(�`8��ᩕ��-;�zPK�b�X:�,h�Љ���4>�v� RpHf�����<�s>	2�ߝeC�,ܬ=����Y*�a�L�~y��[����r�Ry|��}D�"M�K2<m1�n[�9(S.P�Z#B��J�j�f�2����p�sOi��1��`� �3�-�EsC�tY�a��7U�B߳5��g�L�4L"%S�#�D�(e��h�j�J!�ʴ�p:��|��TN�ߐ�Яz��ݞBE� �W�1U����F۴�'�\�ٛu��M6S�j�Y���	C�_"���������K^�jf�mH��[A�� ��z��2���O��8�7�BO���F'����ow��-h��ht�Qk��z_��O]�����(��18/c�n8��әGz����G�����޴�V�h^?�K��w�hH���:�����)6yOKT�2=��,�u�"M;��}�j��Bg�S#�1�c3q978���,G����b\��:d�;e��R�׈fN�2h7��0���D���E�����7XNy���%VQ��ޛ:p�Sִ�"]��NE�)#C����P,y�Xve��kU����Ƴ4�Rŵd��;4P��16Ì,��!y-�B��`9��u�Ln���4��m��Cgː�C�C��`��z��H�9�}��1�f�Rb���o��א2g�\��LT�Om��
)M�5���AH���B�|e��!N�.0楝�O.����[��R�aKw1JW�� �W��IYIf�煾_�.J	�[1F5[Ō��)xtk͚>0����q��B��~U<����h�B�shwM�
�q�>����^��k�ܖ�m<:B\VY��e
h?�sw�q����If�k��[�4�W6�����Yz8��V�x'P
��,���l��w��A��DLOى-$��x�t��ڮ�Y��g# �8��E�Pz���礷��ZB�(�š�hEtIn�����vy{v������,�q(�nU���9�x�B�5�{���3$�&��z�ǭ�h	{�Ʃ��6a��������^����,W��rx���]��y3c�}�7O"D����gNFc�TH�mT�ei�Y�?%�g:�T��D��fU�n���{	���I��x��Ԧ�����}�� Y�K)˨nu'��0�(�NL�ܷ���a��^��~�oݒ�q�#�_բ�l�p�W���Z�6Y�yƙ;����SK{G^�䆦��-W���_CS�l��W�G��{)�=���9�8�W2O\ɜ,R��leaf����>cm��H��WbEJN/�'��Q����L.u��cI�M�sؘJ��cd	q�:&�h�o��,�i)jL�#���WF�@�R�^��i��/[,�;��١?�ݳ�v���Y�l�J椽ă�F��ך��<�0 jā>66s�}���R9��e�q��c�g/��C��?��'U�LDR�� t�+j^�_�(�ۂZ���t�Z�١��lb��ƒ��[��H�M�8n	���d�c^��%�z�z�2KV�ʌ�v3��\����h�,���^(7��>���~�Z�������-X�R���q���yi�)��i�ꈣ��s���=��,QC <�������N����d�@88>���? ���Tՠ��~��|�ty�U�;���&eIEOѲ*t�V��d.�:�@ʲ���קE����w�K[_ tM��\�S�獣(
�Rc�G+�%X	�E!���~ ��|�[a�Z��	u7�[�ͬ�.��f����M�SM��?�;�=�0́����Fw��G��B�w���I�.԰����� +L&%��T��3�a�I���tAei���s�w�,]$�'�ѝ�b�+��Ĉ��,���M��e�5�Ҍɫ� j��P��x� ��o.*�F$ŒY�>������T5�X�_k(���ʧ��x���S�1>"��מ��ɭ�8_�\w1*̡����}����y�qfّ�����H��N�9E�᠗+�n�����vC�x�eA�u&���c�)vYq�=���(�Gg�Ӿ��l���EÁ������oM:,3���m	�	d?�pϗ�͖�#d�A��r�-�dUJh� :W����������P$�����@��U)e�C�7�X�dz.���g�d�nE������T�R]��X%0��/f]��m�j�㨴ݰ;g��;����@��8���ws_rc=��yrn?q���{���&,ψ���]��l��ur�VIxV
�n�$�ŁH���`�h<��t!J�j�DV��8uIn.fV�j�AUt��v�4�����l㈦5�������h)S
_h�j��W��ni«1�Έ�5cʫ:}��?Q.�R�uH�^���7�@G�����SLL��E$Z֬ai����F��D�eۈC��T��Q_��|^)`��xZ����&ڜ���["_qV.q�d$K1�7�m6j<�5�������x��/�3�����#q� r���3���㻋e�J�8�x��\�W�����d�HF����b�S�A-7o�.h��s;"l7Η�~V"���c���g���j��)7�O�1}�leg��-L�=�o����#�ٔ8=���-EEF-H�$�0�B.�)��J�b5c�BcF��L��IS���N4RtSI�`e��_�g����Ne��%F�F爴A�2t�٢���+5�3
�N1'���L_M1�nΏz6=���,���X7��kX"t�Vg� ��Z�䟧���0��m;m�s#}�����ｭr6�~��{'��.����D�9�-��X�o�Û�;,���_�m�f�+{}u9AL
��av7��a+̯PK� ��T������̞�a�UViV�(�R�KgD:�!@�C@ElH�^��J(J蠀�H	���K"5@(ϝ��{�����+�̙3s�53���+�ے'���~���y"�~���W��\$ڶ������x��������w�@��d>���C���$��;�PbXjl�t<���0�n��+4>�$�c�^H�6j�ڒ���&;�hS-�F���������%H�2�RQ�i��o{q�['�~�_�>!uG� !r����)-[ljh�rέ^Xo�q�:�g�����Qn;�w`d�1�}|���逵B����G�f{�Ƚ��������}�ɞ��K��'��y��&�6��B�tc׸7�{<7��<V�-������0�I�?�����X����hi#��'�7�`��N{������@~|W��l�r����j)a
"�-�,����9[�����V2��{�����4[� ?0F�'0��z�2���e&��_�݀����ZFG����N~�Br��"�Ux��/.=1QOq>X;Q\�����)�~�y1�_����sf�j��35Ʋ@��\�ʊt�..��&��\����F*���ƥ�u�E�F@���ֈ5�<"��z�3��K���k�����[�@$:�H�-X���Dń�}j��j�2ݾ��Xi���r���˧�Nn[���{qJ'�)�B�R�GX8�4�9OV�o�'�Ç]쩃�n�����eŗ��L%{��x+��MS<��ypݡ{�2�Vq��2~�Mm�q3B���A��v��dz�B��d�U��]( ���Q�wґ����P�/�LV^�;�Qys�_�	��k�1^����6�~��0�W��ajK��(F�z�"|��־�F�$T��-=PA����q��<u��Y�&Cy��Z癆E�qX��3�T�5P��J7��hI�чC�KKlE!�>Ã-/{/�&��5������̼�����~�����ΉW����S��:T<�k��]!�>*�������F��z�9���41��8��x�-�x��!�>�>}S-���{Ve��	Tu���N��G(���H	H�;q����<Df�n����U�Oԥq��yD�������e�4qt6��~>(Q�5�g��!�1�#۷YmL�^	4ۉI����O�������<�s��9J%�����҈]=����\
�S'�፾��~������U���♵�3{����T�/�~�� ��c�z4:�MF�.G�T�ѱ��щ�a]V�R]�+�8 �?v�:�z�R�#?���RC�{P�Xo/IL(���7�4=b��Հ�J3�e���y~���֩~���X�^��3���ޱ����f��o�GH��͏z]!+I�>��jC5{�6:����8�N���	��[�GһXq����=��re�߀�f����$,���e�}xu��U��,����F������P�s��X�̧6���Bb��7	-�GGQ^������$'��Y��n@�IOY0�d�<�d8�XA�W�ko��u������ʲ���[��#��,,�̌Uj{]��=�?D�4��v����L<�����o֚[S�ŧ;�U@j����b�X��P�< ǡ��Fq$�sx��*^v���YM#9k�w�w��o��+3��'�ф�,����	����&鹼�Tc�j<��^>|4DX�CK�)@ȪpuM��Ad�8`��f�����!}�����d1����X��=o�4�n4F>B�Ek��{����@�hHb�^d�	�z�AH<�C��PJ�ݮ��T��C��
����t��zUl�R0O��t�q����<��|4!en3�pJ����d���p|����2O��ń�Rs��k&c,��*iu�Y�(��ա|���څz� d�ΖY����/E������Oa��+�F�j����=�R��OT9z���Z|���7�7Z�?L�Pn�C��T9"g���������M'��c������=�3}���L���+TV*����UF�P��T�*?K����B���	+��{v�����)��^m9jd5u�8,ĸ�-�b��H�t���h��:LF	`�4쒤����	�Ĕ�v����7�'Ƹ�!_:n�;%H���o�l��U��t���}��)'�:bzu�'��;�%�=0�\�~x�;x�ܜ&�����/�l~��G�k�+ո�ܺ�&Ǫ���+��zmz�^(��$oD�=8.�� �-�^�~��Cr�{M���'�ķ((}<�@Z��n6�¥M<||`]��K�>��bx�zPEn]w9�Gby,�^��G}J���)r���"1�|����'�0�2{���2�%K�s���*�i�ٕ��(�}�zd�8��t��>��&�m�g~�~�
նZQ\�#S�F�h��ه$(�ZU��(�#�.��i���W����4Ѻ:wȌ�~,�Y�c^z��c��ő�^���K�7�u�y50��#4�>}VA�v"S#f%����ۅ؎������X�p���Mr9K�ݡ��E'�Ā�C��������(�TI.	�۽��`��5V�JU3}^�~��vY��ZG�\C�">0�9'uJ�;�o4���RFܫ`X��O5&-!/�Q�.y�>5٫�0���2�f;��.[6���U�(G2�� BV1`eYZц�~�����)���F/���h�N��:uNn�sٵ�厠��y�������#��]o_����6���e����1�#/]�����|��ջ�չ4�v���~���P�a��Ѓ&�;Q�w�)[�����O��*B���Qn���`$� ���jtU�ã<�X��Q����k�#��p�y.��w��EEH"�;m�P�k}�0Os����[4E�Ri��3V�#E��=|�����Һ�(g9i����w�p�6-�f���Cd��=�R\���ڳ�0#��NQ#�����p�s�S���o�V�!������U����*_9������b1��$�NQ�@��V	�K�u�����o�y�l$;�e���ϳ�U��ɜj!F	9�V��ݗ��.����D��/�3_��
}8�^P�XN��b �������z�bcޔJ���r~��jhvlW��7cxs�C��u��Z-�r� �����<�R����S[��y��^wD���M�[?P8���s.%��Iw�>��l�W�J���FEsN-RO6��> ��$ؙx�R�*���FU��.�. ��A1vt��.:襇8�`�۔5�T9��t��	cr�C��a�u4�G�+g���W��g��E&7��K��84��V{��;���џ�4�߲�E5ZH��FL�տ:5�$v�f $�EX�{�r���b�6��x�/w#i潋@�.yv��� r��ّ�a_	���`Us�9��������L);_���8.���=���ȠI���v
������hN�!�������g��	�M& .����Ti[ߑ�^�#s0�s��T�+�v���}i�[��/�A1�k�UI�h�QM���2�to�evr-���v/���#���Y��t�_rT7@oV���'�M��(����p3�N���|��
wD�P �1.�2(�=�c�̙�Ŕ�>��зz������J�A��ސoP�bh��Pqb���"����]W�2�ۿ�JT�i�wL�qE�1�����0���SW���Q1��3 ������;�a��ӧR��!?�u���9c}0�����r��7B�����~��Z���N��s]�c9L-���W*�ɵD�@K�Ů�k{Q���W�>G$zAH+̃�_�U�B�RP���v��#?���^S'��:��~�qEM�����E<��)��E�Ԯ�a����.��ħ��Z3W�<v���ǔ/��\ĦZ-\ ��������p��
�G}�ە�u׭��2q����Q����l���}�`����<lڙnA��g��}M�
筷4-�g?�MH��2��Q�.�Q���T�݉�;� T#����`^.��&����͒�*H۩���TC�ia�}�����3�r���L�H]�+`<�*�^G�
�[  �߉l��^�mon+��|�"��ŀ^f�)�7����l1R���7�h0QXC��u���h��zG�-�և��0r�f��˫L5{s*"ε��R�����vy��xB`X��lB.�W���;�~p�>��n����;���zM�WX� ����8F��Hߑ̩������ȒX�Բ�a��+��	6�[hW�t%@�tR��Ə�&v��Ét�	��&��:�,�M���F�� DX�MJ�&���Zۥq,}˱`1�D/��K��E咴�V#��}S;K���i�K9�&�W�1|dJ���q ��O�%�q��L��V��x����Ttq;��f�j�!-2k��*�
�dNr�iP*��Bkk��
n�}WV�b<0 ��
������i��qҿ�B ؒU����#��Ђ��UZ����:�LTg��������V`@�q~J�����X��2#Ӏ;���9o�r&\w��9���u^17h��)
�4ִ4` ~�k,�Z"�U� f�� -�/���{e~����$���T�h��8m��Ɲ�''���2�C�K���A�߬��q讶�����n*e�n��G6P��ʸ�x)F`F�I/�(,���D̠�r��r��~U�+ kX7�Z������EIZ2��W�&ҫr��ן������(�U4V�ֱ��W��̩�O�|��m$�"'� 4+��v�D�4#n��?�l��� W����X�I��;]��kS"2�˸V�E�������l�A$y��Aƛ��v8��Jw(w<���=zt�Ⳟ!�u�v��R�(�"�w��Z��L�xH�c�=�g�� 'o�I�> 0A�a��^��$��-�a�O�f��ծ�Q�G����������l�;�ĖZԾ�i5��y��S�І�9�� ��P)Q�D��cӣДҚ�S؉���sh���4Y�"{�E�Z���5��Ch���γaͭ	i�z9�zS�oX��i�c��H@U}Ҟ6�u}҂&�L�}���à/���Z���iX�P.��R�噵�$�鋁�wgg��7$��;�[���|�/�#?��.�����h�ꄱ4 ��3���,��tc���	�W�WG+��Tyt��{o�9Udo�	�H�E{pB˙R��I�C`i��6���˗2�e_O��9�TJ�P|i��~�a����ѱey��Ch��fI��CS�w�@��C�1[��=.�%�8�=���w|�z%DCcȍԷ���b�O���|t[!*��&^�a�xXw�9Z��[;w����Ŝ��� -�ն_ޜ�1���!�s"�8���hI�wd��a@�Bj���JNSL�;| �K'�_S�3��~T!LL�:�؏�P_�W-�ù���?Uj+�ے���Ǭ?�E^e��+αX�z��س��y
T���v7�K:�?G�=-D�1 ��"o*b>���(!��^��b&��������TV50��&����٥f?5	����P�\��YQ����L��u�VʐH��uX�, q�J�q�������k}�l�-���7;��G��<|�E�Nud7��ܭqX]w)���rj�x]��X�T'��(�F?FD�8ӗ�:��݂p��8�$ }���@��.=��kԚy��[���G�بe%G �I���������dJ��8�Kj�,bd�4E������#{u9Y؄�6N 3Q�Mg��͗�ĥiAY��Wˏr�!S����4y�5�Y�q��t��Yh�4笺�������
uڒzfJ�D��r��<wE���>�+P�۵�.��/j(P�������M�$�KE�W��B*�C��� .�[\p@�������߅w�m7�>Q~��Y�V�.0<&|��CW�TW�Zf�W�'��>�B�%�g� �<)w	�T���nt��>�h�� ;K��KQ�*����}�QQb�7��X�p�^��?��1�>�w7վ��/m�5��S��'����ݲ-��X��n8J˝�ƪ���%���{t0�Q���m ����.<,�� l�Z��4n�YD(��F,�A�z~�V�VKp�5Q��̒��F�M,���6��BV���Pŗ;(1�-:�ȞN��:�����5��Ue��r���aX�׃D��s��c�~0�ۂ���b)� �B�:�O4�ރ�j�{n=���֘��[�!���sl��F����玕�)Դ�y�4d�S���]y��9`/ �k|J\�N�L[�n���]�3QH?[��/����>eV��1E@'N?���DxC	��M�J%�U!g���rk�ݿ�������<�������y�ʹ~�y_^d՜n/'s�*A�<��(��@�ڌ�4��� ��� �O@E�_�Z���[�@hꤴ>��mv@p���y�����1$Y��Z�h;���IP��a��<2zϦ+�u���l���n�KI����7��r�u��;����Wzg��izA��@[i��L�>�桲�bVMу��� &��13ty��� g�A3Ji������H�B0���Ru[����'÷�ty����ĽJ�����/y�e&�GH+�#���*�wI��
��V(�μ0u��a��}N9ҟq�*���zMW��9�����pXIS��u�\�`�5bG�lW{��(��:�=�A�C����tvw�|M��cOi86*�IP_G�H��m|��[��ZA�y<����*M�����v�Թ'A��#~JA'[�P���g�2�h��q\�S����.�@��1d �Jl����#j��c֙�����ĭ�H-t�<SDQ���b��u�]�{FX�񡬫�~��B32,�PD�(3F��t�=b�t�E?�7���PKXq���O���J@����r�y�G����>���"�3'�Yj��>��7��B'�?�N�v? ��_�MF� X�\O=��2������2����ώ���&^^|��8�M������g���{���<��8�l��]��4�cy�dSu��ӮM�#�c�P��M7�S�MC.������ [`p�IB�" |et�'�����\r�؝Iv0d���(����s��K�^e��� nZX�l���k��kd���i\"v�>�1�g��q[�,��)����e�k�z.N��c�^*����q�f���$I� K �a�H��['�}��l��鄅� �-l4^��5\Um�NP����8Q�[�|�]�N��sV:yB�;�u|���x(��]�L�-+�W-�f})��Q�_>WEu!�pŭ^�-2��Q;��g=3�)���L��3RP?o?n���W�uHb#�%�de�����qj�h �!��EŸ�c>�m���Lp
8kQ�ss�7aE̬j�������߉��CH�kO��4��^�'u|��Oz�B�:����qY��{a�^�����,/8d���m�sZ�E��u�ϥb�Ll+k�Pop[]B���g{�fN���b*X�kA�5X��_��>h�o��H�p�eeM���A�3~�7qq�/ӷsg�)��s����g�������t�	�>��9�z��˅�E� �)J
�L� 3}��2U��HV���R�
ș��|M���`�7Z�k�uQ�Mf<�����F"%�I���Vw��)#i��4����0�fn����#CW�������HhG.T�Z�l!���]Q�:KQ4��W��no���DB�i�ʶ�v G	�v��U����s:�tS�L�jۜ�+���������ZT:��k�u�$�"=������ȍ��2,��� 5aYWm�CKJ�xQ���!��`%H0DA3f���:��)P���t%Z�άg}a�\�s��t�W�D�������c��W�Ro1�����o�+T�.��u i��.vc�C-�9����(���z�C$��.��FB�����k��a`�Jx�~ԇ�1�y��A|
�D�����ҋ�EK�D��~`9����'f���%if��9p��T�R����;h`�X���.Z	���
$'0Bw�en� \��������$Y�� ^`���	 ��er\����Ux��V̮1pH�K��i��.Jn�I��K�}�פ%b�Ha���
qB�����	���=���e���P���n����A��Go�glv�+�+~_�Q���c,Ș���>�Ǹ�% ݕ&�S5�����Õ�����I������J�k.���.RkR!1�X�H��~�\��KW������F�BB$`�)��{Β�X:�ꄐ[�����MkI��	�@���J��`�ji@���/޳��$$�4qs.��k����Z�7>�<�K+�:���	�<�٫7��������(��Lˠ�j��6b�ī�m6�[V�H�U��<�I��Mg���+45�.��ӡ�<=�wr�Ɣ�d�K�;Q�{f-~Ӌ]��_~ZxC���d?R��m��rD~��Q�� U�U�2�7Pß�K���
o�:�ܲ�w.����
?I��(��:̧"(
�Z�J`6��Ƅ�Po\�����t��9��G�gT�W�
��b;0��u���@��6CQ���̭_����M�V����	���Ã����gy�#�:K�l�г��do �vH	,NM�ZY�������ޓ4^��7P��	\d>�U��ȶ~'UR L�K���r]B=Q�����%6Lkp���٭"����1����B1��> ��E!�j���~l��'���_L�:V'�w�߯�~�3R��oWw���b���dy���OC��M^w}޵��@%ÿ2߮�:�*E���׶]�+�H���h�(�M���P+x� �u�B�;��/���3?���H�#HI���8&�<�n���������˔��t�Ft����
��ftwp7����֓-��Dݴs2h��%L<C�9�C�+h����_�Z�Ǚ�h�Ub�9|�&�+�"Wn�☍\�;��Ѻ����*ɢ��ב�&�}2k��`�\ؓ�p���	d�I��L��}R���C)t9���-�	�g"�F;
zN3i�PL���/3���(u�����GLzc�#�;wm�>���,ga�����[3�/�7ҶGʎp��Hr�+��H�TL�z����,I6�䷙��*N֨@�8�����~�^�za��*��g��y����٫��	��p)�?�
p�^��-9���j��ͼs��D�'��t���T��u���Nv@V?q�[P������uT��3A�^���NUM��DV�����3�|d����}�TM]�V�gtUi��N=O�a_��eg=�܀vN�5p�a9�b�ؽ�x]n0dn��/�I���xk�g9W�^�J�A4��=������˓8�+r�x��6�M�3+�R8��,����P�u\˵�=�j0����*7J2�B�ܿ�&徫B?�_Nb�>�y$=�rǉ�JkabJ^���l���i>|?a��S�H�q;�P� �b̵
Z��f��ʹc�!��@�9��ș�M��R��I�>��@G���hډ<m�W-A����x�\��w�[��؀�E�/v����ʠ�6{p͉������]��h��OL���D�����K<bۃ_w�o� ��ױX�A�|_�hyž޲R��0�9� ��ѓ��®j��3!{��*q_C4`F�Mv�x���_8��d9y�'��s�s��,�4���Y�QCE=K�c4��C;ٕ�J%������`�/0缠5�-k��~lU��;M9�+i�sc:D-_��1K��:��Y����a(���QYY�胉���9O���E9��6ׂ.���kvw����f�Iwf��8�'%�[v����x���!�`�Vpzy�ZS҂���^$���u7�$3'm��@!#��j�~�;��Ꟈ����;�p���#���m|��ע:XJ��Sg{!�
B1�0�$H��� 2�b�U�Q�u�ө��^E\KN@p��R��܇�G�M��N�Ԏ�l����A�c���)���lI�D����"ő/�DM(O��Q�b(��
�U,�=�_��9��1�6�Y�K��g�i	����#{�-�4�Y��:
�'�M,ib*�./��yQ�E3�ֺ��"������ɻ}�����x8�}gl�j�nnHR�E���#u+�����V��f�(�����VoY�ȕjQFg�}� �s�<X�yp#*���9�ڷ�)O�@̇˱���`~��Z{�:�S\�$cEn����(7C۔�i���״?DSNj^v�H)� t�ċ,�H"�ě�h��JeU���U�k�G��ѻ�q��-x�z�%Y���8��:u�mZ�������v���%(�r�
���Q{/:� ���	9Oj��#�Ở�� mk�sMh��������˧�%Id{�xuz:�������u P� @u�|[�%N��Ƞ��h���.��t�=��1�3`}&�9q!�o.Mw��lZHf=皋�G]�S9����������'�CB��d=c�{�eb�cM�c�=���W�T�KT8!HW��@w1Npi�M�si3�ǷҿvF[H�I�%�n�81�Z-lp��ϝo�7$�_6I��t^\�_t��uկ�Յ�WC������_l��1:�zrx��'�$_V2Ɖǻ�h����+���A(�3����e|`����8�)�����ձ�
��q}�e+��KI씍?_@�"��.A�S *^�qT%��`v�H$w�__��Cp4>)Y[�1z��<����v+�1��TwŽ����1`[�k�TT��{�Kz�=1J��ޟ_@�[�:Sɑ��uI�T�Ro����Y�������ނ6�;`�
K������y=�m�]�Xp���B������@UG �ĵZ�&�ڬ*� ���J����6�󛓻nSM�&$&Y%M�[y�}j���<��f���\���D���<8��B�si�F	��|w�=4�$�U|�������8���d<@�_���n2,�J�R��U1�nod	�[���E9��F��`�\�F>���QV�E����P�K��2�ךmt���}�@�N���	(xQ*=P~�u��{?����s �B�um{�����Eo	�b)3e�&Z�7���c�'�QD{����'i���mΟx�����GoJ6��g,ZvҠ%|g�*?5���L��E�fW5�����_�g����?jp�̑���/��\+Tc6ԁ�?#O��@d��h���w�cв~��(���gil����S@�}�@z�R�6�{P�T@�g�tg3V����*��o�$�/_���v��,��~�ʭ�j�eY4�q�����.p�&.��N+�(�i�Z��ɵ뽇��ӱ����w�����Y�|�� �	1ʿ���6c-��"@��(�Y)��1QH��3�ɒ�J��4�@�ˊ<Q�	�#YnS�ލK�בv�.�;��kڋ]�c����F�0G��~~Y%Ij�����|��8fm�����U�U%1Ě��_:�>������e{��)�1��ۈ��l9 ��V��?����Y�����Y������h�� ��g-h�
I_M���Af*���z�^޽sÉ��G	m؀��IM���Z��쓨"XCcttn�Qu_I�r��K�::E!�n�9���>�a�
,>c�����wnlS��j>�t�E��R���X�N��Q c����C�|������8�e���+�jlb�jm�i)G?�a���"����Q�+��hjL���*_�K�$vF�K�L��@ͻ���?�v��e�Tl�n-����������ip�fP���F$�w���Ā\�?Ɉ+e*@3E���K��L�����Ui;���x�V����h��R%v�����VLL�@����y�Z�91���*�؈ن߰�|����9 �a=E�;�nG)� ����
7�
���_~$�7z^r{�b�P��X�=x��)�P�_��b����	�m�Th�ϵe�Ƅ�(���>�y�l�����y�ߢ>#
�n������jsI7����⭶P��X�o7a�NJb����B�ܟ&>/ǰ�����)�U���j�Ij���&��ct¼Iz�k҆|H�@��N���޴jv�o����S����� ��W%wxT)"M�[��h(��C1�9�~��QZk}g�}"�^'+/S��kbn��tSi�jLs~�:)G��ګ�;'{���k���n:��̴���$������sD�32V�d�oU��$�o�l&s�[��1�..��o�{����s_x��n!-p��d��W�ͳ��ފ^a�թ�&U�}��M뎇G*�Y#	Tb��;,�ڿ�ϻ\�>� �� x]h,L����Ag_��]-���5��a���/��n]<�A_�'�t����`L�c��|�K�����5}?>������z��(���������X�r�h�A�en:N�+�����Û�_*qQg��";E��m|i$�S�0J[��7_�ۄ7��.�?�l��%��)˕�PX��)�<���	��S�����I7j9�R����=�m��Xj���N1�^��K�x��3��9o��j�H.���:�d�>�v�lҽ^�-��j�ݹq3k�Ok�~���������0�y����jˆ���ζ�[��N�<�d�J��[����cAA���npk�AD�M	�W�R!���(��R���2���*�t����hK�)�ܮ�B�_�Z����ߴ�;�����C��.�u�rbf��y)	�9�bא%�.{h��n:~�~�Zp�ALg��6{�x=w�K]5���@BN���5%�iÜn��/�dN����>����z��^i2u��0�gb�c��r�c!�UöQ�W�6=W���v�`=�B.�o��ow���q2z��X̴w�{�Z�c5!��y-t����*�\hU\s���AIo2�Kk��_��OTu,�RttP �b��h쵛w�t�������0n-����"��l��s�I�?pW��*^ĳh��k�[���J#L.\��H��E~ގ�aj�1x�'�<�+�}������p�Ixn3}B�����$S~߂�2$��_^ɾ�#�I�E��z]ŗI6&�]�[T�Nb����y	�Iy�"��NPTT����ъ�t~�F?5y���X}�)��;l�JX'#ކ��o�тs=�;�e�D�7��UG��J�)�STUϾ�=��Й��p�Z�tդ���ݯ��R�?�w��FxF�Џ� �}kf��Z�4&���Ղ�}�T�D��2��{�^$�b�M��9�m�	��AI�Z֓ۮ=~�:�0ӱM�1���E�)r����Ia��P��� qsm�
G5�˗ώ��zę�V�*�;t�h�
n`޲���u��χ�SV����.|b�Bk�ϫ �b(N���GY�8���_em��� ��1��%���+�^$��l������'���Fꂲ���A��E���w��]�r��j �b���պ6;���1U���,0@�1)Q��9tl>m���ѳf܎�g�B�&\���������ʶ��� �Mr1�A'�r���Z�����I�]L��%���?�H�s��J���'��	s%���bd�<�$zec����#c9�Q)[L4C2�#k���%D���U�u!�}w�J�o�g�m� v1DW��V�>�2��&	i���s7�����U�̈������:�lY�c阊�=�Џ�8h���l�s!��GG*���o�FOqQ���?2�x�B�4#���]gY��7|��7����K�v3農���B������g�M�Ea��%���i�_����V���8�)�2_��#� ��ƥI��D�1�W��}e᫧:���_��hp�RD��a���@�|�M��S\���m[��@�u	��
�`��)�M_x�W�s^����D�*_:\��8(��y�oC)^}��eͷ�Q��i�޾ZHcDWK�A	@N��-��L�"�N���wr$�>~�������D�."�N?��!��<���
�����:��L��x"o�:��f鄇h)=� ʚ �[��݅�@���R�	Q�>%��#~~�{r�� ;8d��戀��q�w�������
Y� W�}-�}��XZ�QS��5z
d�M!7��'}Z��\� �lT����ga6u>+������������O���s�VcXYPn��s)6.�����ut�o������mV�<{F��z�ա_ �ګ�,�S�qQ����x�5�Pn��K�4]��@�K���.�)k���v�cJ�Y��-}�s���V�Z}N�]����h��b���,���~׾(��v@v��R�sXR��V~�r\��W7[���"wn��ʰ ����?W45����b�� ��ٗ��Z�N�փ��-�/��n~�.=��Jox��3��ɔ��3�wҹ��(% ��++&	(تr�t��]��?���n�����7��)3(v�s�Vc�`�z��qq����f�á��jy���Iw_��;�4�8YX�ה�Z�(?5���C���>{F��?��^AK������Tr��s�9,�����Ɯ�3(�%���37�Ş�4�ݓ[U���#�0�e�w��gcaYC�݌g.�=:��2�(��H����7���p��-���4\!���xk3��M]���/&J�b{zj	{����5��w����י����2{8��]Tp�n�q��ʋB�p[�{���9�����_���|�6RRي��8N]o��\�.�N\MJ�v�H�ON�֫~{�3�?�$�L�:a��>��Kg�;�xx��gKFB�t���?<\!y�>�f�[Վ���y��]�>�
Ƨx�ι��}{�оj[�f
g������S<�{x�)��(k��?cM@��#��%]��7jD�9J�y�@.��k�م�Bm]������F�]�^�T�2.���IBy�7���R�u�q5?n	yU9-cWS��zII��0K{��'���'��n5���*���ollM0Y3�<t����!4
�.����F�oK�G��.<̪���/?D_J�7�X5ʫ��v�>���E��S�'y�ؔ�j<��:����Gl�?f��.�m���}���z�����:�o��,1,M�n%4����.���KL"귶E�v_A\G8i[���r�D�W涺ԅ�GF輸�="z�:��d=���������aGBX����
^ʷ���&?���r�5���8>�_C�i_����?�"�|���z�v��"���Ԛ��3���P�߻JV�{�s|�gU�ľ�[���p!#�c�N�z�TH�v��1���pm9H�v�B����AJ��#�w�,YzD�r��K����Z����Jb'ٽa���-r_�o�~<��`SP»���-�p����x'>�ɲ�E�E33潊��rΨ(�ƭ'3��A��lW��C���X��ٵiji�����H�[�Ė��Jaۺ�?�>WX앞�w�l��Z��D�T�<-�_�*V!�i	Jmv��m���j��t�u���C�_nT���'Y��mM�ꉂ��g����>-����Zפ�x���_�,�O��H��|�o{/�b����L[���_��<"�l��'?�˾�j�\M,�IQ�s��s��~�Ob��U<�M2���A4~�G�Pa���#W��F�ޅ���w�%�����%E�ƅ��������x���p���Sȍ"������m��C��x��4g�l������ϛՈ��t�oWGc��#�q:�D|v7����#�"�voI�Ռ3�;�b��lz�N�\ˇ�/�O{���ń5̣̜�����mf|�!�Ac��=jtB��>��j��h��־܆s���y���KT�R��q��MfW;�M�m!�T0�Z43:�V^�^aQ=ȦT����8we�O�<�e\<��(����}��5����|����u�gK�%��E�=(R�Ԛ���bW9�}-���6��VZ��Yb��g�k�с��G^�ֱo9]g��S<��H��~��j����h�3)ɫ����@(TM�	��Z Xa��"a�_B�����@|Sb�.Ņ)�6~m���w(.�m�X1uxL����A���џĐ2�G�FZW��?�O|�7	�F��?�U�&]>�sv�m+H���I8X�w���?�FtGe|�}�b�/�����F��_<�3lZ��*�/�E����r��<�Ɛ���K����у�=���D��6��9��o��v����j�Y��cU*�)�oz����ډR-yE�f+��3�zi(��X��_��3��ok�&?��lY3�=�Nd6�t�L�4��޽M��E�I�?��Αз�J����ixX��{�����z��$�6R���[�4������S T���Ӵ���KU�%��Ψ�W�M�Tx	,�� ��d�e~}i�8M��(�O�P���hG�	�1�d������{�$���F���u������7�)�1�ѓ12�E�=j�l��vzq���>*�u=�?�%Qf�OL�lם�c�<@���?�]�����<���l�RG^H���v4��t��3-vj���tq�n~dM�xh��ɮ.���pj1���Vt+c��L�4G:���sc�k�+{����j����XQ����8�-Gl���m$��8��l���v|eʝ�����͕���:��#�f]@��A�v�+	�}$(E}S�=-9A���66���۞�7;�20�W^%�	m��5g����t�������?��l�o�(IGw��I����P��gr�9d�o`2�'�7r�c��>��-]�P·���^c_`_PA(=��]���c��:$��͛6"�YE$|�ͼ���!gb��׹$JX�IND��1�u�!�?��r=���7���5�+q�q�s��[{۰��g:��{�A87����Iv;n8u�՛��uϓ�_�M���>(j��h���GzsPo�fl���A�Z	
��ƩT����������ݽ����o��z��?���P	݄�N�R���q�pJ�ZH5�r�Ƙ:��D19��\Ɲq)Br�}3B��m�����9��k������}�?>�����y��콟�_{?ϳ�VLٝ����*.P�;0ݏ�:.����FO'��H��Da���`F֩���͟�u�\��I�J���,ª����&��o�t�4���d��U:�����:�[W��7�ݲ'�����ډƇ��i;�;>&5e�C�'�'��zm
���F�k,�Xg&H{�\�C�~}����'�Y�/�
5�I:���c�'�Iϩ]nM:�i���h�$��@pAn]D;_˳!'�O�l)o�LUG˓��RU���ߚ���"�Sfg��y_@UJ���h��NgE��/�������'��E��gwr�����x\���)z�5P�'ڢ���y3V04���.����dX�]�h�[>k�컵G�p_����Lf��yJt���Zϯ?�4F8@__�z�?�vK/�`���^�8��y�A�/��o[M�%�(��Z5sp�����8I��_�2&C�����2��G�h
ޅ�s�g��]���ۍ��>���Ά��ϕ�� ��]5E��� b���&��������a�|�̳�����CPt�E�J���8g�޲��:���d��u¥�@ae_�Ul�ǯ$[��?�����\����}��t���F�ڌ��O���ࣇi2�"NǨ���UA�	�Llqcf�v���#��NЪ"���+�n�<%ҫ�׹Y��g����y'�e5�>��^uv��YoO�h�&���9���{�c�Ǚ&���\�oY7.�\p7��[���)���m�������7��Q�98��V�ŗh77�^�3��um�����g������Y�^p*�mK
���	@`�~�}�EX��~��>O�+}�Y���IbA
D��2s2�������o2O�y>K�P�`��B��yv��EJ����[ ����%C.�����h�^����0Z!k�CL��I�ͤ��F=	f����_���cw�4S�\���'���Tz�'��'�0�՚G�ӿU7�o~� �FS��^t���X)7c�(� ��U���k��,�[�Ӥ�+= ���`�F�דB+���D��t�v�?���|@�ƓPG|2���Փ~��SƊ)&���{[7�"�@˴8�(�c�d���O怈�g�����q@�M��O�Y)>j�h��H~T�>ɲ艕���"a+%p>�7�T�fr���QRt<�Cz��z��{��w��o���~s�K���ۊR@����wΒ�4�[�����S5�˳��5b��i���/�O2��^|������Tx~T��Fd���_��-W8���z�u]�Q���|K����I��hY�
ώ_n5�~O�T8[8�P��~z%�T�	n*����� B��B,����`�f[[2く$ō�hy�������c�j��)9�����09� �š6���p1��,�1��ͼ�m�/��^�nlf8h}�������V��t��&n��~�|ŉ(�ɪS��Hg���xxc��s!uN���=�ƎE�v|�}�9����%o��?L����ݦ���_�s���!�{O;���..������ڜ͵��7�z�:P����9��=��=-��'� �jՃڳ��9Okt���aߌ���o�l���VJ��������v&q�*�|1�χ�o����~Cm��L���"F���JF@N�e�1ӑI>x�ox��s��������hw���{i������K~_7�7���k�δ����&���|!S�Rq���\�|��,а���*l���ϵ늏	�K$���*>�9F�5��>�0_�G2�/���G\��ʳ�>���Zڕ�X����L�Gd���H������I��N���;���*ߖvfpW|��4s��������܇٥>�أܸ�������<瞄�ŮN���m l7�6�������J=�_qk���"���a�ƧCS��L��~���)���V��ǡ�M)K7���uk�~�>��큨����^����qt'}xTK��usa\H�Ю��J}Ŷ2!N���`C�R��(d���hE�?��՟!a��q�#A��[�K"��7��;��� G��UT20$t�wxR��}�r�r�s��m2�t���i��0k=�px�ϟ{�)v뙗/����s�(���K�C������1q���e5_��O��}n'�x�o�X�����<�t=LD"X(����Z���K�O�½�i[��g�>��$_�&�>��l�a��%���. r,�b��2����k������l���}�����ot�vvޣOyf�w6l��a���Yh��"�M>M9�_�P[8�Ԧ�DȬ`<�=R��a���x�+ ,�7R5���fT}���#�xy�;���cJ6G�M� �D��u��'&�/�,�����QR�L��'DP��n��D�ٚ���|�y[k xW�l�����X+!m���(��i ���ތq�M��hG���zN2�Iwj6��x����Ĉ�?z٩�g��˅��?-�SދAH�5�l� B�3�1�����3�k�1NF�Ue�.H��L	ءj�\�X- �ۏn�p�yߵ��n;��#��������������4�8����U��YӳG�d�,'����A\���Gt-��x[|��R��H�����﵏0����/�v5���9���P�E9�����P�>��X����@b��^}�c��IC�ӈ�$����������+���<�F΃�+[72��l�0��
\�a+)�ux��e�m1��ƺ�u�h�[��L�Y�XM��������ӗ��3��k�Z0f���C@!`�S*�A+����Z7�g��,�3'�ioUS*��6/.����؋�>	��}��f�K[I��?�"�ɍ��a<~��ļ疵`_1 ؆�U�4�n��)E�iuA3��$=�+6œ_�B9�#C[�8�2Iغ�wC��ĹsN������nss�P��=�X�@�A`X���S�i��'g��{_�Bj�UB'w�ί���]� @4?�zB������/�R}\�A}5Ҙj��o�X����l��%7��{BwpL��m��|�u��r�6&�b����`�UL�Y��_����,PnL],���L�$4��$�o�W=�9e�_,-�?PԀļ���WuR>�V�� AD�Y�nA���P�X��ԟt)��Z���i�4�DJ����b�ߐi��^}b�Wǅi�a�����҄I�M�"��>����R��<�(w;����	w>;��5�w����eeV��D�����{�d��e+T,h�$�	�:{#n�6IKK�)����B4��5����5tjQ�@>oz��}6�$�RxM,w#�5(?ϟ�F,�r�Mq%-\B���>��s�wFNB��40�չ'這�Q`�L�� ��љL��C�V�
dV��BZu^�Y�u}�O�KY�WCrZӆ�o�]a�''�o�;�U��Wjv�:W;t�g�Vl��FEn����ԴND�Ű�<�[��S�g�kX�X�)�n�ԛ"�+k�^��9O�..+P�f~���s)��ؓF'C�`��}��(��6*%�������u�t�O4��t������ɚZ�JZ�[�7��U<�E��Ĺ%!���f���G��PEfN+�PI1��� ��4:BҀ#l��(��$�cf���5a^�!-�B3�c�|���{��ú�F��ʗ3+G
���6C�!�tZO���#��+���Å�BZ�<��5:�Ҭ�75�|��� 7��C,�!ۤ ��҂'G�#���<*��d#���A��.���%��#R�
<h�l�ş/�ѸXo��}!��xmh山�~?f������j	�K���T���L*N�Y�%��0�k�'\�|2+���h��3���ڢ)��Y���O�G���˚�WlZO�8>_��j��~Ya�ƶ��_zA��yV�;�����[s���;��{����V�j��g=)��Q3�FJ`%a��T�G�kV���Ԁj�H���� �5/��DljW�}���(���%2,l�	jω�Z2U�iB{���j�$T���wz�F�a�#^j�Z\�8P�w+��Щ��Ǭ�=�����}��mJx�{��O$7��ܨ9�bpPF���X����f��{��O=z���l t�n�X�MǨ���кɯW�9.t9_���"��B��ǫ!��n���9n@GT\1tm�����i7���V�D�nB��Ʌ4��G���H��\�
-�3׌<�-�.�DӪr�����SI�������)��^+�����,4�{��f�~@\;6г�"'_l�v�#�
ǫ��`��DO�z���;"����SRܢ�
�rm�w+�_E}$��yl�~����ۀ�����tsV'�w!#17N��j*L��oK���"|q-��{��>�>KԶ[Lc�����S�T�]��R������˚ׯ�`F���dq�����JB�>�D�)B��:��4����!�c$DǓa�(� �ɳ/W$V-w|ծ���YRL���]�矾Q:R���bU�7%�L�+�WO�
��Q(o�R�Q99�~��q�Ҹg7�CZA��Po���)��v}y���Z�rO�)"H���+T7��V�Mm�����˰(�>�+�`R��o}"&�[pK=�Ӆ�^i���L�d��0Aǟfe�3w�:K=�-�d��I�[��e��E6!!��sH�kT�%��� �5fz@�P�*Z�8�<V"�A��Ʌ�6E��y��\��KlZ��$�:>��R��a�nn������Zz���7��i��X?ہ�� ��d�!��`gٜ��ѭ�Z3����(��>������q-�A�H����%r\ͫ`|�^-Ά�{�&T�_h�9:FS�Ѭ2�(�G�C�mW�\��c�����f�a�CT�%���U̬[,������Bl��R/SV��]`[� im��]�>s�Y�%�]S0��R�u�kOKG^���(�Y3U^؊��M	@Ϊz��"��~�ȧ߹{W�ۘ���Lor��!)�=��c�F��ӧ��iXx��͔���a���ѐ�N�}c+��b/� G���� ����`{V��2�|U �=�Ɨ#�6Y��u�2��~�)`���{���/�߁~w�7�r^��4V�E=��_�%>p�YX���?�c��� ��>0������u��}��3E�w���afE�z���kR��_��?���C(��l{���S_������mւ��unF˧�O���u%��v� �.`F��� DM���^�%���鋺CĕJt�h��{�lQ�SW>��Ea>*)�����c�==��}2�����|���as���3�tm���aBF-ͫ�xh�F3��b���^���ga�HXt�~�p�6}��9_�#�g��ܵ*%R�˘B��R����ܓ�(�b�"�Hd$�-����@�:��u�jJ\�����|�F2X1g�3W�}�2�HV�;|��9B�p�c�I�TjO��f��Q�7A.����K��~]U�=C(�z�M�R���y��y*�	���\Yq�l
X64�3��!���O��q����琚�W��g|j=Vuz�%�؇��,�����҃�3����L��]�G��3���O��T
��e�y�ȴ��.,ww�u	�<�y��	v3��ɯ�:Oɻ�T��t�dV唴����罋��u�dn��,a�i��ʩ�Bx��e[�b���)�;�RU��*_�GP���Щ�wa����>�Y[l��`LF�ɂ���Cuم���l��k]�S����0��#ֿ���3����)�����T��1cp��Bi�sv�r�?:��Y��������:���!2�j�Z�u���@��/�I�i� �«�4]��f؜�F����Z���U�u���ԃ��o��'��3�<n8�X}l6Џ'�����_t�r����ċ�OXz��_��M�^�׏�su�{�7v+�G��(bkk{Ğ�|���%�7l�~�=0���{Vvʜ��� �����J��y��^?����zd��0&�o�`o�s��TϞ�U�����b@��N��Tw��n�MJr_��.����M����u�<���f|��v <
j�*v�S�޿C�K�4�q\�:�8���Tk�K��{��}.��Z�)B��wq�F0��Yr|�c�]����
X3���gW�m������<(�[��E�h"Ǒ�{�^Y�x��V�W����}��<6�F�C�x�"{�i�	Nj���.�B��J��4�����҃�е`
�2�!��xSWd��^�e�6�J��>�,B�^���8�'M6F'f�5%%� ��{���[�o��#+��؇��rət��,���ڑ��+�'fĖ��6�N��q6@�����"EIOz.��,ao�b@��q��{�4R�~�?5��4�,f52[i�+	���z������Dƫ���\�}X�P|��EAa�OH{�P[/�%�	y�$ ����&�!E.̍^�ڡ뢑|!j�VN��YF�U��}��s���\\5H����Im��I7�SS��>����Y��&H4n��-���n��Z`2}����%��κ���vɁ
���1۩X��v>M�rt�H�w���n�7	C0W�h����X�ʑ�{����t��3��?�������"���s-(B�w^�<��vt�S%<4�0]}h��D���M�X����|ĵ�&�T��h���_�%k�������l��I��0����=i.���\��s���`���%ȷ�����$`Z6�TU��"�X�F�V�m���i�|�F�A/\N�&
:�`��TJ�}� �}T��Cb>ח"T���&ȌY�ݳ�z��c��^���D���]�ri�ң#& ���Gh����se��7lN��Z����vJ��s�Ņ� ��Qo�x� ����e64t��S� )z����Vn@z0��M�,D$M��{�������ޥ��1���X(v�ц���#���^�۾�%Rb)a�:��WV%��mY�����-)4JA%� 0��A5y�7����\V�8�)>u��(^����v��W���"���@jV<eb�>ء:�Hzj���`��j7�F���f���1�E-�W���U�E�1ʾ6���Y�>[�}�E}�8i)�S
3��^fq2EØ�`�8��pA@�n&���}|դnw+e�V��J�>�}�������Y!1-9�s�& ��Z�������q҂.���+�\|߉��41���>��؇}7y�,�/D��-�D�5�f�Dqx���9��Q�� �&FNZ�����`�u߿eG(�X�r���a(��l<�����F)�V��G�|���ZJF�%v�-܁��қ0Nf��E�C�U7����k�)���.�	���g��z���+;$�k);ʁ��^��!�S���1jb9)��)�>bJj��
�grD�����Oos�Xo��G��i�:��W�����6z�73�jx3����>�?�e-A�C7B ���b�7���J���i��\$J`,����R��k; ���Y���S ��s�K�E*hҳ�@�\?��V/|�uQ>�x���{#<�8"�1[}U�E�`$N��E�� �g�@�{1_��z�/�]�� ��"��i/뇇+9����,�}�*����R��M��e�a��c��5��Z�
���'❵�Uv��n�ӕ�A�¨(��m;�Y�0�_Kz�ѓ�F[Q��:Q��#(gzx|��!{Q+���=���yxo/0w//1�▎Z?4z�������'���dqi!��D*���mr�:�ܴ�wD���&&���k��WoK���r����63�E��,R��rn���c��͝	�=dN3#!&�n�@W����b�����>�+��S<�,;�]���^�]�Hm ��r#�	[C���3ZJ�	>�}�������$_o��jh��[P���I2�
�4����_f�ZG�o-��g��Z"!��^+����c(���^�R��ǣ���9i���]i��[1~���'����]�߆�g���7�	������}�l�qm�'8U4�Gk�~]��'YA����5��e�.ktz�\��!$�U��o�Ё���'��81��]���g�ֈ��J�^���C���$EkT#�k ���a�������l�-���T��Q@�Ĩf8�em'�u��~���W�S��)�; o���S�̛�����1$|]�����`����f��=�y>T"v����4%�	��_�2o�e��bz���8(��I��v�ˍ�}�/��W���G\ ��D�yR��L�����m}��Yk������l`qT�_�(�����4g�'�c5��$j,��(:�e��CN���ڏ9W4S��e�?&(=|>;�d����N�	��%��oQ��){\,�V��8���o�:˂��8����]�q�T~n�|W�"�D��M1�l�!s�Ă��'&�ɛ����E�r��9�F�e����:^]i]�a$��@��;�yM���dh@� `�m�x]*�X���:�q����o��K��U�R
j��S*���4���5����]��oUi��;�»��	����x@�Z��y`L;��4��t�A%qT��b�����D�j�t�"�s�L�!��1}4a����`6����ں�n��\D��j��I}��qك�[�u'ʍyC���S �^!`�^��v�_�Ms��N�%Rx�U3��}���{%�(�d^�ӏ��ij��7�RS�X[�b��U���m�P_
���������*�[����*\T�<X�3 �I�*���9uX;`y+ሄz=��I���;�{N��H����|ח����|��u�d��G �t�'��T;$E�b��D=���8�	��+Y'�&�e�� ��9qq�e���	f	���`���gR�s][lr�����f/��g �F�z�� ��a��K���0�P'��~샧�Kn�X��w�̙i��Y��S��>|����v h����*� ئ'tPE�?�wݙD�������WM��-"�[��x�s�p��]�������ѯz�}Q��;���Q��	��=�ܓ��B�k<����rg�fҽoT^�����o�^� �l\���2�U��i{�g��R��.�=9F����#�e�R�Mˑ�T����/1���8����y��3�E!�ߴ�Ij���uj��h'5�%�GCh��}<��HT�y�� "6��v;`�Mno��L�N�8�W�#3f��<"����$>���W��*36�g`���i=���s������
��;�}��p�d~���>���/�X�ґ�#�Y�9෥��H��W�۷\7zntspEK�D�-�)��y�F�v ����j��Sƴ�X�76�HW�e�������\�G����v���7��7m�����n#_�\ch��D� �(6ࡏD�e=4����	��3w܆4��3~>yl���F�3�9���&?ieluh]g}���`F5�[ۛ��(��ۀ�����f#<N;Ǡ�d�*@�a��Շc�Ѳ�_�� �B�;��%�~uVr���?w����"!O�u����u�>ƋH���;̶d��q���s��6��7����2F7G����>����G���3��TQ}V��1H{EP0�����n�[b��(�::���v�F�@~�){�X8��g�A������04V�5q�:��ow�\�Mֻ]��I)"��:ڤ`��C�D��8�ʛҜ�R�����5ЈQH̰�޼3��K�Kqr;�^�0�0S������k��<�q��R�K���s'-�NA�S����5�þ�7�3��K��ݤ�X�t��Ge_�J4P���U}���jFʣ��G�ň}��:��v�%[�Ja#0W�"^�*����7�a]Κ�Κ#�\�F%/?��MΥ�����=A���:o	��<:-�����ژ���Gci2��`\�|ձ�'�{�D���Gy_b=[�d.����VD����B�А4����������1P��a�r�S�a�`[�Pp#!�Գx�Y�~�$K��3����-��̓�Ԩ��H�� }��Dzwb��m>�O�/��X�q�X���A�/�t$�f����ai��jC
�|�����2���(����u���;���v,��JY{m��.��|b���4W�z����}PaS|����A{9���Hj�9S=��d���xܰ˸�ĘZ-%�A�L�~�86���ߗ Z:�au�5�w����m�tC<݂���v�p5�v�dp�*��X��C�1�TQ��v����'�.����������o����E!���Щ�N��3��D<ץz#7�����6�Br��yi m�w�MM)q�5�y�H1��l�����Lp�����T�A���:��+�eG51H�?'��Uu6_���8�/��X��9�t�`�Snա��	�XR᪏4m������� �=!��F�*�Z�6�<��Q��������,r]���r��52��߄�J8�G���=�$MDѹ^8�������� �:�aX�My|����z���
ER�]���W
��p?���o|_�����k��:*+h�OJ2움���*�@�m�{�~��+�Ƭ��D��PT˸/٘s����\6���^N�2%)�.�q�XRv��Q&:���?�Q��DZኋ����}���_E�|V�^����?��E��[ p)�y��;��d�*MØ�1�n�؞�����v�ϙ��4��qJ�ӻT�sp��|4��J��	���V�fn�H\.҃��jg��_\|�$��?�rں�0�m?/a����}��^��h�ƿ(��t���k�志� �I��']�J4H���;�����jo��ŗ��'�-�]7MU�Xz#LD��]����mZ}�1�!S�J/¾�`��{� �[m�?th\��� �ɣz��=���}3�]�_z?6GR���f�'l�U���������k��7����Пa�
���[�A�V���ǉS���#�A��n <_�0n:JT���q�I4�+�Xd+��i�.�xa��2H�BQޓ�X#}a],�����]��=#d�uo-kݸ��vK<��$�j�oi����xs�6�=MbQ4l0"��k??��x{��8)�H��C��W_E�n��%���{!��/o��I�w�{��p!���&>53��>фk1G���,��i'��7�6\4T|�z@���\Mx��&F�'N�w��ðBb˗���h+Iɽ�Kwţ�<�C��׋ݒ��eA L�^zw�T\�܆�ҟ�|���˫>^�P��\{z���8d&.��nMP��������(d�����	���!O�\� HEU �w�/�ﲯ�1c��P�}͞���CQ`���!D����1=���\{㑴e�������p�hq&I��0�}�� �5��J�eL����k�Y�2a� מ��bΨ	ݪ�_)?j5�;c��L�]̪�`o�I_�m`H��b���	����1*r*��j�[ťh��V",S:ڶ
N��*�݌k��V�HDJ%���胦���H�sg}җ�˔)�:/�}�ʦ
K�ݓ����e�U,�Q�H����Ef���x�gJ� 'e٩��<���jЃ]�������`įu�o����n�����3E{D�*S4o�������Z�٣	��r��}��	�Aفm�P�\�y������YK�,�x�]%* `�tg���t�����X�¨�5��(}2O�^Sai�Z �dيJ"��8���"{QZP����0���2�R˜?G����e#Y�8U�m�:��s��_}~�Ud�'54�^ ٮ�L����S�&N��2��\�����ŷ��c�.���f^cƷ��)�Hs��M���$�z�h�y��M7C�E��qR�<
�q#IƝ1={�`s��7�],p%3���4��v{{�,�r�'��M�'�	'.���F�+H�к6�a؊�pA��Y�ڵ�3U���>�o���1M�w�G�{��ٶ��Z����:���W�e��~�J4j�'�Flέ*ܕ��U�\vE��*���U��n��g���S���½��ى'$q��|xF�ڹ�:�J��f�VuEF���w/�Wĵ��h{�J��WK�4��Mpu8����g%&��$��vfA��M�1վ��	��O��_�`��&&G�F�*FH�$	��|����H�x���>l��ths�1�E�W��4r.�S�E�CH4�@ܩ�GG__ �
��"!�ta���Ǵg�ܶ8�D���˗�V�L�卋���$��,�-:��0>��0$W����eCܫ�io�z�9d|�m����hCJ���B��L���	�P,�_��.Bs���t��kĩ{T��8#*������۰�ZZ�6@���l<�WѠ���Ky����p��}�8�X����~E����"ި�<�y�V�_r)a��zU���bo��4Wb���`CS�=���3=t�KZ��;����n%����W{�n�C���ӹ�2�UA�կw��R�N.i`�������֣Ao˽�߷}��Jl�Ԑ��Xh�p�7�ё�lK$u$Xu-���ϖ�@�>�):C����B�m�C#��,��ՆJ���x�i�HE矛���� G�9G	�&1���#���ݼ��Ǎk,bP�[1_���C_A22�n����ry�e_i�!�e�}N�d��
4G`}�"}���J��������6��mR�Y�m���/�Z���àU�h�rgGY�* �j;m���їL����Yg��*ۡ��-&W��D�\��!N�}�U��s�� 7�h��o����@f�ZC�6\�.�w�h�o����&�4§�W��v��##��
Y�c0t���Z �Ԕ�i%E��PgE@�m�ކ������s�O�⢉��u����O�v�؜k��<���j��:ۉ!���]�����!�F�Zs�L�gW����d��q�BJ���Z>�<-�!����0L��0���b�۪�Z/B�%��|�O������>`�� \�����76�喫'm����������K��y�g�@wF���R�)t�^�5�S�TO	U ���a��Y�m7��R^;-�Ь���T	�Q����zH�Dq��B�]Hc^�"l��f�O�^�Z)�cya�G{¸��B��u�Ĵ���?1�ϑ^	���,2V�C���n� ��.���Mz��sj��=�8���P9sꋾZ���}=�U�q7���%���O�c� �c0�=R{ч����m6t`5���>����:�����u�P���I�2��*�����N�b=����H��v���~rɋpibǗe�v�i�r��Z���b���0�� �yqV�݁S�d�r,d��1m���҄{9ֵ�DZ(���R2�,|\��ڒsc�=�V���dO�w���#dStj���h�&v�_�}Rk� �]W*����ۣ��/�rO�)�E��_�t��P�7����a��,�ݟ%����&Bn�~N7{6?��i9i��;�x�o�ϛy��)���9T���	�[9ۘ�n�Io �@��� v�hZu�_@ j�(�3�j�4O��u���ȥ-7'	���+�}���!���V)��5O�b�{��uV"��~d�3N ���r�z��ί�Q��#����В������X�nx��(e�s�7�%�?��P�IW&�6��;��қ_έ�E:3�=�8�꤬���2�/4_Y���ߧ�����׫D ��}ޠ�A�h+;��t�Ѳ�E�X@�m���	9�1nP�?�L
V=Z�����X����Y����W�u��x�x@Ơj�kft�j�	~y4���z�ex��.]t����(w���&��+Jl�����M�O��]R��q��R�ĭ��7�<���6pV%��������G^5Wf�M��)�ϬT��Y��2C�Da5Z�J@�dP=�z�33���z���2Kmt�m��k�s�B6=?b�����V�Ikc��&%V���3�H���+]��Z����%3���:%H�z�ǘ�{�A�G� Ys�#l#�2^�#ߧA棲���C[�N��j���� �NʃQ�
�����iO'`����T��{�����k�=�g�f��sfx-m*$�`�tn"��/Y��ZWE9�事�PGH�H�x���YP����w�n`Bt����L=�m�F���^��~�HHo'!%��49��($��P:sT�������L�d�͇�͑�݀���PG�̱����+���V����=9��t���+��`R_�R��zs���� �'0�`A)V�[�5��ZTd�Fi���������� ������X��^��|��e�OԱ4�������9tBy��f_j���T��{5��)yma���x���������s}��Y���f��Cp�9/ׅO�U$�������01ƹ�w]E/'Ӆ���ţ�H��U;)�4���b`�
�i���f��|�X�g��PX0X� ���JCم�tb��g�c�-̺g��n%ƌѬ���O���.��t��I����)!���>�k�{��7�h�0�ހjD^�C\��qx8�tA|�5��	���H����#1��F��iɍ_��YQ���A�L�^��`��B_G-e~����5���_�Q'��J(D�m���<��Yߕ̨pk�%����e���uoH��?���`�2���fφFN0�'�Nm:�8.@FP޾�H�wG�I�H��Lꋏ���}�y~�U]3R<66P���J��_���,�f8��J$��H��O��*�K��sL
��u�=���g�5�	���wc?�\s��h�K��4Eь3�"M9��������0�l�{��w�_ T^�t��LM�v<9���')�8C� �I����'e�f���'�|7����/'�WS� 5�P���YA������JU:�^�P:{�T1,�A͝ȒМ�(��$:�o��}��b�O�P|����`�I�<�b$��˕��qEE
��aM��77ш;�H4���)iR��p���S�qf��0��Y��+��W�F�%9�(C�ṫ_�t��ѿ����	��ōή��c�-QW��LR�x�c�ל��f�ƕV���9,V*p�'-��n2��݆�B]�	z	+�f�+�ޣ����b}*�	�=W��Z�=VSR։F��h�U�q��
���K�ߪ^��*(�?��E��{��ĵ9yj�K##"+�.J ~%)ZX(9��:"L��A4�$z6#C~_wwNBy`NK3G[��:p����Az�ii. ���V�͖2�-ZL�7-�R����Ou��}h��sYX�}���s�ˍM�����*�>t���Q'UP�a�\`m\�s��te�PJB@Bش$e�.'�i��t^d��c����\���!�D]w�VL��ޜ,�|���ׄ邗��{�O�h^6�+A
{y���\}]h86��U�h}hD�B�4b}�t`��8�MO�ֶU�������i����t)��R�%��Ғr�{K<K��྄��̦��7����jD�b=V3�9����l�p�2��vF�ЕV�k9wlT�*j���GA��p�ݭ�s
{���p�bX�D`�0K��Lu.�NV��C;�G�����Y�0.�ngM�'�s`|�T��f�V���kgBg�ӛ[�Qw߻�;nP,S:"4�p�6՟������	��<�t��> l���X��zx���ˏ?�˫��߬�$8D&|T��U]h+�R���l��]�>��x�5v~��O{s��|v*�Pws�j@�y,���*s��G�M|���snO�7Xh��ʾ����{�J������y�����[ <B����L���* �J�`.�Ǌ_J�.�����,�>��d��@#��G����Re����0p�@�1$$���h�^����a�U�.'�n�9T>�G�A�GSwi¡q�.���I��$/�? � ��i�����P�x>�S�$�z;�h�x+:_u	���x��������tb
�_�v�G�q�"�8k4P)	����HxUF�m����wO�X1Qb��Y������v���GS�M���ͼߧ���mJG�����i}-�"+|#9�����
�;+`Vn�~�>Z���l�WOn�.?.���u2�������Vɺ�J0�H�N�)"�����;Ds���f��9`�7N?�ЅZZ'�����n��[o� a?h�0�*������h�ޱ�B`�
ޗ�=��t�I���4�M�������k�ۉ-V�=�Dm�+qA��	��W��O�n���0p��K�/��4�������]��� �}_�@��*���1��5l*����Ƃ�&ٯ�f��.����*k_p�@,��ۉ����P�+�g]+,S��V��Q�>�Iqد @k��F�/E�'v�%�u�N�գ����9�c��O��cLf}��������ߞ��9�]���/�Ɠ�{�n�������~Y*������#ɢ�*`�D�㼔�����0��d-�M��Z7;�����ߕ�޼� �?��c��tn�#�>s����l�ވ����엞��Y�7Ȭ}5Ij���_j������D��ٔY����2�0c�޿�N��������|��]�ީX�T��RV-f�������o���#�ϰ�-þ��3�F�G�$�e5�T���?6�������6W\l*���*�C����/����|#��ߏ).{���>�տ췶�~��ҩ��N�ߊ8���3�5�g�e�8l���5a����N��i�Sn�=�ߗ��������+�~�0����=��3���ϰ�m�.����m�����ޙkn��G�r��~S�s�7R@e�^��(��ݭ�W�V��h۟��}��T3��g�E�珋)�8���s�"�mr�]Vd�|3ӇpBrs�)��q(���3o�w͗$9�M��F5=Mj���UG��8��������ًp����rox6��Z��a1�>I�r�I��,�Ň�����F����w�W-W���&��pO�zj���j�Ղ�$P��N�#�Adǒ8���AA��/� fST����g����^���<�ͭ��y����xT[5�S�TE�SϩVklQZsK͢���O����Yh�h�1A�UR51��HB�)��i{�{}}�}�+�p���k��Z���p�=�5�@�ը� u]Ǆ�LW&���t�8Г:�[K�M����$��mi:��ޅ]<��%6{�_��lȵÅ�f]r�	�F�qY	��'p� �.ߏ�~��}��ZC�;�ډ�ۉ�3>2A�n�����]#am���ƹ�O�z�|�.+�P�Jb.ީ��rH���Ύ���:7��Z9���o�o��_j{����	�_4B�gu����Φ>L	l^|��d�}��������>��@'�����p��yz�%'.���[��]���_�k�Y7�d�p��|s�I�XfR��L߷n�"��YꥶE�Ie7��n~9���5v|�e���:�Ӊ��9�7�K�/��O��<���/���#.k!��뻯h|��O�Pp�ܔ,p��喽,ʓ������� }U��s�^8�)����lqs~d��T�?�w~kOK�|�Y��T?�5-��d߼��������ѿ�\�%��
��.����(I!�g�T�W��^�h�e���������VZ�S�K�A�d���]��)X8^�2�,p��xWAA@�&�I*� �VzA5_�ۣϾ��"l�L6��T�oW^}Ex{l\;dg 6m�#�nO�s{��eZ~_�z}sƓ�A3�99��C��HF�S�u\��|�]r���﴿�h�$I����g�wc�m_�°f��-�eT����vR��>�_��ƈKm�oH�CS
�b�vssË}��3T��<�j�����[�@�Z|3�T\_�������f�� ���=9��Q�	�/�WB�D���́[)f�\�q�]�Y ��^�}�S�����)�Ņ�6(|���%��ϡ�߈+^ߦ�[������/��������%�V����@�ا�jt��>yr�V��$Ss�RUk����m��G3�Tm�ۇ�U�J�>����%DN"d͢?���KY��֟�s�FS�'59JSDX�<��C=�C����ӂYYZ+��И��	u�����E�A�o1�d��'="�������w����?Z������T���E��*�փ���K�Pw(��5'��]D�sq��k���"��]}iq�d��Q��k"��5��lB$G'��k��؞��F���fA���ڵ���OgT�?yr�l�=Ҧ����$NR"[��@ou����}����z3�z5�,�U���}���\�n����Jq��I@�tW��Ї��B���?�+Gy;z�7�+�Ԭ{m��cj��@wm���@������`���FbRO��Lμ=x#2+*�㇟���Y��&��Oٵ��͠~Zq�jt��уS��f��=~IS��A�/�=�}�H���hE����M�(�C�'������ٷL�� iZ�F!��[[��jo��e����j��Y飊dղ	W.)�?�������_�dYA�`�Sc�Uo(��m��qO�,�ig��3z�z��/V��m��TZZ�4?���9�U���$mhB\%wHD��%b��{<8�m�\բ'�w�tlpr)�3�����<�01q����~I�"���������%�v�τ��1Et���}W˺��?!s�����07�di3O��_��W���`j�f"ȃ���	�
�26�x���ʒ:z�;���4|�N}Ig"�=7��Y{^���+����_Ԉ�KU��9�X����.8����T�t��r�c���R%,�P)���@�5�Ώ
���m
��TM�uɹvpZ]�� ��⭍{Y�$��waV0`)	���ƒ�:X�Z�sC��s�hO��fF���u^}�=�6���R�I���¿ݤ��ǍU�������b�=9t�J=�v8HQ�B���O
��q�E���=�[ex���>�Ao��t1|��J�5G'l���]?���I���$u�����������������v�>x�@[���&[܂ֿ�9��mM����v�����9i�u�u薆�E=����~)���3�O3�!�hǱ{��䛥v6��z������%�%�����	�Ծ�t��n��E��>U���`W�p'�IuX�$a,U��)t�Č��Dg�����w�����=�P!K�U��$�M���F�Dy������>��=�S�I��k�c�S���p  ��#�oe��0a�	#L�������@�ܸ��hJ��/GН���c9 ��5@ôxH�<���8 �H����C�K�x���ֱK=]��'5+?^��џ���w����������DS��ScfD$�|��������;m�^n�aǋ�K4�?}�<�/���һa�3�Y�qs4w����⇒4�>���n�i�	A���zv����ծf�?����Y���W�x�6ɢbs��&7�B�V��A�oĀ�������Ɵ�Q��u����$ã��;�Uh�%��T�!
is(,@|��M'���ß�酐��"�D��� �7�y�\�3���J!�&w����Qu��í���Wy�v��'�!�y%����#�̴�X��c����>��p�����^}Y#D)�]����	?eR^&^ff���N�����6G��'�Oo��î9$�Y���ݹ��8��;\-���[%��ݳ6H}���a��Z\�18�^.��D3�lDP���Cr���ZkiE�sm�n������+}�䉹��1�~��0�����92������ <˾�&������ -D�7k%Z��L�#�E�����w�Xo��0�Ω�
=k�q��_1j8���D��+f�v{5��5ٯ�{\( �4��7�/\9����8�l������_����(�"#ü��EH�ϸ�<�V=<%PB)}D��,�$q��x�[Tm�)�%�mb��%S�Grm�%w}"W�v��ҙ*a��惘DB4w�CN�|����bSf�Q��b|�1�:m�X�|��n���יU��A*�w�*ujT�<S���ZZ#���=tu��*e�7C��hR0�Nx�4��&��e]y�x�.�f�Xӌ�<V~2f����3�O�Z,��-ֶ���L�6r�~1�m�m�}��s�暓0�w��M���ɾ��,�@*��b�2c�@[l�>Y�`��g�'B��rX�Ȣ���)�����/��3����c����/�kY�m�5�{"�-��>�Rf&�U	��GA���2�^��c��E.dw2uqL�B���T�E��hN�_3��V�k����[�e��ڣ;��Н��&�ٝ8���Z��l�ަj��JqFxt_~�ְ �����#o��&�c���v[f����s���1J�+�X��Œ>�SGrrl�~G�u;�Ʃ���D0����cE*���B=ټ�����!�C�X,g#�pawC���fs�v�/�m˄��0�� !ם֩V����\�;�a;��67�§�;һ�^G���'�a�,����t��n(�}��ճfN��#�,\��Er�VT
Yf���d)��O2�d�VM,c@��;T�Qe�f)ə8�2@�IJ����۔�*�N��8�;6�ؽ�'e���.	}�Tx#'��?�b�c�mx�|Al�����,�	}��"Zى�x\`���O�9���`C����������F�=��5��� )
������:����N��4��fcw�>�;6��39��Xw�J�����2�yy��H>�
�v�?�f0�W���������g���]�����f��3_P�1t�+ d���	�dk0ʁlf����"�V�L��~5�{�Q�ߘ�̼c��.�
#�D�_ˉ@j~��^l��j�����'�儢�5��^��$��-uc\�g�r�]����Y����M������P�u.��Z�����{���-�4n�֝e�ٙWtN��\��杢�9*�]�ӣЧ���ۮ�ƹׂ�w{,8{5�"efHh؇Ң2��0ـS��ݹ$�n�^��Z�N�H��
_j��l�XTk9��[{qKA��R�&OfN�[<WL�޲���r�+�O�1j�j��S���9l���S�m�����D��:�ݿSu��`~�&'��=ͅ,m�l�DC��FqOn%YS7�[V��p��x]��1���>�;�jԗ�;����Ѥ6�1��kUz1���qqCJNH%ǚ��\GK�	�������\�A��^�ugM 	M�����e9�˖�=XPM-�x���2��n>�������:b�H��5���2��՘��Y(�xԟ��:T 9D�*z�mt��+i�X��\uI�� z��ǵ8S�L@�'�btfek}"���ev>���XQ��ؙ�'�.$vDe����d��%��GJ
<%�A{Ĉ�I=��s�c��Ow�A�9��U&/0��CL>�,Y/$,�\���<3ݮ.�u�����?� [ u�&]װ;g��;�-��*�-sQ^�$���W�oHƬ�3�q�A��.�y�_�cD��S̘�U� �Ͳ�"LT��26���j`����\��TT�n�}���W��g��F3�d�W���pT��l{����I�OOhwM@D=K/0'���)�0J�4P�S�W!}�K�)Q!f��NBvO��<M�u|;�z|�nb�B��v��ޠ�m��{�D���y���߿��h,��?��Ν\�սy��Rh�t|������,U�������S08~�[�1�ԯ͐���?�e�x��.�̼_�'B��H���j�話��wm��4�WoG�v~"<�Wt�r4j�e��wU�Wq���ew�֗��-t� ���	��Ӂx��o�'L�j����<�J���yIN���{^��n�h���qK�"E#�I#n�(��N�Yq��ZGE���¢W_��n�y6��&QXO�q ���O�����*#uZ3�^T���wG����b趖ჱҐ�%��/#.Z����{x#��pb����kƧ����ݼ&f웋�Ђ��ϖE��|������3!��'����_Ϳ��L�;C�Ԍ�1�=z��t��>��Q�eN��͢����g�*Zգ��1L�ϸ:'\o��/,��ll��b��DN\i�0Ox8��	�H�[[�3!=% ��#ѫ��^�-(�Fߜ�Cki�B�o��I�E����u��x�E62VN��%r��Au���u�;����L���2�3L�����r��TV$!�Ϻc����0O������{رp��v�ʭ/��M\�
���;�V��O$�Tm$��Y8af��t��h�'<"(�M B�M43u��d�`�Ma��R��j��w�<�u��G�=(I��셵?K_n@�v�;ʉ�W�D�j�|b�ݖ���.
j�:�A�S{�����N�o��q�q��*`��h����RJJ.A�u]�hB����z�f.d�s��ctl����z�3l��a����Փ���eO�'��d�@�Z��3
PT*A����f���e��:\z�$�DEAQ��WM�>�O<��Cfm�wU
Z����5��Jm~<3O�bt���$�N�o��6n��6��0��k'V⶯H�*��9XW�2��g�y��+&@�F�%�0�i�e-��R�]o�?��&вB�e`(M�m[*�w�p�涎=Nlfp���dt�.ݶ*��p���ԉ�ӆ�@:����4$��tL��R��!�q�,x���d��ڌ|�d:��`�5y29����5qq�5��!�Yd�7{�v	b+�K�|�v�c����FTZ�m�#a�4�/_�e� �/#�v����a�P�ѕ&t��l���J�K��!j���~���k�������5w����<�8��`��� �	!vyA��,�d�.�N�~=J~NS������dr��H̺b㥟��p�?��Z�|��{Qݕp�bRmbo�+����~��+�B�����M=��Q�.w��8�T�y��_b=�ۋTer;� yC��h!(V��f��qW�'��[K(R�"Y/g�8o!s�'5��Ѵ�(9<D�1ƞ�%��,g�Ɛ�F��~ff�K�z5�����S+��>�~J~��x�3���T���R<�Ee��G
5�n}
bo�.���nFq3
��[����<�c���&���a<(ry7Ztx��y���u�nl��-ѷͿ��
[���ʟ����-��4���̱%�T�*��%�f�y�(�$�/�a�u�]������Pza�#���~m���{�}vV�#��\�_x�:f)��f�L=�0e��nKD����|0�js:ٌ4p6C��ֆ�R-��^��Z�fyGQ���J���jf�F�kQxC�Aʓ�/�8F9Ue{l?��N�����`��_���;WM4D?+ׅ	d�,��2�=[�fr���� �U���~;ZE��%���)4?��V9��)��.1+w��8B�WHk���=��T��Ly
>Ez�N�r�F5�W�������H̥8�"L+�Y:z�Cjnxv��ȷ��1En̒K��r�+����2Y���ȫ��ayM��a�mwXޚM{�-�`b�`�c���2Эz?� �"���I/j�_�L+�u��f\�^�T�Y��������0�|W1$B�=�HA��6��TB��J"�١Ö@KI��	x�L���Ή������"��A��'t�W��2*v���IS�����K�߁A�]�b	\F���Q1��q���e{��8���:�'���c�x�g�� OZK�$�Pc�r3��2j�M�%Q�Nt�Ԑ���VO�^�j�Y!Vr�(@�7�5�����[f*���
�����������m��#�u)�̷-*��R\,� �-/a��h!6�jR.%�9��q�³gVC�b��[�za�]^=V��|��a���D7�~#)�v�>g.W��cl.��x�lCﲣ��k�<�1�J����i�G����/�{8�E�>�S�l\G�y�p�G�6�S��?:�����O��C?49��}��1�~�f$�AZ�c�{3U�r�iu|k��qc�(%=�5����v���S@�l�'��PK-Zk�#˳��fc�n��+�)�FN�I��:��3W�n�z����E��_�'Z�z	e���i^﫡L�N?��M��P3H�VRUM�؍�%Ǳe�r��+H�k�N��˰��#FO1���-�?���jo���}��:_�S�^���:xC�_Oج:�]�ٓ��g��r��,�N��^\ꞥDН��a����>�D�N�/Y��mG(�t���nnf_̧���堈6�娲�����F�U�ҞODVI	"=����W��NO7�t���;M&����l� �󁠤w���C*E�{8n�]��Gd��ΡWA]�zT���a����+6MCm5�8k.�W�?��_�~+���*���ǆw��J�������\'?�":�fz՚�pv�*5���#�FZ	�.a��4	��gR��v3	+���t�}\�st$U0�>nWC��NR��ݶ��(��Y`3H��&�Q~��P�q��C�]+<6� j���3�#�Ez�'����#����~>�=ȃ]�ż]lB΃@f���<0��ք����K�C�W�<+�_v�b�ؠ(e� �Vt�0�_"]"�߅}-�[�[l��zڱR��IG�m���H�Mqï���Ս�I=���K�W�1�fF2R���-E�p�g�Q���xP�ɘ����Vɇ1���3�on�s�������g{�p:������pe�`#]�p�������DT]��)2���L��WQnE���w�Hc.
֕� J
�ftn�º+|6���� e^��qX�9lq6����F.�Ojh>�I�KU[��u�h���ӭ��ۄ�g��q�Q����Λ-= m@�eη�\j��w#�C��nTx��>��T!��Pԛ�Y6��_RD����^�bH�p_�7�1�O���(��q������_�H������\Ō�Fz`~+z�Y�֔�ȣ���-@���*��]q~���<����߭4j�m�w�Q���V��pr�S���߃�� ��<�i�Y3k�='L�X$d�{o�Dy�݈5���cI dmȷq�2J��"_&�P��@1.T���[f�ܵ�������a�G/�M�BZ�C�q/�r��,��[�qyǂf�*77;��{�`�tH.��`ڧŃϓ���_�8�P�zY�B'�6J��5��M�J�A�^Oʋ������(�G���J�Nt����k��U��V�����(w6�Պ�z�w5SQ��h�I�hV��1�p�d~7;�<�_�du7�+ �,������uI�?�z����������Yt�c"l"'WS�ϝ8H5늘�	���HN6x���dV������-�{� {�pv6%����8kt�p7� e5�W��?��z�
�������v�������P��2�2[�TA92��r!�p8ć
G>���#=��_������OZ��}��~)l?;��|y����a���u����(�q��K�ȵ/��,A� ߙve�'@E�{dۿ��4��&4��SSM���ZZ^�w!%WL�;������؝" u�$�H9����햘;�
�!4�eȚ�3S!?�<t�ti8IF����`]:�>	�3��ǖ7l�f�t\��4��~��N����w�r��c����_�x#u�_����ɳZ��I��b��ꄖ���vba%�Xk�����tu�J	�-�h�٬ow�7j���o�qCah����)�H�<�]�Ш~oCU�z�9�o�$TQ���C�;�\�(L��%�ǖ񏤽�i7� _~�_��y�R�cW(�b4�x�;<��� �:�����=��Tk�>� ��/�F�wh��[��6�81��+�5X�H�h�u�I�Ѻ�So����Yg����V��!VkK��)��~��� ?�ƣ~�� :���%��>%-�+�P�-a���0��	��G���J��_�SG��l����'0~�R]�(u@m��9{��EN<���������؝���ME������Y�Cm�_HB���"V�I)����_,����<�lR`c�P�~KW���H�*$*�f��_� �+�{NqWJb���xf*�����y6~�)��i��`AЅ���\y�"zQ�# \#�,I��Wچ�Ӯ�����&�Rq�˼K�oU��Z����:oFZ��\�@�|-�k�b�`��MtFE��Y�K���Oriƿ�o;�G	NN5�y|*Y��/�p���7EF�	�Ǟ�=�$~�lYBm�_�\G2
�p�<�mnϮ,����St|6�s*@k�����{�Wbw��[F�Z7\�L�*�^PNg��.���F�� �E�:�e��A���2z�D�di� ��a���rlde�:�J#��h���"Zcy���P*�4Bi@f�����J?���Ķ�bBCw4�G��/���f�6ڧ���$/�N�J���Y$K�Ѥ1�_��O�U��;ן�k�e�����iD�|E��J�BJ���*�����[�T����>u�ii�0xmR��A=܁��<����s?4�TA��D����c�X�Q[xr�VUl�h��"��]?k�kM�aC
�}(�V�J=̚(^]�/$�R����C�6�Ԛ/Q��i��Y��{Є�!���ΊC1:9H�>�����!l���n����Q�<\:���)����*�U�+�����������6&ix��9(����qC+L�΍�Uc@8s%�T2v0�7�A˩���̹����`��*V��Л+��VT����^���0��.٘��,0�P�4F��q�ИF���O��S\�/ږ��L8�V�Q�9�/� .���rnqo��
T��e1	"��Y��_<�n#�[k]�>.��>vV�'���O� ��&���-j�|�Ρ��5� �@�Re!�z��+`�*[7� (�ӄ�Uۏ����JrۆL�@�oR�}��P���#�_��Qб|�X @�>�;$uW�¶\�&uw�0�q��9��\]N�K�⎸�A����87����� �X� ����z�t��zS�D�k�F��_�PNe
i�g�e^{]�Aʽ��0,:�|�ʌ���3�h_v��]�ê���6Sd�)�̵.�P�y���sIy�\�1�x����A`�a���!���>'��4r
bЖ��>S-�}��H#��ز�z^�?^\���q����C����o�}m��ʃ�џ�.��W�[[��,Z ����V�p�+������Қϗ�Z]W�=�,��_��:>�v��0c��q�SL,��G�q��5�YdE�O�����|F�D7n~�P�5�W5R���=�9 ��G��+Ud�LT�? �{xp�q����HQ�m���{-�`���s/���SJ�}E����g����>���,�7Ԥץr��#4�-�����|�j���sL���GO��f����󸨭f��f����ك��ґ�JM���vs���ʜ4�Cf5��Kп�"�)���@��i�*��(;"[�(�S*��L7�ۋ��.����e���@��e�y�� �^��hU`"�1�����	&�&ڣ����/�Fq��M�)�׺��ҥ�ʉ�;����om}ǆ�e̓���j�ϴ�G�����2���x��k��L�-���T6� �����<O-�|lYr�+�'��9�]�R� `���Bf�*��!ߣ?��
�wy��{&&d���\���o�Yp���bFֵ4�)����zs9�a��Ȋ {�c@�{m�~4�,�{!�ρ�g��x��A�8���ep����'swyr�&E����-�@�[J��B�^�V5p����5	���UB��G�!7\�]��5ֳ�|�@�GY�J9�y@�K�1^<I~�y��36qSS���%Wb3� �� "�1Dn�����ח��J��D�w���^'�N!ڢg�K�k�&7e��o�풫��9���)�R! ���{�E�yQ���Si�='6��i[tͼ��H��K@��K�m?rEma��}'��,/G@�࿖�p��N{�<���i�SX+({I]��3�s�H��e��G�/f�W���H���xN��y�G�^D��Pv�z��$}#������h"����j���c �8:����k���Z��|�]@=��K����%�����`��N�/~(O�Qt�3�R�Yo[\ʲ�![�B��:��d�83�Y�4��T���LZ�et���@����� 2��kw�oq�0,J���g	�0��u0�0���^�i�˂�*,����+���H��4	��ACz�v��X�ir�?�?��ȓ�F`|H�g��?�{q�{��G�b��;E7�^m���:����G�
�4�/(ؑwN�f�^�f�w��cU����y�ds��G7���ݏtԞ�N���WSi�p�z�r'��J���t�+?7��M{�#��h�ս��s��`���=r���z-H+Q�2b�~p�*��{�����L�?w��.q��.g1�A
���p��*['�]ȓ>`}�.&��7
��@2��4���8����쯐���#����M��z{qhI��Q��lL��"B3����t��:�ʝ�G�
Ƈ�-���LF��kDq���lD`SiA��f���~��������;��}�лY��zj���^�%:��F����z6fBV�ٜ��t%�W�[����	� ������J�!b�/���������6m!���N�=� �� �{^&�v��� d��QP���%�	Ɠ��%o�ςS
��؝�����������JK�edyY�GZ�j�XiS'v�̣p<��=����>�tA�'��a��E@�~ځy��4���>a)���b��+vB���p��3�T�W��E��Wm��:6p�n�+�t1'Ux����"�����&#��9���v�ٕ?3���N<)� 6j�)��?�-�o�
��|��N[�G�����!��4�D'OS�"�t1�{�D�S��Ʃ�B](�xf�г�X����H�q���\/��m��D|#╉ޖ����N6��`�!�.>�/c�S4+D���RXA���;ςYd�7��X�a��_;�=�h�3�[)a���_%F;k�fL5���j���;�~i1_������<�=��#����gv����/$�@q���κN��@f�63_g��L�@��|����C�.��IX�n7��蔢��j�t�h��`<�!����������՜�;�.��x�2
�0��\h�c*�zw�h���p��\b)�~q��4�z����VW�^���ȅ��'m�MF�{�hi^��b?J��ڝ�u@�w��3�}}0��	3�T�m�g�ڨ�֞8�p�3z;�����xS8Y��2�w��0�a�oN����p�Ei�����Y����ɨ�1�e`��m�>"ec���}52��_�\�z�Pu(/�Uک=Q�o��]$H�Gw�s}�x9��<�I�j�w6��犢�Gp�3T����.��㹘���EZ4]gY�� :d2�{��j�n�~������޵v�;��@����.�ğ�S8d+/I"�Q	R�C�!��w���H���CX���f�^��ۏ��+�vI�3�ND+��t�kj�N\3Y�K�����v��0�/i�4����AK���8H-�d��@���Y�e�g�]m�m9��б��D�?S�M�<�
u�~�a��H���<�R
5׾��i�C�褵R�*��F�n��3e������r��Dۗ�R�ʐY�*�}>�)}jL��S��Y���Ԡ�@w���u��'�-OR͛2�H��@n����(f�d�L fƫ�5C,qN��5�ng<�W�*1 ��L٬�'/��-�ႇ6`���j���������Z�&�!~�~H�C/��x���w˞e͈{����/%�>͠�OzY!���R#CЎ.2�{�5b���J�9�X�ny�b��.�eu1��M��~-e4<j7W	e�i�[oK"T���P@��ý�X�r!��nM�h9�����KY��?��L�f�CKߛ�z;��������[ߦ�J���Fr���.�z�	����m=�#��v���Ȍ�m����k���y1����9u��V ���zr�-�G�tג�X�Vʍ�0�A����]��^�
)�?�蕧[�_hVwH/���
..4,��ڳ�A��{iz!۩�Gz�![Ť��c����{k�`a�M�hZy�t�<nu(d�UC�����p}�g�ُݵ�'�ζ���z���9v́w_��R3�]�$�Pj��3�������пR��{@Rz0��E�����xb�ӎ��y:S��j��% -[_Թ�ޗ�UBu1�y�t$�ݷ���� ��z<<5v(ǛN�f�ڔ����O���z�Z���P��uO��M˃�L��ol\	S��z��f�����[N2ʫ�����J�R�U��y������- <S��/�a�153qH=��v{�ͶBݦ��j-��	 ��b�&#EX�R���T����'�O�*�y
�W��g�	�y�\X[�|�(ң~FIUYF�9"M%s6%���KT��W�*�
`��-
�%��lci�X�܌���:��C1]|z�����J�$`��W�]8S�vkx��Z�s���u��$Y�(`+I�!�����T��1C��f�"Q�Fu^�6�Y.��y3�1� ����Ol����HZA֫(�D	�d�L�%��p�f���$�\�]��[V�W ��+6�&&4��+@1~�Z��z-O{>@p�s��VK�v����y@�_��zַ���6B&��TV��焔��Ho{�G��%JU`Uٰ� �̙^n�(�-�s��/]�J)����=�Oq}��A��7�<3�8��rO�HaPް��&�H #zM�Ғ�%1����c�e�=ڋr���x �^�a�w�ә��j�`3�N��PK����0�{K�E����"�(�F|��t	��λ������,�H����"�&KeI�%��`�Ab'�xdL=Su�V�G	4B����:i����GIU0��-�W'Ҵ�SQ&��
hֽNhF�J�@�;��ktR��k$�����Z�0~n���36����sB���Һ&Cz��t�i_U�h�\Ph���A�C`�<�V�Ԇ��{�l�qM21�~n�Dn"h 7���6x�i�NШ����a�$3?����H\�	Q���$=Q Y�A'%��h��u�h���{7K�8Ԓ� ��T\��S3���r����� �gÊ ���U:�����}�i�$�Bl��{���ֽ2z�
vA(�6��/w����E5v#�չ#E�����Hu�K�H�"_ix���[_6�nN1���6PU;e$1�z0!��x�9��$��b��}�/�m�n��/�M�<
��Q���B��ϝ�}X���i�\r�^���V?�7pJ��5x&���F?��ʘk����W�j�/��߉lH�a_L 2a����>m��*1�jN�m~��z5���;��0o����ԍ�o
[��;�*��#�Y��a�o�"/�����oQ_�i"�x:GRGf��V�����4���ɒh��zc�A㺎�����ڣ��f�ߎv�y���~Ot��]�:(YE�D�9�AZ����ᾡ�?������q+01SRd�L���}�N j��ro2��^�G�qX����]�z�1czŻ�Ti��Zr��F���vF8~�/�5F�cJXF�E�1`��4F��<�{�06 �e��E�O�&��o�ɢ`��ř(|�GV=�@���+������P�)
ڹTtL�X��^+IU�裷�ĥ� -Q�m%^�����P3���~	QO0G�h��~��N��9u>9����e*sc��f�H��[\LZ1�$*Ze){k���&��W��8㤚"y� �0��h�)�H:�cV�DP���4�.���w��x;�=��]����=x;��RA�?�i���;8�!fp�������'M
4F�/.�i{�+�����T/�I�� ���7��Ց]���kc�w�;���?i�\M�5�W՞������q�����f�=�X��nV+j�1�F+�d�B��Jco����9�����v�vx���2��� Q�`��=V���ܻ�5�G[9���b�ƀ����p��9��a@ּ( =���v�e/��l��6rZ��4%��J�3JK��V�A�Am�RV��S�ɇ�˜���a��g[���_]�6�f^��|�b�a:���v/�`=�c&J.��9SC}����(q/�6�ꠜ�R����a.D]C܄d���c��I�8R9�P���Pl/������C���@��.��[���H6�$ݲ2������%H_0,�Ŏ��GɉxY"�w
��9�@�s�j�k�C����̘����>z*ūξ,��y��j�G�ι1���]}[ߺp����s3�v��t���^���������w�ؖ���NN��'(|^��<p˃�f��F)�т�+l���)r�
c�����6���Ț���[+�y�J�m�\i�����]Wf�M�ׂ��vJ�(%V��{�Vrs�M� ��v��dm�m�0*+w¨���ˤ�����8H�����Ҟ~f��7Y�Ǐk�����^��-Rފ��%�VhJ�v�{�{\N+K��1��_Jv����p� ���Q�c[�toA#z�b{d$�wi�>�Y����z�.�G�3:zil���O��X+�&�Rtu����Py5��E��F���4���ww��}��K�X�z�щ��O~��d�R�rY5)�>�A_W�����R�Y��<�a�E��:Y��zsuh�şl,q�`I����T���b�7�ʖ�=���A��n+� �h{����>B�푄�y����*r�_�
��Es�F���^����y��ɺ7-��>[�Q���Յ�]&�f����6�ѽ��̄�Pf¨������S��d.���,i�j����f$��A�<�6'v�*�㇢v��D�F���)aV$C��&���QqV+���_R�:j.hyN)h9C�=��W|�����Q�U�	���W@�璞ROe�J���X�����+{���ґ��_p���\�1�̝�W9�
+Ujp�.�����9�1��;ڵ�ԁKu���y�o93�Y7��:ܘ�<W}�Ē(+��n�Å�wIl���OE�Vi�^�b|������ܜ�Įy��΍N���A�_Tk�*����bV�R��Ƒ&H�bɗ1屒�1ԉ�#��d�i�W����xmף�(��I�]ܖ6t�s%���T[�h�U�����[|�����ֶ���c����ɛ��~A��hVt�\�er3hl%�LK@��e'��;�P%���C5�@��p�x��'��;�]7*����X�$u�����/3��˦��~�t���y�m(��l��d�H%�M1�k"#�+�o��f1c�Ƒ\�1L�|.��Ws��]j'�K��"�u��{<30�8_���;��z�ݮ����q�"8���QT�K�>�)S�a랆�̾�~ZM�0lTi�AC3�$���\�Q�seWK�L+���ԙ�e�Ɏ��96}�!�ڐ?�F��{$���~��@�(Q{��z>�ꮊ��f���?d���x(�\����F��fdg�)��9�RF�z�mv��5�d��c+��1%x	�}����2������^�S<��?=/-��K_Mk����Ύ���M�z���V`|zBZbxse��ٗW��^ҷ&T���HĉW
[��[,xTG��0�:��!_]�Ç��WDU�UN��@Ȋ�P��>���z!��z�b[�l��� "����v~^��z���0	�ʤ���ƺ�ݻܺ��Uߡ`cc�\n���/�Nr�z�o%Œp�h�Ou<��w��w�>씽R�͗�r�lw�D~�HT�
�!F=>q������N/5&����+��`1�Ȋ���V�Ni9(է���2L�v�f{���;�����q���
RGP�bA�"(]Z("�CB�0"HS� �I�t��PBI��@����n��������keɊ����g�}�{��t��d�j枣�i�V����&��O�\���+��+D�C��,��^ee/�Ra ��>D�I)ڌ����D��/R�lqr6�\����[����&ꚶ�Z�a��V�� ��و{%=�b��Z�'Gz#ON\�s+c���UyC��w7#e����baE����P�N��_�ߡ|3l��E��:NBmH�7���:���/�?z�{<J��k=�yw]܍9y�P�,J�5���?P�'��3 �i^��{��Si���9{X�@S+�4k��t�Fڑ�/������lEQ��������cIeQZ���*�\��Q�v\�x��
q�^!���;j�yz<8o�"��N>S(��r�|E�m�C�����J�X1�����e� �ܥ�4G_�w7s۩kG�F%H)pW�j�ޮ����&��>�x��J(�li�?��?Í�)����!��L[o.r�yG�����.�&������I������5���K��y�|��?a�.����몘q1J`��M�J�n>Ӳ�Q��B�Qm���G���d/�Q�(�!1i�O�X⢒/�s��VQ��E��K�(����/��X$��g���]}x��V�og�kF/���]>�P��u]n��W��P�� ��f���qn?u�>�.j�ʹ��(3�8)I����'��� @���XD/5[f�e���W+Jt�cJL.��W������䣸��O�xY��ᦥ��a.�y��P��Z���\k��J�>[���!{y�r��EU���s�u�~���u?[T��,
�Q�*��ل��h�����9�nϚJqf`��P0��>�!��@���9C�>H9�`V����)��4V4猤w�uF�Ĭ��<X��D]�U��vs<���7�GA��*�}r�C'�����c�%�4��C5��ӱ�=�se��.j�I�e�PS��!z�RF�t���,Hg�i96�W������i�$�Ѷ���:^����XdGh��=v��"���w��t�K�ш2��T�)1
Y��F���{�ܼ��H��3��
�Q�1��}���`�k�u�|��4B���"�K����L�N���<�ȁZn��f�pD�;U��õ�-�!:��Vݗh��?pr�ߟ�Y\�$*���w>P*���NQ�1�_��1�q촁�)DD�p�6��<=^o�`�:���@���ݿ-����`|Z�fG���s:�4��� �i+q�,��S��V�!}Z�����}h�i4�x�&�l��K`�^�5.tH��ѡ��}���k_tb^���;�y��ie��8NL:�wL6(��֍��ҀTs��R<F��.#iN����X���q8+���������w��i��?��*�[�}PR��q��g�������
���̃zs�'��Z4�z�w�_�@H!je���A	e�J�탇��ɻ��G�L����S�1��Z���$'3f���L	-��9��c#�����n��.z4f�q�G��6�����"c?5đ7�5��Ke�;ṉ����u��U�Z5�H��27�9���,�����J��@������J����×y�xL�����]���vr,�.{cR��渂��ī �^�tP6�	��KY��὇�	`f�h�(�f�[s��M]�yFy�f�V��"z�$ZS�^e2Ҏ�����2>y�0�Z�ir�x�n|�]�}��#���sg3��둲�Ϊ�!K�����MZ�)�1f�[R{is�IPCPw6���J����f���!���<I�ؙ��GƇg�? p�q>��_kt�\<��]L��q�~s}B��KİF�ȱ��������F=���K)�ŏ�l����p����u��vW����R�?���3fGn�i��S��G���ڵ����|� S�*�P��A��U�~��D�l-"�d��� 
S�X��~�_���pN�������2J_��;Q4H�u�W�/��}�<�kP��N���kd�Ol�Q�m�\X�.�b�x�����͵7Fܗ��)����,dʹ����X9�%ݗ$�c���v����Y�����`�wJDw��;*���S��3'��
���d��Eg����߄g�|�b6侣�!���'W���8��A&]���##�4k��ٟ��6.Au��H����l[���+�<�@�Q����^��F(Ezb��^��d3�X
D��7i�!�7�+M��'��/y��B)>�z�<1j,��p�A5�p�I)���勿�����[u�u��BϏ׸�\� �Zף�����8ZWv&�'�g_w=3�?�����B�tu+@ �����2��U�ox3S=���d �4��0��=�2m͐Z�V���嵲)�1��t��.>����ס�Q�܍��������N�,�⏦n�S%��(Z�����Vv/za3�����q~2�I��J{�9"8�`I�0z�[r�}e*��R�f��'�'/a�o~�i��z\�\��tM꽪�\s�x�h�� ����2Pk�K+�K1�ܞЬ)�Va�Prk�k�]#��	��Y�)i�$�jJ������`�i��J�c�^"�8����זi]��I�la�T~w���н/`�W�f����U�^��� �7�׽/� &7��I���i�^V���k�U��m�j��!6i����71�?�5�Ѿ�W,��i��8��Nm�ں�w9;ưA����������[ d>{�c�5��8�m0�A��Kz�'�����tլ/sqG�J}�n���@��m�ɣ�C��ۇ��؛�_u�Wd|.]z��=$Ӕ-��q�r�%Π� �z�8ݒF�[��I��uh���V��	�q(+��;e�hȈ�:d�:��wI3��g	ʷ_u�[)C��a�"�v�s,G? !_���z���9�^�zUL���.����O^�0`�l��ܞ� \�BX:��̬�ѠO�h�ͲI��eR��p�5R�DU�	�d���:��#SNC�����,q�*?f:\c���n��w����_<�Zd���] �Ru�@�ߺ�ӵ�������r�>13��Ǯ@����p���њ���N�'��b����z���'�����i�JP.��̨����5;��H�I}P�����{�Jځ���t-�ı��3tM���]�;���F
r��ݍ �.ǘ�uՉ�D�"��s�c^3kO��6���a:�n�>(�9�JR�t���N�Q%U��Co�h*����n�Lrܨ���@�K��3�X����ҫ��<�;���}�%�S�$�������]!�/���}D�b�j�e�+�Q]Om4ǟl�O��0�?b�����س�49�\�l�ޒ�?\]���:��������ջ��^oVn4+`�B����ȷ��z�Xc��_�K
�K��^����f�j�X,ME`��%��	�:�)q����4mᵧ��G�����W~�՛���"\jZ�����o,9��*��`S߆
�Mf"F��O�b������zL��ͨ�*���/��]���Wb��}�W%V���, �ߕX9�) ���A9�K�N5�ĵ�O�a�ٌC�51,�Z���1%JZb;F-��S��	�˼�� GF�\��g9�|����ËΜY:�y=L/�6�{?�\��=~�������<ﭜvñ���
ïUU��~u��*�NT���ri;������/b������P���ZV� � �[�O��>jN;�P�Ȕ2�����(#/�o�$q`{3|o�#26 >��ma�	N%���Y�(䫋�ah@�c�+V�\�gb�����o�_��j��?~T��	����?�/�6�6�]�o���9���@yo�oh��CQ�G�@lt8��ȑ���A���ʹ�Ъ��X�`:��9�}W(+�Q��$�>������ͱ!�:�6`<���e���_i��s�?ڀ}�@�|�$�?jF��V䮑����,����S)���r�?��Jw'��U�U����Q���8W�N��&�X�G�ư��m��C}*#�K8�ssV����jUf���fc�a�-!�Ce�;DGJ"Y'vW���.�rhX�������^���?��A	�{A�厾T�
�O�����u��όK.%��<)!��yZG,b�h��у�����f!\hZҖ+ХV��(�h�w�"c�M_�aw}�CUT	�2���F_Z�.��ӌƽ�yČCE��R�w�"�_vm��'��g>��E�/�}�o<��Y�A�!����Z�/?��hf�`�:�<���| ���Ŕ<�iоC_S����OT0 9[�����Ip�\��*˹a@��� \@k(�{|:�:	ޢ� ��۰��{�=��dasQO�~	����p��0+��P�22��5�7@��g���{������O� �^�Zyp��0��L���?�,#��*?� e�S�,sW"[�,9Rf{�=d]����u'��fݿQz��l������p){>e�X˥6o�E',i�6��(XL-�W#�x���zŔ�P}�]�6(�޳}�n���W4o2��\��ֺH��WRc��m��$ ���Q
MK2�%|\8eտQ�}�)Q1���zԵ�2�>�8��j��z��^1}�����2�eʹ�7�.�qڟ��M���dյm��� u�)�����a�M�������=����_7�b+JWh�:���r�W�uP���7U�w����� CUV�� WTu�愈w����	���ܟ�N^t��c����s_�P{1I��~�_���<)i��6�7ȧ�{��h)�x�U/5���?�������1w�����n�߭������������֓l�O�C�K�Y�:�!
ލ3�zqzEg1^	�������x/ �v���x��g��f���N�{+3M��vj��d��o3ٲ1�W8��ǆ�$+[O\�/G���2NW��\UK>ET��C7���?2?��0,l���Ľ�8�w�(*Ų��vW��5�W��M�/�¢~�ňdۧ��D�o��$�G[&=̔��h!�-1o;ۗ����aˮ��&�k��Qs{�V�`�O��p��Ɵ������;��#�9����t�����W@�/��owH~�p�x��5��%v%�3zg���A�6Q�SZ&t�����qWY�[9��W��Ų���B.ގ==n�������)L:&��Q�����h�z»�h;Qּ�����;W�a��m�QD�T������S,֦f�����%(ne�*?��a��D�\�my@2Y��\#�,�lu�������jWŐM��#����H�����D~wy�A�$���FW�_�(j�`ߝ���@ݐez���Z�kx�\ڌ�8�Q��h�\��E���7���92�6:��)����������9E���P���Ĥ��\�geAtX����i�������ZnƠr���`���g_KI�3�t�3�ҁ��]dr��ޠ���y��]��H,9oL|Y���|��|�e9��"'1Dw;�;�8��G(%W���=��v��i�*c;P�h�I�\`y�ܬ��s�gl۞"���ִ��HO��~��ޜ���YU����Z1c�g�瘲�����D$��]�Z�b
�b�~��t�Q�d�B���f(��HC��xGQ���	���F���\�@?76_^��?��>N�q�Kg��m,Ҷ� �<"�R}������o����gP��F�R�ҡ�����꣭m���R�Wá���\���0ky�H��V��e Lw�ri9�)��c�3 �-�����)��W&.J/�s�g<�����Ыls��<�1\j2U�� ��ņ�7�����N�N����QwHoC?��zC4o]�:�zk�=�<zGٙ�q�zo�}��Ϸ*^~������KtGb�&����v�Edh�%N^5��U�k4��M�Z����������f���)Bm�	��O֙"}U%�b�2��k�ş���Q��h��lu�+=5�c*��@�T�'�2C}��J���B���9F�AHZ��̈́�_�=��{�P���m-g������EHL/����5�Ǻv b3 ��Ss�vg��|� ��k|ʛ��N��W��a>�J���c����p҅��VS,ϵtEx鞻2��V�_M�{����}���9h:��ל��m�%{�WЇ�
$��:��K��8�@�#>6Zn�w���z2��'�܍�5��3ф�EE�[�nI��6{J�7�_o�<��-����T��j�����jr~uy�;�૒*�$I:�O���E��}�TI`�_/{HS��p���2�������K?����I�����a�?N���;	�7�����������@G-b z%��D��G�p�Kwg��$D&��_ ���7s �@	.�C7��[w�/wQT���w �FA�Yo^WۏY�r�d�C���U���S}o<A�uD��ZB���g����!T9`I�IR Dz�|>�����[�h�*2[���ϙ���*�o��e34�YQ�)�.", �Xx6�*8���쪚"��K7= �<M�����%6�E��y(x���rկ��Ϩ��J*ו��t	|kJ�P��2��֒ɪ�QTdÜ_�ͪ�X��=�1j�2cC���QXS�����?@X�qEOI��j0�|Y�W��Ԍ�q�Q�S���:f.���Η�'v�[늬4��Us9(Hp���%uЯ�-�\��s	�S8e#>�	t�_}Gn-�gQ����M�b�|Pw��b�@�����n���T���#��d��J9PG4����e����0�G?P��j�X�'�Ĉ��x�i�}��(+{����3�xi�-g;�^�`<��q��P�?�F�V]�,�^&ל�œ����\
�FJ��MO�ߔ�u�u���z�?���ܷ?]�AYxv*��l�u�S�x���2W��E��r/[�d &������Uwj1k��@�:r��#��$�������¶䭭ETz���̓���k ���gi_��~�U1[�Y��J&$��Xi]U#6��
��͆xw2�Z�^��)r��"�N�=�Պl�����X����嬩�t�H���V2�,�޽��f38�Z�0�R{hX�7&?��;�����lFD�W��J :���b6m��4��R�a#��=ee����ѧ�.�h����I�C�} ]M&�p~���74�G\7��|5��n�� B\j�PSESp�>�A_�_� ��R���pֽ��ՐGa���W���$$��2"K��n��.�����K��'9���APa���9w�2&�d��-����Ɖ˧zoh�$R�����&V�pKbR�E��l~<F|�� ���N5���UHH{#��#`���q���XOm�:�V����Z��not�Q�Q�̀���!�ŲKq�����j�T�0�E���Wr��*!o�z��/;}� 1{���u��#:��s�L$tO�֨aN��?����=������Q	�[˛�&�����n��u�'�I�m=�)�Y�K���3#&F�댈X��Ӎ\�-��^��uC�̙�:iRz��8�%p��30��ev�~2��G�J{g���y��_�s\6I�t�s���_0?��ڤ�F!#��r��Q��Ɠ^��#��sk��(�����}u�� �-Ǡk�5�tE�pB��7Yf/'o6dvH2�����i�]M�uJ��P�)���`:-�nꭽZ��wT����URo���MT���g��f�=Z�.1�|~~���nq�b��Y��g��
���'2s�s�r�o���&��䜹�#@8h��ܺ�Y!��J���K���3���`*V7��}^�o;'�5�RY����N���Х�:o�Nѵ��e[�����R,R����w]?4k�q���O����_��\;��"q��5�߇�z�}qJ�Ѐm3��t	/c�Ύ��hG*e�g{�T��2A��7��')E�l����F��ҴkY��4����T?l
�q���^��#���6�t��Kw���s���ً)	\��J���ye������A����(H������d@벇㞿y���9|g�y�!V�z\;}s��"Z�'�_�|���_�d��S�,�	���&M����y�D]���W�/��M&N�#�fZZ���R��Ͻ����SJ0��m��}|�_���$�6�*�W��rC-�$v�r��A��Eq�>Cp�`�����K�T
Rn��~�a�3�=H7����O(Ÿ���rk�f2||<�T���� ��!z��a� �3�_�$8�s��$i�tӧ�D�hx� �u�A?�'���a�ㅃ��W����f�%ۋJӞB"��^�3��M��:��\|�U!�F	Y��)h?�l��3�3���%M.s�Ik	����0��8��U]�^`&aZ*�{�cqi&�A�n[�����qy�J-#n&܌�@e�v1�&���#�W���1����k�Яj�6��1��KS1��*`�=��gZ�B�H���ؙ@��f�;��2�e�U�y�߀#l��y|g�n//��\'IJ��v�?fu
���+�ҷ�Ƨ�wė8D�"������q��/v� �f@����� on�����A��R
�l�oR�o�0G�-�S���B��!����y�XIm|���<�i��͕4�R����U#m� ۥP��♚6o�R*���è�̆`�M���qބ�/.�����=��Y�x�\K
�>c��������E���p�n]����B�������u�ܗ�������O��Yc/�� H]��}(�F��o%cDW��珿\&-����6R��0�S�2^�鹙�f���&���E�-m t}��N��N�ė5M�؄�Q����_Wl�������N��2��T+}�ڡ.IH~�h�n�/'R�` ����oh�%��Q�L/�Vl�T�h��Q��x�ВG]�.���bLm�^��m�>Y77[�o�V��C¦�3�����'`����m�A B��՚5�(�]��'k'" �p��w��N@MY#�V��%�Ϡ�N��T N�
)�qX_АL��p�>;H�4q�+6���������4V����^3����o�2��4�&���EƸkU���)3$��ӋM�P�~�@���'����\h:lPR����t�]x=qn\!�( �+������@~w�{F��L����t=r��6TH�#D�Fٳjy��͍"L̥�����Ӱ����;n`� ���t�e�+Mޓ� �W3z����\�A~�5�mVW.�l����3w�03��O��������N�DYF��ƕ 5��'�����ڨWx�]�E�Si5��~f0�e�����&fN۸�n'Ћ�9���������z��i������`*�ST��S7厧�Ⱦ�U	t�i||���.*�\~U�65����i��DH�|Y�����׏S���,Ges�ёV΁�?#�H���Mwe]�&�r:�����A��4Q��,kܜF�#�'�y!^a�ѓ.A���l�u �qW1�JS�!��o�'q��ߚԯ�8����:��$���a�����u3c���4x�����M�_�6��Y�?�SY�x�Ϡ�����"��|��-�ʍ1?��k�{�2U�ݛ�ԉNNx����m��\�e��4���T�B��n�:H��W�6�x��W~q�
�Vn�LgF@�:�u)k9�jb�&?�����6N��yip��͙E�Y�J��bʊ¦�~��� ��/��1Z`X�"�F�6�d��,��
�|�fD��Ju��gԂY��UԿ��[4!�J�Y3J�����0⽚r�y��w=��H�quW�[�����~�П||�A�!��LYR�� �0S �D�*�4��+z5}{><kGU8ڗ���H��Qܬ�Ui&� aE[��0TG����J�MB3l�_�2��Z��(5��A� '|�*IP��YnH��h(���F�����,����u�+]3';i���BO��@=xh��>���	6�����1���g�Rt'�}t�S[��i���V0�zEF�ɟ���R,�k�r�%����dY�B��}3���."�;�4h&j./6����R����Ƕd����X���/�>�����$���',�|+�vu�U�gE,u�ƿ��?�����O�p�T�;�)������c�^��v������|68r^i����Gz�tT�l��	�'�7��>ր��D{�.�y��vhy��*����s,/i!��S�Ȓ~/P{ݝ�f��m/�Ww���6�B�z�u���g/ڡO��N�M��θji`�%���j�r� ��sv��k�)MwV��x�,��7�s�;@�5i�^�)�K�|C�# ���{O�r_K��?��0ܿ���^�¥��#��#3r|���EO�c/▹q%���p�1y3�!�_E
���������g�WvB���,�#l>1& �,�de� �Pm�"��h���+i l�3�,��B��3��&�vb��]o�=�'/�o�\4����*TX�y�K��B:ɏ��'ԯ���M&�5��(�U�{�Ŷ��G�rz�|� ���V���4^8:Q{����dչ��b!(�B~�r+������5^*O���~��ɤ�V8g	��n���	R����cy��nM��������^�ϥ/,N��6L/W��U+>�s��Uf�S��\Ƹϯ���ۚ`/?9o�<u�r�.�K��Rf%q�hm�$=��q^�L[=)%K�$���K�|?֟Zu�8�K��kL�C��[T�� H��kS��'Ҋ�K��?�0"�.�w�̾��+S��DN(}~�g���'�H�B����S5
�};�M�������/F$sҎdX�Ed�]F�iQ���sJ����,e��]U��9��;J����]��R�O�D9��{A{EU��y�p)�{��Z	
�(``�� ƽ��O���^�YX0�_N6�QC�LB:%k���\��T� #�%�G��u�4�&���i�VL'q���>2��Ksfkg��>{��[��@��f�������E�JbQ��W�>
��4H��3%���)$D��0�Tt�p�tN�o�%����%MD�a��C���=�A�(7Z�����u��:�"	R<H�Y|Ë�R!����'b4��U��̍ˏN�|�B�˖_��Mp�.C����H8%��&GG��{�3��V��EI��5�q�OV>-[�-)J�d>V��XE�F�V*n��6��+}9��,EL�Tfi�g�3�������y%��y�������0�*�pR�^��<~���ک��9�/B&u�{0mo���K[~�����Z�%�2�C���)��ű�Y��Z�˪�
).���A�F��^��;_ά���:�$L�����E��둯/��{5�E��`X�z�R�@<6��0H��z�k��]q�V�b�J'���n��nU�\��0g,�i�&����Wd�l�V�F-��(�|�뮲���l���	���ݼ;����&1�ġ���n����9�����r�X����#ې%���@�=}���n�:�vD����?H'�/�6G,����p�F�n�F�����N6 �@���_���Z/%\�D��q�y��� �÷���y��5	���F��p�=�Ҷ����U��ϯ8k B�M��G"��H�Ź���3�\;Lw{��6��VW�DR1]u!�*K�;>�[������i���gF�^��LϺ*l�y��B��:����������
J� ��=��H:��'9�Έ���;�u��T��@o�ǂ�A��D-ʝ�B��X��l��X�@��p{��=�̓8$!2D����������3P��<i���Q��8є�4�=�D�A��_|��l:�Vd�� �<v'�z:���x�
,k��6d��fH�:"���	)��z���NtdTc�q�%^��+w4y~�Ԙc$���L��W�����4������b��O��'z�%���8 �x L��]ٴW�]��J�*A��%�����I�U_���fDnŨ��f��.�pˋ�����1V�c	���g��HYY1��io�PT�Q8'
�Bb�Ҳ������M&G���ҧk�"�jmѶ@�����3x�X#��9�b� ��ρXJ��6$�^˟$�N��47uΥ�Ϲ��gP]��ʡ����P�Ŝ�a�߁ ��_���1�Jz;�2���Q�S��ŷ���ߌ�.��r�:����]��d��ż��f�$�sݝ3-]t��ɷ4C:��H�w��1������a�z'�,[�F������_f%%��V���w��!G�^�җ�o{�j��[��_�g��;/n�4���4�j^/+��gN�{FL*��b���W� �_��6�c��1�S���m*^��C�$��6t5�rL��-)��{M��5�{���/`�k�]m=:L�����_��hСlBGLP���w+��C��&w�	@X��$��<r�~E��ޘ��U�����@J�dL@�
� ��VH�q��W�7�nF���5���W~�O�$�#��II������Dˤ��E���AZ8Ǩ�]����V�Sn�&7���X!Bj�VD��f@��+9(i�%f�I�$��M������,��u D"��ñ��ν=PlD�h�u%';H�6�P�wi)�����n�N�~�G��z��wY�d���k��3X�Cw���{��	��@��5�"/w�쯟l{d&�V��
{����~u0'�e�e: SD�QXLۗxkB�X����Q��;��sM���j�G�D��W�'��b��&>��u>��d�bP4���� P&���6���4��IUc��Q�����JV��ý�$)
�n�����n)�sc
NeŦE\fH�g�y�9�G���>e���&�)�],^}E��Y<�V#=�n�_�0�����۫����Ȧ 3��̴���+a�@�#N:�~�%CVIćfBhD�'
�Ô�|�n�΃���.��8����7�ߘ=%�y�qY�ݡ+��C7Y`8��ay$-ר���p\���E�\��ξ�#d��q�������`.(p+�<2��˽�V�!x���k��L��û'�@9^��`����ӽ{;N����:C�y��>,�A*����
�1e��RFPqJ�8O�5��`��$��._����-�S/q����Q<���;B�մk��31��]��� ~uLw;☮����u		U����s�0<��BX�f%�<�G������%&����>W�%T�,B�K�#���3��	�3I3�%�iO�"�`AN�b��1E�(y���=�g��ġ�9���nsTY��H?��Y��ʿpc��YWuDH��]4���i�-A�atQR��#e�-R)ɘ���.V�NՊ�飯�w�x��h����OP��Ec��{���Ԁ���-X����\�,�ݖ�# �ݞ�:�j�a�#!�>J�3�ʃ]�G֒
��a������n�ʾn�E��*���m���\�B����:ݞ7Jr�
�)}�m���<J+�b$��c[�JB����t�^ȌN�.���3���lSZ ���ҵ�~-�C�깯]�ժ��p��������p]����"tJ7N k�,�\,���7�͸����g��C��o[)nѕ�yѰ4/�Y�Io�ai5�dS��6:%i���4ʼc*��m��2;.�4� 㵛�(������k|��{�]/m.Ȁ<��mFB8C����U�	ġ|�:O�]�����̮�����x�����b{�z+���ʲj}#l.�Jl������HM�%�5�0z�ɨ����=Չ��6/���U|X*=&>P��ճ�31?X)����巼.�6pp[*M)�(-z?{&�<_,?� *���q�@?C�#�'C]��T���O1-r�ôD��o'3Z�{h��EIڵjm���%�#�������K�|��GD���!�Z���ZY�%��g\
����&c�{��}/�O�K��}��8�����')mHfns~��&�1Vޟ��:��%�����?�9e5Bz�W6»����k��зd�mk7ca!������D/��^��=,�&�
��t�����̷���y�Y�NrP�b��L��C��(���]��N9��l>��sѕ1�-,�&�Czˏ;�~U���2�?�okۢ�&���Ncܮʛ����x���
mkq���Q)��gp���-s�	����������W��cU*!�h�/�S�;���DsNc ���� �w����̘^[WVtR����w�5�2���jwJ؏+�����C[���ؿ*{�hd��/���+��J�@V����&��Mc�j^�F؂��ß��{�Ȯ(��ͽ�Ц�X{�γ4>�e��on���1^�Z{XPi�/�|�?qϩ��T����+���(�N(����'�
V�{S�d�v�_$ͻ����oq����6��fc�L;��8��T����/,�<[=>4���j�qR�����Y�ƨ�-%����d���m0&�糺]�LE���vv�l�-�ki��*c�4�s�`�1,�ԫ����� �>�ם�"7�D�W�G��]{��*��?#��}с�U�~��2-N7�Q�=/f}�<��$9�p���9//Ĩ�|�PS]X���F�G����k�9��!����@f��ֲ��!i�����������;Cz9�"�񽐲�>�ԥ���v	�,�u��2T�c|�r����U9r1�o��_J;�p���OJ��=�1��q�g�A���R0K[�칎5����1���s�-s�3Q�r�aa���~[U�dg�<|2w>U��m���8��/΋�ñm��.s.S����g��/���sé��SY���TWt�i�3gX�OV��ة����՘�6�h�|�ϭ'6�qR�)�z�#����,���+I�s�z��M�D�;�S�~�^�����|T�f�(쳷��j�x�������i�(r�YIe=���	v^�������#n$�F�sk�ƅ~{׎�7������d��[�ڄ4=��p�`ku�*e��lԋ�jmh��큮��d��:]0��MF�zi��ib�l�5���D)�Hmwm�f�Gn��B�c�{��ws���2�:\,�4����>Bǔ��W�,�B&Lw,E>��>0��9�����z��nHj�g�z?�^�$�¬S�{P�m�ELҬQ�����_������k_�S�W�<����.�3�r�����u�-+O�؞�����L��L������Com���&co���)�`�gq>R:Ye#��o��u��t �VV,� ,�I9���E��$Nn]�Z� �^A��a�l���f���$&\��D�h�"L�\ocTOTr���u���`ɕ2���<����a[QNp����
H����JxZʱ'�|�e�~�m���կ*N�A�6r�p�Z0KW�м�MUg�H1ɥ�n�~�3�c}��!=�rEq�d�d�Kki��3||�IzoPM�}H1c*sVp�i�4i�x�F?����5Ϸ2^��H���"<b��O�MH<���0��Ǽ>�z��Ы��D����3�a�q��B� U��*�iȜ�d�wb���)�Ǝ$��j#�v\_��)�n;Zg���b���}j�'����p?�� �5/ν�T���V4������݈�v_���2�����l�
��E���G��E�|�)�d���
~tr~�<���f8�p���S�j[�Q�����7�
0�B?<�Jxv�;��;��V���u���P��?�tlvƌ�[L蕖&��́�N��63[e1ۛ�� ډUʈZ�qvK�-\q�i8u�v3v+��uՄ��q��~�j��Z�)�����ZM��I���&8N��|�� �v�x=[�){�W]�#N7E�^�^oc�ԏ���w�yv��w����q�D�	D�\�#����?��{�]��k�:�-�}z�P��5�-0��@�eT#�Է��E.�C~kDy{�&�ׇt��K"3�*˨��钦�?�.�x�vD�ˤ&ʅ���f��<���/~�,E�偪k���3A�@z�5�|z�E���:@�i��t[��)1����O#\��~g.K�g0�]\0��)� ��O)��}�����
 (MD���z���7˘4��c�ffC�����#��j���P��Wm�͗�<�-q�iؿ-� Z�xB�еq��L��ڗ�\��N�c�jĩ7�\���y��Kt��E�H��'�}s��'�l��6"_�D���3�?b��i}|#8� �n;�Fr�sR���x#��Ɨ�f�#�I��F-	�e��d������UiUU������+��=YR�}����6�;o����#���e�[(�w���oݶ��
Q�j'�ouK���b�Ә~/幎��_�g�s1��b���J�p)����+*B�ġ͇��'�?�A�@ �N�(�0������a]���R��}�x����1��k���$c��Q?���i�"C�e�ʇ����.����?v�#L<[�P���,b�
 ��P�O%�[]�2N��~>��>��>�ܡv>ힲ �t�
/�H�9+��5%N�^2�3�vu��Ҹd�*�4YH��K����Z���w�ȓm{���{��Y�aa��5ٜ���7�0��R����q�2�i3�h��}�Wi>zB����ӭTV��0�$O;�ܪ�y���*Y����x���>�Tf{�a���D%-*'�[KL��Cs��ܨ~����������v�ND��͚=ɮ�o�𬁢
�*�_c�ׅ_���<PI Ç��;�9Vhjz�76�6'e�p����U�j=U�8�@��X����=>�*Z(�y0x���[�>ܹ�p4�*��`[1Ϻ��oU򄀏�wF��W_L{�"��B(5qUh�&�3�{@��5=ʕt�.��Ӄ.~���~H�
x~a���oy�7-�v�*T�G��T�^�q�-����N�>��ʩ(c����[�E�>��(��"�]�Hwwww�H��H�tw�t.�KJ�s�����?��7��9��3s-�Ar�!�5n#.�d�ɓ�6=�����kJ�2XxNH�{��c�D��dP��*x��@�ڙ���4��8����@m�PCӡ)?sQ�ʐƓgqA������������̴�Y��I	bh��+�2���y��^�9�#ܵI�_�`��@������EI�����w�}�c�'��g.N�7c؄��w���*:H���Wu�<��t�+�߀:��/uB�ٷR�����W'��Ӈ8X�?W���j�^yF�X;�����	ˍ���c�:k���Uo�v��YH/�|X �cC�~���� �74zœ?���ķ�+P��k{��l.+}�}�:3�[����!������L	�����'@Iɭ?�wW��U$}�l�=1}��	j0c��xhp�AM���Iқ�Zzs{���
Du|�="#Y�L� �Z/�����)t����g���{p��e31��D(c[�+\t� T5VLD���5z֥y;�r�k
̃J��
��~��cT�n���s�&Q��F!��"���C�j�@B�L��9_,�h�T|ꌻ���a�N��f�j���W��jiB^�������P4�8�8w>��L�m�W������8�f��Vԁ�t�G~�ກl�����G��7Ѓd�X�G?SK���	��ҶtO28t���Ԋ�Ȏ���½��������FUh�:�=�����ıi���Lh��-lI�+TJ�(���#�C?��bY�z���MnU��)��a�d�}Ldn��z�d�����g�+;�C���9��kJ����\@�y^��c�oX�#��%����Jet��u�M��rk~�d�jXG�*W�Z���Y�����"!s 5�G�!��
`_��"��q����?>�I�H����{�����)(��=�OY�+��Dy�;N�������`�,��2��rS՚U����)6{<�M`��ߩ����v�o���zkG��'u�H�������Vf@�E*�Ǭ�F���B��s�d���ij�[�ּ�Z�c�M���c%�Q�]���ۤ���sܟ�������)Ъ�� t�X	�9�f�i�z��φ�|���{|�w��籱��K_i����zg�֩˃���ƚ�r_c�K�[�f��r6�
�ausm�d�Z�^���=-^��D����V]n�����"Ni����6-��dB�Uf�����O�,C%�Z�a%�� ��� �����*��څ�|�61k����eE�5v�e���q9���Q���/�xG���ݗ����q.�J����UPO���ԯ�?����&d�<�	�Lc~\�3��T����hr{�0^�'��A��~��B�-/��K��2(K
~�ɋ�d� ��Z�CX�wcƖW0�3tT+�!X�L9j�!��>N}5VD�R���Z]	~�?��$�#f��U��n��
�l�j��4T,���F��4� llWs�U���j�O��ID�7Zpfr⻚z��4@eS}({@{%�^�ymt�(`}4���:���H͌������\��n(�8w��@4���	�=W4f���'�TaȦoC{j�<ҧ�W^w/���BB1��аq���Yj���sFB�Ԇ����F+1R�8���������`� r*�ŝS�1R�?a�Cajн*I����4�j+������Cp��D*M�c	�vTl��{v�����񩎟��w�[���Ų�'�pz
����l�!���������m9��Y��q;;\���e^U���E�22�V���~��Û��'r�a#9/�)�;3�Y-$� ��d��Y]74��ΪTTg�-̶�<-/�<0�78@�R*A#_��e�\t�[1tF��}�+�C���&p*���8����JKN���(��plͷ6����}��ڕ9�i���;N�� �5��VS| z+��Va/��+'��[M���[<��I=���ߥx�x=�l}�X�C��;Y��5V@-�JD��<0A���"��Z�=���.��g/|�"��3��r�7�ѷk�� z�H�XUnpU~�'���+��ɔ+k�n��C�I�Ö����.�q'������kw�����U� kk�q}���tҀٜ�/ᡝD�R���d
�
�!�C�%�4��SdF&�o���.C�ߍ���rO�u�0t���3e���JQ�q���f@�*�t���
��������P��}�v����E������R���Z@x��zm���ek:���fʏ.�����d/�f��{�Y�ur�h�7	�!�|�V�&�� �tB���i�rq2͊E�*2��0VEZ,˓��9x���\C�dЏ)���<��w]V�(�yNo�gp�n�s�k��n�n�}��#�e�-����W��8�@\�3R
1��h�oe��g�kA�)�p��H�t��Qs㆑==_p��Q������)ee�p{�^0ۆn��I�a��U��$N��O8��	wa�-È���_��V�[�)����Xܑ|j��N� ��}q��L��t�@�����4Z��8��Bm/�њ�<���,`�V��#��������M��5_hXfO�.���[a���M
��
��W�@6J���Y_� ��n8P&]��y7��"���%�m�������U��]�0Z	BJ[`'��G�:�	9e���I�a��ڌ�8���c�I�3;����״�m��*t��~�>�|E��W����r_��q&q5N{H��ю9~����4�G��?S7��?��BvIQA��σ��ݽ=P>��@n�'֯�����͟
�5����Q�W��ƫsN"s rJ��;dG\�ї�*A<���	ruQ�r�WJ���.E�	�=����4G���)�#ψ�=�t@��Ҝ}�`���r{*�*ù����{�ѵj���h@s�����ٷ��q*�݃�4d�״�����W*��
\q2���ί �����k*Ö0���
���W	Ԭ�h.n��T��Cb��}�(���5'E3��$��?����M�0[������uzAKh�?*�3*��݃t���4���k#��q�qA��vf�;"�o�/�"�Q�	hx���V�$RJ��T	���F�u�ӌ%��| ��J�!�Q
W����t��Jv��ȍt�������2�3g��������G�c�l���ex�����W���p����f,�kݥ#����PO�&�!)7�Q8U�2r��C%�շ����R0�.q���j���G�����Ucr������N�谢66$' �қ]�,O�z�w��u��·y�>����s|u�^�H��a#DQ�sU�e�To]rUO�YТ�����H����tt�����Q'�!{�6A'����A*3ĉƬ�i�C=39��������)4�G��ǻ+[�	�u@ n�2N���8(�p�](���˯yt�e�M3S��Պ�/w6;� ���6%\}�w_�4�mٺ�W�P�fV��'��y ~y0Ewa���=R�q�gW7z������ae��c"ѫw���h�?ƥ�Ϧ��.U� IT#NYh�ɣ--`�������W�:	��(~�E���� �W|"[Z|=X�&]7� �x ue�?��p�H9��e 5p�@ha�)�����\9ΐ��HJ�,힉�B�MsAxyN�϶qw�:��|��p����\pk�
���Fe�ۤo(�	�S �Ɲ�Na1Ki����o�Y�|29�/�kG�W8��|��wq�V���~�����;�K"έ��M[n�:�*�~�aoX��Z����{U$)���1��<E����\�2{qO��Ǚ�&���E�����M����I裯��0 6TH�u�T���00Y>&-���.�P�5��q���R�_�!�i��8��X�$�I�	x:��mDң'0:":��_{�]�`�\�En����Z8j�ۧ&����3���ۀIbc�Վ(O 4$^qi� \B_�E9тk�%�|��S#2����)˳i��d����%<�v�RҖ��it=�NX�D6��<�@t�/NU���at9.$�;�.�pk:�I}c�byV��;K-���k�d:�������~F���cK���@�GȖ�u�����hAJ륿��l���b�}4B�(p2�\��I$O��>�>�b�7
�w7}�o��������1)�D Va4,�@X���Ds��^e(~���l�Z�WMD��� f�]>5��l�hx� 2�`N֩N���?4�خ��I>�Ur�����~�@W�/D�M�t�_���<̶c�ڶ�� i7�U�a�~R�;�u�+O���I���/Z{E��] ��
���1jaL��S�M�&I���g����s�w��C�{����y%x�AΪ<����s��2vp~��4���`��U�;��t���㑷��R	�W��>��g���Q��P��׆t�1���<�ኍ���$#��_�zFx\���T�nZ�3��5̛~d�ʐF�Q!��x�]f���o�����#a!n�2J\G�yy�]�~�&��'�m�%�7��� �P�E�����[𸨈���`xn�����T�_4��q�׍<Mʖ:�7,�ˮ���b���pұ7~�ģ�={��S ����w�l۾��懖���7~��QQ��u�u��@��*e�IK*���Y=�x��꧖��kD[:[�C�K�Z]TX�����@G ��)��X��<Z�&&�x�݀��؏3�3/��r��������E�(7@g|��6�(lrZ�W�@��F W�:R)�!���S�hL^R�/�ѳ2\�=�K1
�Af��dL���DĈL���_�ﮩf�	 �1wS;�N�2��_mQkO;	cwFg:��kܙ�پ��5qZ^o>	�o_��9�K����udT�#	KP���K�ihy	�Zi���Z��������;qF#䨖�~��d��@DA����hd��u��������A�P{�SV"�yl�>��V�1@���k?@���e�q�+C�:Z�Q�S�E ǻ� �vxs� ���x
�	-��l�GʤM}!���F�q��'6���4�����~��)�qql��Vx�OTx\�A��_�J��pS���=3��;N�Z���dZ��Ądh�Z�� ����!��N���J�D�/����<���ܸL�=��#��~i'۰���h)�j�o���p�N<��"���>3�If-���k��g`�O�aq�w�HG�-I�>31KDB��n��@�XE	��o�%�����}-�Wʭ�S�Gvo��`.5�v�o5��|�}jt����N�3�!�ip�nD*� �$n���hn��I���߂��,T��_c����B��Y��� z�b�0>�o䌵v��M�ew8n����Jc+]�����>gG���Qڗ-��p9�Z�&�Ą6�T{�����dC+i���+�]���39ύc�Yy���1�Z�J���^�����ܐ�~|.������wAZ�ҳ�ͫ[��h�/���[4���d�s� �/�/�l~l0���
���T�k+�"�DI�!�����ھ�^�`U��0K]d������e`I�̼�8W�Avi`xOd������^ű�D~c��`��\HV���o�vu8�n���j��X)�y.�JI?x�S� lo��'��,ז&P/��A|m4��u�	�\���T�K��.�:36�B�в��K�v��꺪pW'���Ru��5M�Ζ��c���TtEeVn�O����%�!̛��Ld�	x+9c��R@8D䜨ن�7���/�e�\-8u��<���#ι��q�$x�;|��ydޙ��'�"�2I���6ԫ�Y����EF��5�:X|�ݣd��V%������]�E��a:�R�V�����RUO&Ĥ{�I�Y}�j�K���:��&x��������)ĵ��@ح����ؗ��}Ȅ��U�++����/'���a'�4�d�\��w?ј���~<6Dܱ7�.+��'�]<qAB��3��+5Ԝ�W��< /_�<`���\�Ӈ�!#����򃓍��H�|�}�k�/WeH=�"n�7�6�;W���WL�5	���E�"�N���1�O��h'Q����S� ���AU��BT��+x�ċ�p�o_�3X
O����[
���4�ߐ� �pݸN�N"睎7I�#Fo�y��BA!����O�`�����)������P@�b�s6 f�KqB=ɕ�:D��ē�v��Z��+�ү���F�z�&ݿ�'�y�̃�ٚ���	+´P�D�lv� =ǯ���OR}+3m�V�2V"�_�q�o-f����*���l�dv�X����3��������Y�RWtCP_!��7@���dnٶ��L���5V
r�Z�F}K�7�.*��.���O�Hባ>@I�����	o�E�K#)q�5��ك��n�ůꚨ�$
0�]?���䚖x#�c����6� �<�m�#�/�C�_�Ju�MhE;�;=2{�/�]PR�"< i\�j�wɲ���>�(\�����g	��<��k�p������h*?n0l�\C�6g���w@et��h\^MXD8�م�d�v�k��ۼӹ�֥zgn���+;t��"��q����V�6d\�4�`gtɸs�=����&� ��l��Ҽ��ZpTa�Z��n�A ���ť���W{|�?	�$_W�P�xº�d��p��xo2���cSS_.X��^��g�E�J0\��C�C�_7�osv��s�p�uWrn,O�H	�w�8�T��s����T2�u�*��[z,��v5���}4㞖S�>b;i��^��Z�w_�9��f�����M�{��>9����(8/Ǽ��^G�/I�(�����'єU�7��ʖ4��>��5�?� v-4#���{�Ŭ��]�"�{ :>޸�r��Q4��/�F����̎c�.Zky���XA��[mG�6S�x5�q.C�Kz��W\�t�����[�"�lXף�i��&�_��-'+hM Td~�,e�q�$��{$<��𛺨�>���}`\3x�k���E��}4	��b��叀���^ovd���OL��tӈ��?�$�.B��mP7 �ۭ���ix�VϾ��%�z������^;n�DM�05�}�Hh���	��kG�+O��-���V�!ϖљ��6d��GJi7��u0���"�Ս\)��y���{?Y�e�˷q���4��
NGjv{��t9�p�+�ScFj$Q��Km����{ �I`f��)&F��mӼ��	��|J<���M�mSڕR�@���W�x�n?Զ_�*FJ�xd�~�d1#`�M���+A\�1��Ź�;�5���r�%�S*�'� ��be��%�]��n熆�� ��B"��ᓲ6b���
w<� �i����[$��ߥ���＊KP��I�0Kq��&��?[<�k��}F�}
_�F$�\@Єg廌��vw(T7�	Q�-�ﾭ|�#+w�k	>���e�_�y]jTJ.��[����_�E���CX�?����pC�iJW��.�Pw��i0H���trRT¿;<�-��Ys�vq_կ�K{q@W������L�C�PE����7淋? ���@^�A])A�|ti()(F��9����,[=ܕJ��|���h�r�0���|)
?�v�s���� �@W���}��z�_j�D+�,QĪ����S��%�!��ׄ_ׇ��u��9�m���T\=D��A��P�
tQxG�ԝ����P5�*P�(�1<��o 6)�-$()��j�4�?UVRQ+6�;�#����b��bkdp(��y5#�	�k�u�pn]g
��ŵ��X��U��{{퀿�`J�ʼ���kH� E�߳&���ސ���ȔwXkCCO���bj�x�]H+�~���_v3T����=��95v%��1��U��0 ��O�Ap�t�D~��k����u��=�: ����qf�f�B��:�f�7��F�༏�	$�Щ
Yu�b??a����2�A�f �鋁����J��ͫ"�2��˽�|ߡ��������kÎ ��3�&����ս�����x�u<�v�x�\��[��N�(��]&b��ӵ��m�[�k[�9���2싛���d�թ h�_�BD���G@�)<�>�=�*_��N)%�/�h�4÷f������"�]ģ.��%�?q�p�Eg�%�|�Ħ�8����@�=��6I�;�E?� ���+�����4�T@-�f��2�`���u�o�(���ֲ���<x����{Nֶ�1^�UESj�p���̬�}�� (l��������I:o*F�yj ��NB�A���#�B��Ʉ��%���h�6�G� �$��dq�w S�Ņ<��(h��@�͢}���B=8�����aVv�/�]���E���.^���g�gq�K��ۀ3����=����4%�g���lG{��� h���m�pd׸\FK��9�(C�f�Y.��"�`u��Ʊ Iȴک��ȑ�實�<:ꊅSE���lH.�w@쪍��6�@��T��-M��$���2W�e�G4��SX��<B���6{DWޯ����a^�-]l�Sh�*n��S�
~{�_� �U1�x�������� �(������>�h�qC�����ɺ9���+��U��Bx�~|G�q�p9�O,~>oYe1c��gYcf�x���Prbrr	�ч��Z'�#�@r::�N��%8����	c.q{m�O��VrJ���
�D��$g-�Ӎ����A@���L�������DV�0����?�7�pߗN��p~X���3P
~���M���B[T7������N �F���>g]��u/�& �A�̟`+K^��@�e|�����f�ij�{3���jb42���`CK$�Ü�����M�7wx����Ņ	�ײm��]�x_hIa��c����A�r��X]яߪ� ��+�������L����a�ڇ����B�q_ee��D��/8�����G��%�η��<op2D_�������Vd}��mf�:�X$*Q�������[i\k]E�-��\����Є��_ND�Y�xm ��R���+b��9���\h�U�+��p���}��Ӕ	��6� B>��Jz	��K~�t�'X��L����,��b���_4#�:��&�+n�VyZ���NW���آ�ԋ��=�TV��[$�GO�3��?H��ᮊ�����]�~����|��wuJ�l��ٳ4��� �PD�$Ȁ��]Q�N�:��.�F��mp�6�ƪ��H��*��nq2ј����Â[��bJ��Wn[(�0y��#m��	�_ߨ����C���]M��m2��.�4U� �Jgܟ����k�7Þ���A�m��m�ݑ���g��.(`y���؎6H	�D������b��|xa)Tak$��)���rXއY�������:(�@W�ڸ���h����5���m"C������9�[�_����G=���.͠dZ��Ij%������a����K�A�}�f������@��C���Y-��'z"p�+��T��sՖ��B�w�c�!o����zoE���!?��}�V��v,����&:�dṍT��W�0����}�_�87���#k���s�4�عa�M���]7E]�஍bb�UC8 �3w�� �8&��ą>A��.m&Mz�O��=&��=w�����*T	H�ޭ&F-g�Ç�cT��:y�
�/��J�Ĵ'����j��4�M��݋���hJ�رL�ɠ�Ez�?�mr� �&��RѵY-L����`��r���ʛ��ӻև\�c#�DI��o/�*� Q%<N�(�^c�������D��uY	y�A�S�����u�mȫ��ݹv� ;���8��^�9u�'��?�03�,�����У��8H���3u�kjsڭ�@�Y�vM� �t�vt���9u~�	�
��"��Q����Qj�ɾF��y	�$�_h��6����x���^��'�e�̡k�y���xh_9s�k���޳Oc���W��K҉ ���Q9�� ����	ڝh���Y^�[�s!���+�(��wg�cϿ�T���͆^���h2�v��1
&�mw8��[:�J�O[����"@8��k��>+[��2n�,�/�Ճq��#�&S@�h�<+)+;HA5N�_ru��+�9�&Aü��-Q@���t����H{����� ]T�o�w~�&9�n9���tU����.��m���FQ
�m˼*莯�J;i�Ze(Y @�����+cW]<ksNΌ�g^P���j2UPi�.^�"L���k�*��vps�~CC�[W��_�y�7�2��AJ1fr�/���a�~�3(�Tpm��̬��t����A��S6��|e�=S&Q��XG�.� ��՗+���>���̣�m\�p�ձGҸ`�'���7�9�g����X @ 4jo��_�g33��nD_iWKf �d����ϔՊLxul���ֳ�'�|�G+���̔Έ~\�����N�3�X1�@C��\8�3<\�8�1�/{�I�5tK��{|s�x���ţ�z`I�2O,Ȃ��� W�ɘ�kn�B�U��Դ�����r!�W��>Z��q����G�O�������$*?V���M�ղ2X0]K�s�OL"h"�`"R��g�	>��N14s&{jS)o�dŸ_!b��n%Z���J^u=��msx�}�0��⾒�]�k A2<����k�o�5�CҸ3��%>�ۉ���hP�=L�Q=)\�M`���s> n����5�����"��.�,�����(	� )$	M#��tȆ�e��ӡ�`���<�_�:�N�+*��Y�){@s�`�^>����=�'!
�<��*��Z��竸/��������hў�^_x]�6rJ),jj��y���i�����ک�}��N�N���w@ů�X��A|�-ߥ� >Y;O����e��\{0%٣]�E+3�>���n�xP���Av����Z{Dr��F�Ʌ��)Ǜ,���L��gT���2~_�r��݋��j�<����<5�Snf�Ӥi(�Ŭ�5f]\kp-��͇��'o''�;=�I 9�D4A������e�������A(Ɇ�'.m����_��ݤ��ܩ�5)Ǣ�)i�,�F��Wk��#)A�m����u����XM�K�l�!�[X[[�x��ƕ���q�iÙkYܟ��[U�)�A���H� �N^6);2!@.�:��2W��2����]��=FP���n�pk�W�Bgw�!k�A��I6NO��B��t�%T�������q�ۼ�z9����p:�K2<i���W��}����r9d|3��?P�������}����B�'�!����L���tW2ˉ�YIe�	|�1��{4��ք������`�t�/P�~j'�YCl�6_͙��>�512}z��`2����\�9/��:�����e�p5��n�;���L��ji��-d���!x��o:�OV��̡M
ɴ�����B� U-�?+l����M��L��u��z�g��=�z6p }x��p�)�������R.�𱱶�9�U����A�U���I_I_�AԺ$Z�r�h��|ŦǾ5�\ݒa_nH��n�q���Ж��/�����k�oa.�'��]��,dz�oddyV����/Q"� 3���~��h����� ��p��y�E�b>�L�ӡ6ͻ\��Q10~�S��n4x���"s-� ��-+dgT-��}�|�a�����h ̗�~>��b!�V��eÕ�3��A�/��)O�G7>�y���g�!�g]ܝ��|��P&���;�R�T�v�,��Z���m��C˳ʋQ��	��&\������ֶ�n.��[%B[�&�/dW�?���P �G�/ЎQC	+M�Z�����<�eKkHq+`�;|��U���T�[�|�0�cò?*���lS�}�Y/���l��y���2 o���z3�rk0��-��V;��I���R�L��7y����ב5��/Jx����pV��9��@��Zھ ���۱R����>�ߪ"��sg�P��i��t&R��~�tɧl�R5��w߆.#������	���s�;)F��D
lN�殼5ҕJ ȧ~�P����{�������5m��r��i|#(���:��	� ,I��l�_�H����o��N�U�(� 0���jz�mk1��"wكi�gF����$���&\'��ۦ��()Y�_ںI�_&��YK�=��CJ!n��l��H���K��xG�������t�&D�!�y���w#�HN{!�|�ʊ�8�����Nky��شj��V�*��=p���^���W��V����~��*Ez~y��%Yk"�/�q�:  6�$��(o�����hw��G����xe�)���o�mG�|6q p�	M�w�?�tw�=��W]���c�*�2�F3J�g�D�2�w�Ob���}���G�ܞ��Z}Z� ����~��~��y���-�U֦q4�϶�ش��-L���@G	�xQ�K��%MgC5�Yk�+����� XhFk�^O7Ϳmy���$�F�2�Y��iЋ��zni��lu���@a�iD�W�����ډ �[��	��o���2�H��ѓq��'�Z�$�"�	٪׹s��Ӟ�T�06"��p�.�DA�I�-����挏���Ť���K�BT���K��!��<�O�4W�+����I�6l/�?���qc���C��	2��(b=y f*�q��@���͖iZ��4���q���S�]�cg�H�K)<es����F؁\�^'�Y.`�EG�)��Ĺ	�w��笿At����V2�}�}��li#��kITT���ӥY}*TS␢��*�D2�x��@d��t2K�����z��aQ��s��{r-��_D,�l��	�y�$C/V&K[�}ݡp�����XW�a����g-�җX��L�]�����?	�Z��ҠJB^d؞ˋ��M"�f���EWc��fae��2����S2���Μ���A��_��'곡��z��C@g�#+<�rf����Q �
Ly��1˝�D��P�ڸ��k�6a��e3�S�C)�Y������?E�W���]{�8u%�~a݋7��,:�\����0VQl;�c��ڗ�B)�=�n|@#N�kƢ�=?6�0y�v�c+�]nUfo ��)�z�,��bhl͟%<J�
�\ i��]un�Pb �"p���B���MZI̱w�@���4�u�Vku�.
)��+���s)&fod�r����(�n�z�lvЊ�����zf�0^����ԏ�O�a�}�V�TE��f�t%�ǈ�Ih�%ھîR~�� ,��4���)u����^[��A��ssW�����~ɜ>����!'��ßta*�]G�V�F6��)V?#d⥈ȡF�T���u����������?�3_|�J��S������'u+]�9����y��ɿ|׭�ݖ��:�?��!���X�D�%nߧ�铇·:_��vVP���H 1g]*
�$pV�g=��1ڟ[�Ę�R�sB.B�w]p$}��G��v?�K��NҴ���L��{�	���wi����ۿ��sD�D�7��?z���0���D�pcK�iЩ���ʻ`�؉�~�׎ʁ��م������a+�[?W�V�Iw��Gp���N��0��쪟�Tz�Y�X��������'��8�z
:S��L�	����ьI�S&$]��&�CK�W��$�Yy��������p]r㥴��
�``�Ud��zt�yo����Ɔ���R���vi7�!R�t�Q�	�ҬiQ4;)����-}i�i��e�gc�I����	^��h��8i��U&�jȕ�|}�5ZQ����K(��\C�t�i��پ��}F����F�+�qL��H�F1��_���,�L�]��c�E/�����,��8�(��4d%��C
k�\���`���f��49b�.M&�O�倩d-ا��D�w�yC�&}Z׍u��Y���c��̃�q����6Z%���#l]�u�ꜫ���s���$�9_����k��S帑&ޱ�2�� �N�ҧ�4��G�o~��|�L���["=�j�y�Q݂W..��u�T�P��#�k�B��Gw�Y���'8]y�~����0�W/�h���+P�mN�q��ע{�KW�t`������?���f{��ls�-��
&״�7����f�0��ܢ��IS((Z���s�iQYH1:���Q��1��|�3PG��Q��Z��/�O�)�YF��i�A2p�D�'{����t�����Y��v���*���J�u�zj�&HXb/��!��{��iGd���m�%�'Ō�B�i��h�5��0�0��ҭP�\+^��lVh�\��9�0�d$��ߨ��.�$��w���b�C���/F��t��2|B�%Ĵ�#�/�����mwwd��P�@X�0�S�l�ĝ	�4��%�d��۪:�i��ڔ���k�nSFB���2�sr"#��Ø��H�s���{��F��[���e���~ʿC���[z�˒��Pb�q��c��x�����S�ï�:�^W���'
�q�J��ҩx�g��'��f_�,$*�a�ZQ�����n��L�"N���>�uE䞴?x�Ǣ�&��ڈ8>�2\}�s.{Ü� ߀�`�w���ݰ�����9����T�Q��v[4���*ؤW�2� �`��}'~	����>5�ꭿԅ|���s�E��s׽��d���N�c�#G ������m��q�-ЫX��AG\���/_�!6��2C�?��sS|���ygJA�y�m��+�G\zګ��S�<���\Et�?��ފ'1�M�����XOI�g�d]X����˒��it�Ao�~G�'�·���jg��[����-No.n�<�C�&�]�~$�g��=���$yo�4�L$_p�ϝ׫��^L*�Ol~F���7�����s]�^�,��z�v@�:�>�۲�>��R�f4d�L���An6���w�Bk�K3Vߙ�2����y��G�ĭ� s���Y�Æ�c�Ŧ��0����;6̚����G�|<3J@$r�n�
mT�ދ�}�z	|z�?���(�=��a ����2T��C�l~�Ȉ>2������.S.]�2���\�����>��n���D��a�����L�����%�R��w6t@�����M���G}g��WO�~���P�>�b/@�֬pW�P�%nT��w,��m��ſ-��~���L�q!:�j�u ��tv�����?���߮�I]�q��񦃞.Я㒾���r}㽑��dЮ~�Lx`3m������7Y|,L��6j4��x^'([��F�\�a?(�<�oTwf��*���	��F��o6��ɮ�]�n�e���z�B��/��t��������־���ˀȯe[��l@�v>��,R�������D��bgl]??�Z����tm�Fp�\=?�>?�z��󪞸byEH�&�#�c��0eΝ�8����� #t#á�;W��Ŗۊ�#i ����3//���)ym�7�L1G�f��Fy�o�7�b�sx��	1d�]�3����Z	���c�$ٝ��X�a¿`*�I��q�T5d�:54~r1�p��]ɢWb����V�N��"$�t�p}�=ީZZ�Bh�'t} .��D��ж$b=�)y/0�L�i�[�*�u��ֈ�"Tӽ��b��ZN�1���XNb�aa>)@\XC�3���6�lPY'|[o���B��6��ȁ���wR��}(�/7o�[yDݾ��
�:�/"�'�3�-|^��`�"H�b(0�|��95�
�#�¢�ަ�L�[₧oHO+ޭs=�ENAh����.������j]�"#ꐙ��sv�lG)ԘU��"�鏜��&���A�o��<Z���^���x���+�(�2��O��z��Jȁ"��M�2�gO���
����� �L�tF����h�0�)$������l���0*����.�?�*�ѓޯ�������v��&f����w��f�S�>�0�Z�-�GT�Q#쇟x�{�9%G;p::iV�  Ym�^<�W��jǒ ��o0������.d�h���Q(F����ڐ���a�̵�x�d��R��G� �K�RS2�oj�=()�h߷|�#z~/����T(�NSuW����XFm~a.]a?�w��L�{��˖� ��F���/�9�f4��GoIA�oګ��w���X YtZ���u~B]��:��"J3lp�b�vƯr�G0�Zu�5�����T\n��2x���Ωh/�^��Ic{�'p I@U�F��t����]m���$�iŶ��
0&���k4��P����e��al�$x��w��m��L�4ô�kd�ޣ�����Nf�Zmk̸({.\�YZ�<��p~SN�\^��gc�ɹxF����Ǆq��3X���%zU��j{��g6�/�_�;`O��m���BKj�Wp����빤���A��d{����>�'���VE��9S>{�r������@�� ����5��ӵf#ٻ<�"��cQ��;ceD>#L	���3�L�� ��?�Xp�>��"4�� �%R�5�0(`�ak�G�q���i5�+9[S,U6b{��B�,OC�ǅ%�h�l�^zK�χ��r�Eg���>L}��~Z���(��1��B2�E��V6� �o�@�����.��@�V,ph��3�N�\w	������m�Y���x���vh�놥6�-#��Z�TA���"?��:�h�����>e%V�t���Ȥ ̽�$���ʄ�G؀��������F��������K��EZ@J$��n�.�����A߷�Z��#k�y����o��_'M��r$��!�)�M\缜�Z.v���j?�]��NH	+��Tܬ��T&�gH|�Y�;�(;�n�)Y�ޢ��tU��+��Ҿ�|lUH���H&1Δ���hX&Oo4^�Lq��P>^��<qx'!�NqN�燬����F���.ý� �[\�&d}�����R���B��Qɠ�M0V�}���ؖ{���(5��0�b��|3������ʌ�j�J�\�p�,�wz���H�+g�t���W��e�mY��N<���W���:֥�Y�ur�b��|O��8rR��GM&�4��z��lǃ+�h��ϝ���=b�ֈ�����FETiQ�&����\�Ye�Oߥ��o0�7��^�S)AO2��œT"Wp�G�& eZA�>��Ppmk�pXl���Ge��|�f�$����w�ܺ�����oa5*;�*��ta��� ���a�a��E�u�h�d��4=js�5��0}-_����>޳�J|;�#'i�t�sOa��b@�:���%�d�����W��)A���fy�~�g��|�y���>k���k*>��'�a�e���E)��wҠ�� ���'Hh��Bt �-,�}�2hW�j6W]�p���>@3�����9>���t����j<�^�X�"�+"��� �8d��S̎��ږ�|��\"�Aw�n�mO���z�����6ԍ��ʆUK�X��������Y�<IiJS:��WL����l���-='���b�
Dr�J�u��{�޽����P��\[��������n�����S�Zud���)*}�ŵk̛:�1�^߈��*����o%/�m��p�s]�R�Q�a�o/Ps�_y�Q8��Cv��qm����U���<�ˬ!�dQ�8r"}��^���E`k���9\�����>Q�X��tԌ�|��4u ���[ܶ W�E��QJ�\Ũ��<e�!%0|E��Oq�&�w�DC�ۮz,j��7�D����7�x����~�����x�!ZMHL��|��SA���8:�����8n6���ک��V
����2y��������h�!����&��'m�����;:�-:R�yέ8L \��I�u�e�d���N��.B'�?���,O�?��	1�zc�8��(�?#G@x>���[�5����\du+0�DW�B�l��wL:
;�m˸A������+�h5	p�@��
!^B�15[���[�t�Ł�J����&/B��V����&U _r\���☈���QƀZgg�_
��o@ſ.t��}�#�2�g����H��;� ?1oY/���P��ޓ������`��*�C�)��r�͑w��eFbϑ+�I��p�f���@���S^J�H"��I��or�{\B>+���I��Ms�su<n�]*����
�����F�tɻC�_����?�'�%�G���AK���ʲ\:C�<n݅�v�לɢ�?�Ԙ���s���ۂ��-��r�̞�o��ٻ���q�6��=�O������3z/^���zN^��p��Z�,���Ҍ���Y�RT���<1����Nr��%ҝX�`�"}���M���}-:F�=%Y�[�vʦ�Z�:��V�����?���`ؽ�=	����]u󦮳4��o��Β=F��֞@���K�I����S#������^
(D��������t��%�+	�'���һ�т:���J{��H���̯\WK`��!B����DX9 R��d����������$m���nD����+�m�}�t�y$#���f眽D3��&��ҷ�z����bi1��m��&����.�d��^�����W�1t�Q2)�A����\��"����"i%bx�ۓ�-�,����(p��&�H�ֺn��n)S4#f	�;��U�CJ�F��P�	��B�%,��i��s�����!xԧKǈ}ۃ_�_}���5�^��K (5�!��<��K08�y�iҽ�����Me�h�9�7+�d0j�o	�"t�'����=6!�^�T�o�2���~g�����O����Pb�|�P�8{�C��W�uнk��hz����O�e��Vp% �]��:�=����O�J]���k�H�j�Y��oby�кf�޲��P�n�)��L]˦�Z���CF8m���t�CӢ;w���V@$�~b��I:��w-�B3�����C���i�a7�u�A+��Z4��Q�H�ToE��k�r���vH.J�t��Û��l1��,X6ʢ&
ۆ��ߏ'��R��b>��!�[E��q�d�<lϩ�eܻ�,7[r���dWG�0iI�\�ދ���5�DP ��o`%�vx������x1}Ɵ�%��
�4<�-��C�CAR����`l���ã�{�jyH��+r(v-b@������_��8bY���̻6��-�+ bm���?m.͠�g[��+�1a������<�)�ߎ�.<�%��	����Z�I�������3Ǳ�!�	/�P$/<���:�%&a�_�6U)�!B+g�9^�r5�wZ]��ճ!�l[���ٹ��/�}��3�0.w.+z��'fcuRz�ߣ�5��LUlϚ��U\��*��P8�Z-�]�4���G�o�]����V$J[SO�����zC�U/t�j<~��l�[LkϏ��d���a�,wj��L�Ȍ�%�E�)�W ��M�/R��%Q/
���wG���k�����N�#/G��iN��8(�@fR�"��S�w��/d������V�#�
�)BϨ�r��W]:�+nT�~K"c�Qm��r�E꙾Iw3��\:Ph�¸Kyr>��$"���~���*�FĹL(����~�$����\��ĝ$wPw���FuO������:Mvj�挕0=d�'���e�GhH��ԵDY�_%_����j���/c���%��eo=��L#"E��j��-V�g�b��_K��3��%N�����P��t��Ɖ���Rٖ�j�O*An��0�Wh�f�Fs���ڵ�}�\���r�n`�%�c"��ӰāR�������������?�{/�nxA�L'�&Ô��i-�8�� ǍC[�t;z�9ƍT�(q5��W��޿���<��.ˋ��iA{T�rM `��qnؕ�0嗡���l Y��Jq ���@���+$�ɂ�V����1��s��c|��В(ϰ]'Vp�L������|��ݛ�)o���Ս���Q�n(�y����/��ŏ��L����7�,S.}ޭ�L�z��d�m�/��>'�k��^tپ�N�$�m�ۦ�mc�ӫi�\)T/�<o�\|�FL3�{%>��W`�y�<���T���-�A_�L���z�B�]L�n�?���E�%`��w��\;�a0�l�z���Y������9��ɷ#�v�����P�Iy#R�W~RI��p�^[���9r) Q=�G�><d�=�l���E3���گ2=r~L�fg��V��<BP�B�x�F�匠0��`�*+�/�)g�iC����R�a�[A�fU�j~��E���"�� ]��F󓕫���у��vr�*N���x!�^�0���[:�b��VIvtԐ�S�x�f���3uL�S!�*���ɰ��l����[��~�/�.���2�������<�Q�0=/�\ؗ�|#�M�'�W�S���	P'�m�6���!Q��j��(�	����Kk�N�0C�|�o�
fTtK�ԡ�_���-��ڜ_6�|F��dm^�q��Ujh�,t�h.{4�s�}Կ����9����XE���j�0ckϳ�,�|���3{æ}�P�t˦���R��ZZߠV�5'Gg�T�۞��9O
nS��,�J�s
�>k��}u����9�|���:Cs�|�W���t�n#�^�����M�X&�Y�����Fn��R��A� ��,�1�ާa{���pJ ^���Kk��F��� ���toM	|~�1~�Q��-��Ȱ���x�+Ջ['���\z��sq�����E�\٪������k�sM���h�4K�����S�BIh�+��O�cCv�e2CS���42uĜ?a��$��+�$�m�h�B�z��g6������K�XWQq�^sȅsB��|s��6��fi�^f��52k���'��UT����rsj:w������=btlҐi��Q��=�G�����"*D�q���e�K���KbZY�t�r5���%dRtXԮv�s��Ç:T���CR�Ԯ��������3@�J}���`/ۜ���@^��H'Jq�Hiw���$(��ai:����Y~��v>3����5�⾰�(���������B}��X�tVq��̅*SM��I�]M� f���f���Ք1a�Տ^&欞��Y��1��qz��e�S=���ao`�-⿝�!����T9W���E�܇����/*���Go`/���B��5Db�+ep�J�|�k�]0��{�[CJ�Z�A��T㚭�?�^6e�1:�O��9BH�0^SY��k,����~����V��n�������A���m�����r����`�f�Xߪ�z�o/���6���"D�H�[o�|4��s�V����Z<��ꉳ��z��PV/�9��J�TG��޲�O�X��an��~�l��[� u��W1A>�`W�/����H��|=�t�q��Ԥ��l�"FG����V�"��������q�}�{z�-�t��#챤�W�|_����l�s���T+0
�`].y�����6�NͶ�;+d�<�6�y�)����M�����-o94���r`=潜:�==����\���C#�)C��Ǜ�U�F�-FS����°W3�|b�<�
��fbh�̥�^>�z��v� �Xq����yO*�p�_XKm��߹�(1���Ɗ�ׇ��ґ���)^�A��>�Xx^8I	�@H�>y=/�x>H��z��ޱ�v۪4�(�Wz�ٔ�>��(�Z_؍mL�Ҝ[>} ��=&�ށ|/?}����=�{`/�i5����M���N&���gظ�*�a��j�h�zę4_�vf��d�ƃh`5��KΨ�^��'���dy���rO��P�Ì�❑>�=z���'�za������z��� �4�b5	��ͪ�{QF�{�*��/�D�6��̙�\T���p�g�}8.,����Y�1�/�^�2اX��/9R*Uxʤv]kW%��~$�}���[�/}W7����;��*��>	�+����'T|@��T��������|U���&�M;X�+��6��{� j(�w58��R��(ַ��؇��1����WfL>,ߑU����ﺜhS*����ei�r�9����=|�S`^	�e���,Ӑ@>�+辌����RR���͈"�[b���הH������Z��xfr� ���G�`�y��V��T;��+�i�X�J2����<�����5��k_�?;z��.�u���� �ø1�^��߃�����3��߽�YE�('W�����@����_9k�iqdڈR���$E�ĴAC}�*����ui��j��j��V�L+����~thq����	�|Xo������q�R��"�UlrY�n�M�kF:g�@!��L7�h��_s�����C����S�ʕ�������C��aƚ_M�����1���$n�y�KxR�:�E��SS;��=T79��{}�|Mҁ�,����:��yv�r?|3�������m[qwx+�a��rF��E�g;	L���5�$���v(f7�Ů�s�p�����']��#~r�t�v1���5 D���ާ�f����w��f��mҦ�׭��6�z&9�w��wS*g�q���b�,QQ;��92PGW�0`�8s�;�I1�jgʖ�6��ʂ�ټT�pbs�D�D��@������qf����,�Ʊ���?K��G�)�^Ғ-�\������M�X{%C�r��6'3�ǅ�d�juN������d���n
<^��ȧeǗ�� P�����q�c81�q<s�f���S���1'm�`�1�܊�"�	���TSń� ⾃�`מ����&z�v�����l��$���I�W��k�*����1��@yZΑH���Wia�g?7��{�x����J������[_��6MA"7��M}{�/���A�4�^��=kϰ��bz��z;gO��4��=���#0ëH�����k�]20���_a��D�g��u�
�7���ٙi���Ov�,5��<�@׸���S���U�2���D���ǔ�p��,S��^*f��n�C��Ȃ9w 3�q�M�/��Y�~��Cئ��J�9�4@��
���\���R��$͞��j�Tٯ��6Uv���h�P0�e�K��+��zUV��Kh��ǫ�I1tC�F+x��oҀr�l!�Gv;���2=�"��?GD��	8|���_<��%7x�|�.i��%.�PW���+��_��&�	��tlK�f��P�k���&��%uqɬ��Bwr��ࡕ���X�䅈�W� �N������o'��!W�Q:�=A,L��aG �*~#�,-���#M�Z;�D_��e�s�#
��|��k�Yl�B��|<�͍��?�[��om��JկWz���JT�����1�u��m���8���^+��3�|�^G�g����kM*�~�W�~��y۶Q
"C���[;^��6�3�H"St��E�d���
���ܹ�����8�/�R�n��������O�� r*�\��L��>�z���ZHjf�����ł�d:�/�?~�s���������#�Î޿~��^
���@�g*0��li�"�-�aA�:3�0�Z<v����g�qp�� f(%�#�7]�}��0}���A�k-L_D�Bآ���£Ѭ'�fn����]��:����h�UQ	��F����ż
�����v:xr�,�^_�r%Ī�2��PhÐ�a�QT�C�{ԧ��В�<��B}�r��a����vȌ�%�ͬ�iv�m�hE5#+E�(H{!��/��ص+�pߌ�k��s��d.�ʕ#]��S?"}\�1[�ֶ�=��ʢ/ʜ����&�QD'��&WnX}�x���>��0]�m�< �w��#��	F�;�藘�;�>��mZ�m?q�)������n���L�C�1B	��uN���{�B��� 1:��7���-����{�w`��e��~��X";�$Ə�����7��:�c�M���^dQk�a@V6p��r.�����"�&���_����%d0�:餪w#���\�O�jp��JټBc�y��l/{�(��wӆKpE�3���QbqV��u|)-���ܰ�� �*	n�*ͤ�;��o�� ����e)�JyF/M�U+�>�U�<��D�M[� ��.��4�՚$Ж�FK+@��]�S^�я
��*��ҵ��q���L����7ez�:�!��-(	����/�,���ը�蒍��{��I`7��h:@�r6τ��3P�q�n(t$p��<KL�`/� ��rä�~U/<�DW���Co:8|w���l�b9�D�±�xk�[�)��]�"�	��0�E�?�T����H���?�ڸ��(���Ip������������Fb���$f��B��,+@9�Xڕ���e��Ĵ{(��ϋ�ğ�+�i�s��F�U��g�>���+6l|Xe�TE�׊u&���>�n}H��G�mn����������lY7X�WNEͨ抌3W��^�.Zr�����a��Q��ވ���	�Py�����������"���5]�߉�n2^��hy�F��������i~��!�֦��lS�.}3<��p�;r��Q�-��'��qK�sV��:G-���er5^��s�g�C��j�0�Eg�q���hm���4�]���f���U"[܄w$�c XȄ=쀥Ό��6;b���F��;5nϻZSE/�I(C�쿋�}�Rr�$�~�5�>dv���K2�XN�![=�:кC&�^� ��>f�D�#B_�ǅ)9�&�k5�Y�������Z}W���&��rfW��'�����vP�Cs�󰙄7qL.ю���r���{+^̛9�;N\�1��>����nЋ��� �ے���u��6���#0��{G`����8��]��F��XX/��F�#Y�z���T�"�[�C���T���en祶�!�>�>w!}8�Oͬ�K8��G���5׿PG���0�;ˁ�^��Y��|D��tt� ��I?���7�D���K����_���3 ;#��B� ��ײy���������a�o+��k&e���U�'���Ŕ� � !�6��a��{�V��n�������o�Œ���C;|�$yr��}3��ے��Tp�!Y!�nD�㬼�;u�2��}��6�D�8pz#2`���iXl9?^��Ս�����c�1iGm�MK�Y��+�����P�p��
~r�9��sw�IqQ�`��c8�g��k騏�W��{�/l��w@�x�?� }�B�Qd���dg��w֭:�P�¾M����yX�¹�̗�>�-7��x��G���$�sa*��Dҿ�ߕ�7�ymq��>���O���~���!�Q&� �����׆��,�LoZ�h��}�����m#
N� �)v�����:hn�k��_�z�c��6,��^w~->T���k�3|,��=��k�2�w���u,v��^��a?J�N@���.
|y�H�(��x���1��d�v���	�D]5k�8�r���{-����~ �wJ�/ƍ��P��t>]0^�k�wS�[���4����E��Wj�#��qU���_�3H�)~td����4���<x�_��`ۻ����a���� N�/��a� ��o��>]z(��p3Km���c%�������Wd�ru��3���`��W�J`%�8Z��������d��4u��(�NV �2�q��|Wz�L�TkF ��ğ�.r�����|�y��=�-gǭ+��p�s�'��A#�(����w�y-�2�����̋�u�KGUF�_q�,�]ހ�?|�[��\΍��|����Լ2S���m^9W�0�f7��9+�g�$D��}z�(�E�6�2GB�c����D�KJb��d���{ ��n�}����׿ZL���%��c�3��� �X�*)U���At��u�h6Mh��4��Cs!������I7k��'%��Q��|��Z,�)�}��f+�{������q����nL��~�[���*��P�0ZY�������_����p%�V��x&W�X�P��Fhx�Q�j�6�9�ˀ�R^���>����|>�@�S,����C�'!# ���ފC�Z���y�G��^I��=��j�����#i6�3����g��������&y�����n�t�@e�k����>[6O���c"��Z���tFz�cR�7t��p$�k�	�LK��x�gAO5�����'!����mf��-��bf2�2�w��mȬ��gѻ�i��H�[�
��X��py�ز�rz�v���+5B������P�'q�~-�w���A�s�P*�La�?Ғ-U�-~:L!>���n���	"�D�f$o��2"'V҇@J�� �����)�s�t*��K����l�\GΞ~���˞��D��X��h��G�|�}gw�~��L,��KK��*�Rf��c��;Lbz� 	�"�[���W,����Ȭ��%�_2c���<��!��w}��_!�;s9��![o�4�yXg�O�[ٗ�G�5Χ��OU�zB�������9�+E��>��^e&��f ���+W�ϴ ��ȵ�^��V����J�(�=����'����i��r�q
�i�u���i���ᎊ�ٙQ͜�Ff`O����|s`� ����[����w� �+`کs�}6���!��e���w\�?�C�@j�:���D�ￅ���������ͳl9C�	���/ݐb�{п����w��x��o��:YD�"H&�E�HJ?SMq����D���#�4̿S��H!��
�(C���*H�
W#��?�##�1�TyS�v(�1S��%n�3��y��ߊ�#D0À��I �3��k�k���2�ϵ�����~����󌚨RwP*���}/�U��͈}��DEG�� ��:�*�APejR�?G��O�%ܝ�zU>"Qԅap,�`���s� J�)1i�a!�7��1�%P�=f����^!���x������$�܄״SlX*�qOP'ܛ�7�[A�[5� �Ў-sf�����f"��"hk��=?rb�@9��8���J��=���d��3W�ڙ=�L:{&\�shA��&�#���$���r��G���(���c�V��y�����)Y�P�Q�s�]3�N��'�9�_�6{�>kź�*����gㅗ��J��j���naN� KE�8!��KfkW���*y��:��l�)�����y���y!�'	f��6k�[�c\ys�Y�$��Ap�8|'EH���z� ����#O�&|����q#c̗�� l��<� ^���?���6D��f�$������6yG�Nzگ	�R����@�������i�hE�[*�B����y$Yh���.X�Yp��m{��MV�鷃膱}II�H�-�AH{�V��"S��yw)lo[!o���H��`��� �����u���0K03�
��'�+��%����q����Q��t?�������3�o`?���a��;�`!�>���a��=g=*������ߙ�c�۬��>�Z��}�͵���{�%Oh����lǷU5�����I���g�6��(��Ǐ�L�mjj~��$N����W2���~�#�i�f��+&��ⓐ_�u�Zu��tj�g�R�����]��\Lf���|�\u�;O���2m���/t㩤����-B8���l��r�O��=�� ;Yw��w߉��u|!��nmcZ���E��t�@ő�@cǊfs��?�I_Q&���_���BT�	\+><G8@���9�Q�]���<*w�D�v� ��^�T�#D5-�(�8�\4T�0����k�w
 ���ް��G��Λ��{�=ʬP��z3e�j/�\=���Ĕ��'�q"aҚ��}V@d�c�+��#K�A��\9ۦea] ��I_=4��
�����.$叶�mqN�/8�x&���`x��E6޼�&�ٚ>�0�!�=�/7�P�#P�hD�É��K{���ƅ�d7/�V��5�.ƗS�:�	+���|��Y�c�%Xyɇ��ĳ�d:J�P�0��������ߣ�81����c`Oj�*�W��:�#��>�q=|Jx�Zw^c����N�>
�C}�	�@��[�w�,o\���T�M�IP%zϝqm`��eC��O��MG�WTF�8�'���=m��;ֿ�x�z]����:D�I�/Q@��� �~�@"��TM�DP�4,}�\��zDTw�w�4gC?;�DK�}8P=>H��S7fL�����_L�H�㺗�a�N�q��8ky��s/���(�e/k!v���.��ueЯ��w]Mo5����S����_6<r�eM���~&U�
J@�I@��fw}ĸN���5L-Ť\��c;����5U(p֐4k�	�3�G���:������"PIz�]����\o������N�N�U��yw���q��^M�/�@a��k�e9��@��1Y�zz@�ҁ������	�+�UBj���#ƕ�1y#5"�ѭ$G�mX�Hо*�W)u��(�X�k'�s�2��_��� h�Ј�ʓġs_=���ύ��ЌQ=�|*������[�P���*�+?�q��1g�#������?S�?���7�
�}��^Xx�B����]$IS6�~�~��S�ݪޟ�?��C��N��N_c��f>@
Y���=����s����E9��o/@��wb�A�7��u"��}�j��?�ɹ�+�
HeR�P�~�(5�x��/��<���E����3S��F�&D��0&��G�d��F��S���W��o8�H�ڀ��[�t�;P~9sm�ȫ�F�_�6�jǝ��YW�nB��\F�[�����x�Ᏼ�%�< E�����#y����O�s �v׷��,���ɻRh+Nw��+������Hţc�}�+��i6,�.pE\��]�ݸ6_��q�Z"�W�Bj��W<W����l�����J;R'�,���b�*�����~zQ�Z<�z!��`����L��tI9�@\�h�:�0�4�ѤX����z��A��� �j��Io~#�*�����L�oY�a:��������.�K�� �DO�~����TCƂ����oU��<��-�:B
��v��iZ��Ιd�p����I*~�a0��Z����Փ��`�u6
��m-�������8 ���N@z���l��`��1�	
v�y�8�x����"-y�Tk�,���Bez��Y+%:��v��I�!������Tr���zFl8a5[��t��g{��"�ݹw���_Ú����%s�6C�R�(��lfDc�������>�l>���?�;L[��(x�7xC�w��]↕ܼ?P�E�\����U�02�j����1{��ry���ʝ���M5��涷o�`��A�:�i�l��y���`r�Җz`����62���|?�G���S���r�p����P��l��mb�j��0^�I ^R&���J,'Iy�z:9q�]]?��lph~��Äd��ML����U;�(��E����~���_��%���h:�5P8 �ˤ�@��X���BF�r�Y9}��ghc�o<��f��̠��6
� �}�$���e�Ђ��e�B��K�j��?� x�ƟnğC�>u(�e�b�U�a*����:��l�)Ԛ��Zި]�U�EЬW.��qz�B���!ί�̗:����jo�}��Ca�8���ֽ8u��0%�!�.���hB�n�o����ʱ�>����{�_�Έn7�G��w�r�i��G��$UN������}�#�e:���!�xs����\����e�2���J��"~):�Ď͉Q�����1K_7�lr�odkmy���z+FRa�餵��^?eҭ�!�s��w�֦��\���M��X�Õ�|g\��p���3xSmί]���HFa��l���W?!	ds�D��ꅑd�PeVS�V��3�x���@�Q���џ���[l@�e6%�-�Y�
ж����v�XEn�$S�P�'.�և�iHݦB�ޝw�^�� ���Y��18}�*��W�:2�!�S^m<ش�~SȮJ��5yGm]+�r���Vo�A/ ���"��"徭#��[��I�K���	 ژj��<����kޚ>���E^�?�7$��T��ժL�k�BHʎ�Y���]��-��&�N��E��Hʭ<:�юF.j˫�X���~��g,�*��9]�M��i>��Y#D�޲6�4��n�� �H���� �95��딒��+X"p8/��Ҫ?�QP��e����������ҍ4-����M���)�E�ځ���g���I�PS�L���2I�2�D���'΀�� d���OZˍy)��\���f������ut����TQ�� �-.�ǐ�X_Q�ߴ)��c<���P��jVƸ%?����K3�����B�aqH��'�㔓U ���r�H$�5�^��A[ =3K<�v}:d��_��茙�FlƋ�5;-�>�;�K��J�hIc��Jk��Z��6���*`2��_#��<!/��#�.�����)d[��[�J���pJ�ym�~|�A�tK��);����ýg�qEKG\Jl���p�If��ꤕm\mF�|����Dꢴ����ͼR�{����bb�k��:��_�{���P�̇�� [WZ+'Ơ��?F��h��,�T�˨
������:_�s(��V[F��ȇZ�@��4���!eѪ�,���/�H�X�@}����.��r��V�ہn�GRl� �j�����襦��*���x�ﷃb_:f�'��1�5y����>�6 ?��b8OQr�$��h�ᾪ�ϙ(t�����W+w�,/d�e����%��Z���dZhm8
]��?o�����.0���\9o�c���͔R�����p��7��s�zoq�-�	�Q��.m���̳h����qHsnY�Hv}*�g_��DA����n��C�7_�ZJ�j�7o����X�!�@/\�ry��с��w���<����L�0X��������J\��$:R�и�F�:Qqvb���#�`�l���_�8�X��y�0YD#UiO9w����Z��ݜ�|��Ȁtz��Q�-�x3�n �GwqW(h��]�T�0e��i)r���c����ed��	���gS��l�y���5E�3FV��E�b�[�N]ɇdf���̙š��G��(���`!�GDF��q�z�)B_�)w�̲����;��j4�!ߣ�g`m�G޼�,�n{,d�VjͣM�X�1�44WmP�e�
V�G�xD;Q���ZW˨�۬�w2x{[���ٗ\Ϝ��_�՞ύ0-�5X��Z�ԭh��̘�ןU �'s)�6'�4|�Hw��r�r��t�ǟ~T8��?���w�qX�����&�eR�Ȱ+��I�akZ�
��nэ7�W&�CbG�IƄM���\����+��-%o�k=�΅�|�	����L��mo2�"�(ZM�/�Ӌ!�O�8t���$Y|�/;���:r2����H��1�\C���u�E��L!���/Po�|~���m��B�i_*d�f��-�N�c �J���|u˔��ۦ���V�<�@G��5��&r����<��mq�#��^x_��)I�2����z9	��7�7P,�z�u�yx�t�Q�6�gr�qB=L���% U�,�,���:�:�O���՜_���O$��bK=���M$I�k9i�;0b"���7������?���+�Z��J�6����r�5��w+l<�>_�T��lJn�qn�-}�\��E�G���ƍ��J%�c���H�0RJ��5_�c �WY#<�؀�pg���|Ii���61͸&#��tC����߳�u���g��?�*��mw7���II�/���\���j֯
³����Y�oBP�;��ބ��E2 ,E@�2./��|/t���N��<`�*	b��Ś2z�l��8�$u(�P71u�/Qj�?z�=��Ӭ�����tk �UX�oӁ�����,Ib���P=DF�"Xt��FTuE��`�rt{�K6_�[{��}��iZ	 1�v�|����+=l~�jv����ߔ_	�m��2g���eI����Y
%ӥar�yK��	0���zzh��(2�l��*�	���ĥ���+uأhz���+8���
I�#!�`�$#�_��@�{��y�f�j#P"z�%��OF�SO2M?�y�J������5��N�N�(�ϳ� $�U�X�d�\W��b��P��I}����֔���wl�	�!�f������f:���t����D(Fܰ wW��窬�gs5�,	�^�Z����f���;к�o�[�擇a,��Q=�2�Wc��<��M����;%�	�Y�,���	ލ�O�.���;�΍Kv&J���m<�wN�1E)��̏���J����t)��(e�{tqZ�N*XI�B;�:J��z��± �D����1��K�;p�ƆK��y?���"��'�(�-w�~���lX~�|���Ȓ�e��������(r9 4�d)�Mp���;L���az�&~]�Ҟz�!�������Ggj=���7n�|a&�~بǉ�<38��$�Aǭo\.%��u^iW��JP#?}9`��ԝ�dF�[��6��@�Z3�{\Py9�@�7jX-꫋R��ͅ)��H84�T��������c�-L� ,#?F7��)���T�X�J���"��l�~uj��{�a��D�Ď��fŔ��n@��9Xc��.Ǟ��,��~U>���)�Tр�aSʜkډ���[��=��i� ��.ǧ��A��|W��TI&��-+��+ ��Y�%��U�TT�LЁ�+���x���(������B�2@2��-ǈ��[Bp�N�q͑�������M�Ӂ��/�@��qD�_%�K��T"}
��G���I��ef�j�Xyw}i��nW��A�,mS�o��l��L�o4�qy�Dp	�[��ҭ|���ˁ�'�ߦ�K.�M�?�����WC��!p8�D�9�[�p��!j������]i�7���C�����Y�D<�7���Z� ! �J��ʂ銒��^:��x�&eǚN]��:+/g�{bȶ� �mL#m��}z�o_!����D�/t��*�����s+ˤV���'/&�V�_K�55�ej��H|/[d�Yz{��ǝ�[qv,*#���h6K˗��B3�؆�^���R߿T�[��홳���.���������A>ws$��eW@r������#YPs�u���Un"���y��~��.�>6x�66��4��<�S^��R�!�����f�����F�&��J�k�o�|����9���G�g�c���yΑ	Hf���QH�������K�/���q���M�w��� ����r���Se��@DX�x��aH)�դ��JST+}`ɸ�W�oʪ9�L�:�Mq9a��猴��4@|�Z��[�W���A,��j�.J�����x6��{�X��y�x+�A��-�צ�iVB�ؑ��QC5k[��z��"@�����n׌_P�����stPu�˔�����o(u P%Ĕn�0��nC��D�#����Q>�'�V?�%o���/a�:�JX535��j�ؽ ��y
�=�����j��h�R���t�o���J�P]��}���<)	�[Y@NU�� ߕ5Kz�|�2��O�'O&]};�}�ˏ�����}īE6�,���O�Y *X�o�vx�2��h�O��V|2���%Bշ����``����N9�`#Q ��u�j�Ġ��tDK&M8���T:=)�	J�|X�VcF�^YGʂ_({� d4	�3(e�����$Gʩ��QI��1)yUG�GT�x�� u��9U��e*K���6P�w����C>��Pש��ֹ�4mg�'V��.y�4�L#�� R*<c���g�y��d=G�������m�fږ��Ҭ�B:8E�+�5�ì�G������aQmo���
�������H�P*�%1t(�!C����HÀC��]����0=��3�ts�&�����y�X{��{����؁Q idpw�	z*�O-f�S믷x�N̧��$���G�3��2|6j�z���_	ٛ��O^5�4��R�R��L�s�2�B�������V��d�y/eB���Ǚ��0�j$ ��ar��](�]�}�~]A]6|xz�I��m��?���~گ�ˣ����lbS��i�ʗ0�A�!Rm����<A4��4Pwf�
D�}�_�K^�0h/-�v&���d���[�̉�6�"��B�']��2�����[4U�%�H�u]�GRԵq��A[�H�φ��a�a�^mF��ۏ&����؁iƖ����wo���#7Mҥ�ŕ�;^r�M��0�[�^��ٟf�/�!�(ls�[���o�V�����Y��H�o��.zo}�2	�d��<���ʙrI�^�V��^ۢ�ٌWA�e�i#o�԰Z�ln".�	6Ԓ���hu���˚�$�ԯ������pA�ű�v�t�v~���m`�!,ۊz� N�f������6t~;FK�yH���÷�M�|�Ӌ�b��Y�Ǽ�_�_�)�D�Q`*�^�9�~n��:"ۡ9���z Ù -��I���s�y/n���1�*wt�,��V�q7��(7��S@�GF<~ ���8NV��@Y
�k6�������1�2+��"���MnWj��d�y\��tu}�5�N+�}C4�7.|~�G��i�2��^���)�e��2�%��!�֦�S /B[Hxmw�4z(�K+�!VI��X�;O]�~��4��N����������9Z�ؒ��hni
a����y�r]������B+����49�Ia���`����n&�-��ߞ�ˏQ��H1�tv�A9��/̄*4�ī�R��wT��ր�\ �e1䇾~����͏�5�3&:2�+C��LVYLĞBY�v��=d��Z�_S�z�\��Q^a�� *}��Gy�S5�ꦵ�e��jZ
C]�{��N����M�7jq:,���
v�g[Xn�s��)�h �I��j�.PIb�-G��L����>�Df7�q'�v��.KV������K�#�Z ��,��k7�>�g{K�����$@�P3��e�vuq���<��HF&�^.x��&@K�� �| G�A�-�`��'t�r���)��3�c��9=����:M&<a����ne����'a^KZ�4wFs��p���8���%TA@^�Ҁ&��-8�fG\�I ��
]W�p�V����}<�8a�U�-�w�6Lkƛ�	� ��B���&�]
~�i5'y�!ħ�B�4f� s}�� }�&��ƀ]�|��Z~���7�qZ�o.xF�1woߒ�A��'GH#����
v�r��:��,�A�'�e�?CE֒�����׮���xK�bru�h��T1��a���U����w\�!Y/%lB��\fn�ӂY���N8�QhҲ���9J�n%-��?��k2�W5� ʢ|�#��\Ѽ$�B���̈%��C�xԜV�+]��`x@P��ߊ&���)����C6a��
I^�
����	}�#�B�&��s7�Pn������a�ҩ�O��jn���N���{�B���m`��}�����S{���2��l�!ť�U�U gw��t$���&&A�?"��,���P�2�KAN~d��������֖�T�S�-��)�����#�ՁB<�����ԉ�B��N�a�k�Q�l�2���n��cy����\M�K�(����їB�b����S��Yx���o��IY���y�\��|m�Cl�;�Jæ�&���:��Ws�/�ȝǣ��tBū��1}�o�����@L(0G:Nn���3A�e�)�,1�n�.G2��  ���c.�"��b]��Zo�[��K�¥p���V/��J)e�(�~T���j������rW�,�u.�v���fY�qS��^Ļ�J��V����w�L�w���:g]!�!�d�zcg-�	��ڸRs4!X���ZX�FRy�UT�����s�̭�N ���tY� �:�3�8��F2��������m�x�=�5e�K�gk.�@Bgj=5���c�Ϧ�����d~�Q�\Ϭx��}%1yݔ#��>�e��jp�i�a���^�~�i�{�@��n�]�UPѯ���X���6'�f:\����NL��M�|&�Jt]˾��2</$��s��AH���ڳ������r�O)���@ql���?j �7�i+ii�6b�݈��ޤ���i�f}f���~�UſU>�ŷ�9�yF���] ����h�0�	�NE�s�ګ�L֤��A.M���i�"�x�>u�0����*=�T��N���4������a?(�
� �ycQ���|�^�q#�d�GZ_2#���DA�ƫi,j��	��#��8?l������X��BVY��/�~͉ʿm�������ͺ��m韋���}��<�z���!���Z߹)���^���(���B{����c|��D���_���$�u�`�hG��eD���XwZ�|��4��I�e9����$�M�����F�W���67O ��=�O�=6��Lqu�8��㬈"!�h.��nd��O dO�U-�4�z�}ˑڟX�)�k�D��]��*>Y�َ�J�����G6���aUd#w%����3��+G����e]����u�׳
�{�� 7)j�D.�D+\zטl7ݱ�a#e��=Z(gV��Ί���j!�]	�NG���8)����U9�t/'`O!���D��B�L�J����R�Cf-~�qC��^��5ʌp` ���C�]M�����3�}��5����'C�F+��n�����8���V��p�B�\{�rX[3.�b�$�{L@�!Kyf8C����b#����G��zHW�)��!�m7������Л��-^ޡV^�܁��ߙ��o�s�N��$��ywL�D  ���!HTTs'�����m�f���̂A˫b8�� �g~�\�j��	�Η��̔9t"^�lb�MJ��1��v�P�+���>��bo�:��~&���븍@4R� %�Fe�̌/.agC��^d�g둺*���M.��䣕�4T����6�:e�<O�>r�{�ސh��<���K��ۣ��P���2�-SJ����Z���ʵ��Ri�$��^��^���K��C���"G�,�O`�ˀ��6�g����ܫQ2�c�o�|�s�X�b\<�m���Ya�~]Tg�coo�%z��	��LW"��QP�ȿ=�f��;(ߠ�JF�v�?��
2�/<��_ͬ�F #V�?���s�����C���n8f]��
}����\,R�O���eɯ/e��G�~�2�s����o��'pO��F�����]��"%'�\��P`�K�'����O�����Lhh�� ��R�u�JcB��r��8 ![�g��{�<F+@��r��S�-}ju�~��ZWL���v�fv�Vv��܋�ɻ`C෠�<Ʒ��d7����>��d�;-��NH���ޅ&}�;z ������2�����Q��30K�JEPb��Ml�����~e��٠��/��m�T9��$_��366gJ+��M�7��!��(�꽅&9����O�,�MK��A���_�zˢC�@m��Z�fue�Is��}qң߃Ҭ�H�2�c�5/:{��t��˗38�0V�~|�Y>t/�ƣR��mr�8szm���C�0���w`\]��:t�K���7d� pf�ds��tĝ&������d�7( kݰ��i�J:�}�.�W�+���p B �<�(��}u}j�O���^�U�Y���=�l�����|W,t�K�#�`� C1�E_��B[u�6s.��uN���'/��S�h�0�{#%i��2;
Y%\Ԝ�O��p�x�&���J�ji��	�_��X���X�dU̯{�;Py����	+����,2��VP�Q/@�P4��K�i�C�̡���{���� ���I*�뜆0i��-DQ+��b�4$0���2����t���^��ɔ�Gv(�c��+�3õ �9c��̥1]�+��~f,�4w^�|+%�ꐩV��V"�0��]T�Q�R��o(�<i��6z���� Z�	��B��?������^����1�GOw��϶b���o�ӿ��1�����W��v�o��dO���R��V��]��Lv�$�����˶C�+K/���[W�ZP���c�Ĺr�)�%��\}~�	K�L�޷�/��� Ny֩O��Fٕ3-�T�vSV�i����Y�f��_w�)��*e�����
o�THpg�D?��b
o6dog�\\�e�G��~5�^^�H���P3����,C~��#+��2���������:ɺ���#���"�TF[��)��HP�MP�Q��G�c�P5�]XGe�xFtZ4����R�K�URs�M<���#�_AK�4�Y���Ĭ�,��5���g�}65)�����
�[ϗ���������ul�;
.ɯS m�P��vW��OqL�z��e����!��≯�s~�P���R?<U �/�e��Zݲ+2@�\b��=�����}��xֿ�g�C�/�%Z86?h�9i{2S��BjB��D�=�����J�̱y�J��Nz[p#4��-L�&�����v��sr����6��,�owj�F��c�X��D�?�Y'��.�{�����uc����r���h�΍�U�)D����=�@�.�z���*�#+zMK4�T�b��9����Q�V��By��Mu1��k+dLŴ��X���_E�Od��ǕCy�|�`hbTȧw����N�����@;㻔�3�;�P�e��
��WE� ��w��٦&�V ��鉫9�b�i�h�����--�qG���M�T��r��bZO�Q���fY����n�) ~S����������c��_#�̑��ue@�X1�`8!��mfjЙ����8bAjUW�@L��n����чh�H	��aъ �m��Η��ű[t� ��5]����	�p�oi��0�(>�Y�M>�Ө&�>~�Tǆ���U�~XR��0�A!׏`"�Y����u�Ǧ(��Զ�,���6_�(�ң�>�_ #��L[M�{�U֣�Os��]qͷ�̜�^ϐE9-��.D�+8�b��`[�r�� 5�xB���|�3�|�9��]�}�V��x�-����ŉ�&ɂ��r,��-zѾ�./��di"�L�#�`cg&c�^���w8�=�?�I}6U�&*E��M���C�<Ccm3'��Y����3�a�#��O�󴓀�&�Ԕ@! �dX�|'8mf�[����C�$�Z~��^lu��S�p���O�����n,B�	�)RF l��F��V�4�B�@��wSi�^WL۪��g��&F�_��<>�[i�4Ԙ�R|ͣ��i,��G�]�V�� ��8�#��2���]j(��4장@3Ⱦ��I`w��ˊ�*��z����I�n�^���HF4�W�xU�m���G�N�mH�V��#ˮ�m�7\�N�Z��UZ�堲SQ���o��D6��c%�nS F�!vǹ��W��k��39i	o�O�6����R��H2^�{�1t)$�������{�!^�9��F��~u�*hw���ж7n���"�!��iX���`��f���`���uh��@�����u�j��-՘I��݋�����h��j���puR(�cT���!�|�r�:Q�E����}UX���`�y�{w8�f߈�!���X��2�.K��x×>� �q`ˑ�莱�>��7�N����܈�	���~p������i`�����Z��J��w"I�W�ࡀ�u�EqY��=)����'%%�[��syj���|����X�N���
׫�I����gfN�%Aܐ��� �0Nu�~������U����f[� �}D�eok��2��K�5��g��:lB\?�x�W]f랩{���H]ڪ�k�c^�0~�%Cۥtj�+S� Ͽ# �>0O�%�W�5��6�K<�!p��=�e�M��ʹ6����jn�{���RG%~�ٯv�D��\�x��?܄^��Ǧ���#T@8�!���=�+��VK4��WZ�yRe �R#�����������V�!.�ǽ�	��0D��ec�pC�@K��bƋ|I�	�D�*����[h ��r�z�*!�;Җ:Z#Ӽ�?�F���c��5?�U�{\q����!���;��@~�b9@���*���{qz���$>7�Yxt��'%�9:�&LP�x{�w�Iі�n��ۆ'�VН9%tߤj�=�yϭ�h��������P_=~c8�D>JV|yW�։�����z�`��p�;�k��\�%��>ư����rVݞN�+
�T�ļ�tR�x��և�Ȩ �����%�2��Wc���c�CR 7�hH�|��͢sb���!�>H�s��/Y�'5k�F>��<�{���ދ'���N�^ށ�J�?��9(ޏw¥��0Fڋ� �a-f�?�q�F��t|楓95���{U��>�T/V���c�7��ũݍjY�����3�W�2�� �Ats�&Y�$������ڔ�Iv�NO���L\Sɵ���5⧃O��񉱭�n���]���y�v)T���	�&��y���	8�/u]&>a������3tC�Pc��л��M3v�1��������Q�^���)�K����cܞo���z�f�{�񿮷��N��^�[�~ ��j������ﺇ<ZR��ƨQJ����!��/�W���$�X|uWu܉���h7��+��o# ��6��C�90n��۴>����̲<�צ�����lqf8 
���(3����M�2��w�O:��nf�[�WȢP:9�lT��d~�Z��];�4��H���g .ue|g�r��NC�d�"��r74#7��b��U[�\ݺ�Hw�Q��a�l �@��ۂSȬ='���y�����f~eO�o�x����R����ѧAV���,�ŽuJ��t���e�)��U])f������u�͈W����x�~&��-|�
_�b�L�Ņ�ҡl��Θ��Ǳ���^���6s±����2�����/;�C�2ϛ�w�.tM&�M)UJ��m�ـ�v��F �}n��*(��F��9/��l5&99�3z��gf�nf��
2zkV̜��zIJB�BT�!�N8���*��.�n��'WZ3C ���봛��N(G��m��3K�X�#�P��_�<v&~S��G�hD��|�i�F[X]	-yqz�\jȣ7�p�b�zg��(�gA�K�u%�F�:g�QjϞ�<�����{�kh�VZ:���{\~��e�27݋�;�|�#;��Y!YA?�M��=Ų��I��!���������f_��!0�7�Wk��|z��lPh�_����+T�i��
�����ƢZ̩5.ɿ���z�r��G㖠�Q��W`�`��9O��w�_���]�R�UwKF��ɢ��	C��b�����ː�X%�W�bʉ,
_����o͈�
rg6�}8��������}͊��e�fH�H3
:7|3>V�4>���YW��i�5?;2��J*�&~BC�5�н����%�k1J~�9:Y$�8��Rʾ�j�B�'7�f�?F�狚w��)�|1�x[����^�y�hN����}h��U�D��1�,�j�T����{�v@�0y���R�7��P�w7~���o����f��  Qu�ˋ�����2��G���I�	A�wt�#�U�B�6��\��w	�^d>�M����n�����я[?�3�˖�Q��ne�Ǜծ��P�R��K��F��[�M!�{�sY�B/K�G\s�եj�LʄYѳcY$����yC�G�������(�>q���(�ݩ�6��� d�~˞'��T3g�m�N�dP�����z[�G�Yxk*�x�̚�ɡ����S���G��V�l)�o����aދ�	Ix̀�=g\
@$Nh���t:�� ��q���l�����I'��.>�3RIc�t�c_���5�u�����Sf�ben��Bǔ?�"����ٖ�[�mv�x]}�T���P�~�i� �G�u���]</�υӦ�����
���^q>��ƪ�}���Q�)е���L��-�����)��%�M�͈��Y@(���B��3��d����)F�H� �g${���'s���`"z�����v���߾��M�{VKud�>͈ ���y�.Kq�COE1t�'.���Y�:���ʪ��2u��ZJ�랛 l��HhU�_yZ}{aV)�QS��%L:l��}� <G�*�P�Ua���S�'��(o�uu��f�i�V�� �mo5�b��f/��Z�ރ�p��Vwk�1�?����az��08�E����g
v�*�ܤt�L�V2�¨�pǴ�d?-����-�F<� o�j ���V�6g��mP�x7�J����V�Ek��d��hN��*�8��
��^8~���@H�s��ש�b��9>z@�CL5�^����W�~!���^��7`Πl)s�#�Dl�7��P�&TC�5������Ik���\�4��|Z��{%�zϹI�4U�/W������}(��p�__����rfW^}��k����m��*M�ӻ�����ף���a��E豞��D����q#8�h��Z�ء�Be"h���N4|H2���<��n�Ѣ�uW���0���GS�
��yA�`Cs3�!��X�h@Y����ў84�=����P
9���ʃ!�%�ҺF1��$z<����LT���b1�Ai�ww��)L^;���-�}RQ��6��gU�c�i�;����'A��v|�����a���^=Cg��i_C(�@�%xp�7�S�D����З�W<�N�R+)֬J�q2t�S|-9 �m�r54��RS���a�m�	�*�/ � ��:9s���&?m`��W��5z)�{�`���۾�U��;*�L�~��u�?�U�D�{���F�;���
��@�b���Ǒ�)�)�.��?�ԓc����U�c Y�@Y�!~�4Im� ĵJRD�u�;g� Z����e�~W�1�b��e4�y��P��F!_�g��]y��B��	�}�A��:��UV={s:�&�i5;����Ƿ�՚��3��KGpl�kT.fD�^I��s�4O�~�TMjݲ�T֩�fU{{�Cy��s���#��H��m���e�#a���Y�B�)gK,�
}�3�-i:s��?�Z�)���$]���T����0�It-�`gKY�G�y�'���o�8�WU����u��	���,{����}�R�
��+8����祖`��fbD�&Qj^'�0��O�$��V�wr�t�γ�>��<|���ҵ����&S� ��bBcT������P��c��Ϩƛ����yف쁰��g��S�����~�N3+�"c�U`e��X�T��ZP����!i+���F��3�����i<~�ú�f���
��f�������w�=�g̇/����9�����.�)��
F/j&CS	 ̀���*3e�����әF	F����'�4C}��e�-+q[�%ko���~T Q�d#����|�@g*� -m0����&�&L���'\hGƍ+>�6D�_��Rי���W��rnm�O�i��v�q`��}�.�f���#��/m�x��p$ɫOǛn6�ě��o��sRvk+�=���gUQA4�^����9��ʶ�^i�^�ɗ-�\�h$(������-�`��"����~���L�.�!f~�Z�"v}}X?(�<�Q_O��)�\���ݲy&,�Cb��gߵ���vwݗ��S�����wl�;q?P�;+��((ʘW�B��x8�Qg��*���y�s�� ��3#���#���g��T+��9��Ļ� a+�w�!_�B�đ������]2�W�[�)ٱ��3~�w�V���s.np[dX��9���s��k�ЛdT�/�i�t�垱�2�����b[�)�I���y�aO�]��'o�w���ν�3�U�P'
k���1>�T��I��$�kt7�5qD�9T_��"{���S��)�OΝ�;�(����Q�$����zr�i?sG�!����k�1&�#Bb��t2���n�NF�笖qs]~3d0���Ob�XFB��s)�?��0]�V�w���2��b�Xv\�z��fl_�vyxB�����uF�d-���e�߃��~F�R>ۑ8��-}>^��x�� a�3�K!>�n���l��>�?�������uwy-䑢�T7���5�-�����x㧲�Ũ�a>���l��QC��R]Ԏks��bSS|�%�;� ~�`5Q��ڀ8MF���+ȟ(���k�J�q�_���P7�ӫ8�@�*R}���Q��aɝ��!��]�,i6O>�*Vp�V��3�x�i����^Μ围�.�P��	Q^�o!V�=����yJ[�pL��_�<���\�:�Uq��0��t[7@6�!��ӧ^a���8���\��d�i���J��E3��x3��R@��fwѴ%x���e�MĢ�ZDD��IxaB�G_Yڤ� :}�e�:����k{�x��g%x����>
Y�����+Q�;��|�����';���)��=r�'����`����y
��E�/�Ҹ˩J�2%�vIUe�l��ݙ�ՙu�7,F��p���,z.�	@&�
]>�C���Y�>_��_�����j�9�TDB2�7X��܊�[<�Ә~�����6~�A�bﺇ�jW>�B��wY��f��ήoU�E>��~$O�.����������Vm� �ꥼT�Y������`�O�3=��?u�9Ҍ�q��3�#�W����B�q,'x��#�Z�	��r+0���ɣY��nzR&X�"/޻�J�?s���%'To��yI��GOG�4�e��5�>U�I�8-/��L�d[4G���|��S�8A�Cl4��2��?8[��z�.�dk<��\q�{+D|�Q��F3�v��ؾy|9�z�\"d�n=穦��}y���/=�w�VM~�bQ`=^ �g� x�[!&9���]d����x�1�k;���Ǚ�fԥ�h{o|�����Y�Jc�/�9[Ѳn��O�k?��x��������V�&ݖp���-�+��3���8q�{*�3;�$�M�,��-��BH�P	/�Ԩ�����+�@����Z���H�s�y�b���t����kް��#��=�.�)�.��s���Jq"�o���z}*J�����ɴ�r�����g��DL�կ���<
v1��G���(4�J�7~�6�Uᱫm�DV�=�AoN���Y�	��ҳ��s��ci��+g�6�����Ta�t�xU��e���T��S@�֓�a��8AhN{����d|�sᆎ�.C{U5����E�
�w��,	���wl(ޭ�N�۾#����	NhҡT�c�����S���/īd���'K�<ݕbA#0̶�Iȁ�<w��A���6����. �'x����}*��?ӕ8�����b.���
�Vwv�2sH|vɼد�y{�pp��c_�_�L��i���qY������-������lޤ�L���7�0鉳	� ~�дl�f�y���v��A���-k�B3h�7T'�}�+���9�^���gH,7n0+��O.�����u��(5/�� ~�g�#���3onz�p�}����;U�^/��:mHO9��� c߰J�A�"1:p�Mɷ��c����7�����k�������q-
_!��L�&&�,e,����� <8��KjCݕ���t����h\���4/��k�R۪��v��(�����ȗ�ڴ;0��V��b��!�\b�^�}y�m�W�oQ�B~����C����r����st��*7����6, \R���)��c6#�ރhʢCC�����GǴ�csE�=f�g�k��x���z��+ռٝ\:�������3$���a���P�k�)txZw�g]?2	��3m���>(�=�K��VtZ?Na��Ȳ�(�\�,��{V��) ��?g�9˦L�b��w[T~���*KI��;����/&�� ��5���=֯0yI�G�rENG@e0���Z,�`������	�ힵ�*��Z� ���8{���I���ٸ�myNm�HCo�^&��ħ�S>|��V�X�]�WQ��*��Sz�/je���U3XG]���6��3ξ�zh����X�):���egN�݂�`�*P6K'뼼]�ojj�G���5�*ϰ�G����i-��ʧ�w��ۂP�}���K�To�0Y�*���<��1s����(�'�Ε���j�r����x�y{��|�P�{�)���W��?��U���c������ک��'s��O�_�p���-挙Q�����8�Ib��J��)�e�߭���!�WS��$����*����0m2�N��o�`7l�`����⸘�������Ni�������+1J��vk*��̼�͏V�K��m�������b����L��u�Y�* ���h�X;_9�l&,��U���%��Ηm`,����ո�y�!�9�p�O�̬��J.`����sX	f��7P�F%e���՞��?n�*���ˍH��/e��a{�W70�4���y"j��c�j�*�������&S��*��l�NOg���~�����@L�Z���>cMU~�{�~a�2d~8�
Ux�n>O>I�<����<�:V=;�s��N� �M��6��ױ.�uF<H��n��ǯ�;?|���T�P!�[��g�nh������n�����[�sc"������;*W���w��/њ�ꦒ$XSb0��7W�,A�Rh�jr�>�f(PssH�#<�n�s�M�ۆ%F���P�p�^[*p.��Y�f�|�Yǲ7���w#�H�e�CaŪg(�A��X޼���r���n,�n����7փ?3 �R{�t]�.*�kY�Q^��o~+�5���O=��2o����x+;���}�j����bb�s��\�lw"g��{�y�h�=o`��I˫ę+��N�rܽ�$qp�D���+`o�Ϥ,T��_K,�Q[��&�Zhk��L����,$YC����q�}>�j
i4���ܝ����duT�he�T��rM_5���XG��U�k�-2��W� ���)�fę�j������� ��
Y��<�������@��4����9�֗��W�_��K�>u8�'�3������K ���ف����9�r@��9X&ӴT�Z¹F1-�r��*#{�t���~��>�7�^�]X��}�^�ft��v�
�� Qܹ)��5���p&T���uY�9oE��a�Z@VB��"U.�)Ǒv���ږ2��!+-�^DS"dvIӌ�O�� �ӛ��xš\�z���Tl+[���\)��S�|<X��&M���1P��C�W�oH|�Kq�?�˨S�T�gWL�Iv���K��~���!��#`�#9��ڣ��U���W�ߞ@}�
 �'�95�/RT1-�T?ɠ�PLo��r�$�ݮ����x��K��o��A�
r���/v�&[�]{��ej��"3��8����x�Zo�ᔹ�ݝ����wǷ*u�7�I��F%��@�2z��dؑ4c��͊C\ ���E��6FG�M�y��R/u�o6��pה	�w�,�����<�@R91\5����ũa�җ�T�}pwTrBP��1�0	K�N���=y�!>����X_�a���������_���D�7�ݮp�P[�*C�@I�?/�Hx̲\[�E�$N���#O��_|���}���=�R��y�xU�Pj��Kl��ȷ�nc|�]kpl�:u�y$xu�X�mw!�S@�qj�n�,�ې бa�z��׮�%��3�����a�/׍>D�������+�o�<;z��ߜ���Q�L�/Qj�8'���D�K�kpT�� .�Q;���䘦��ò������)��C	_�(��ٸT��:��`���D҂E��_���гT�2�MI���B�m{T
M_|׺�������\|X�K�J�����Kfu�ҍ�3X��]�ft�@�����w�ߟ2��u~��*�
,.p�qM��愾&!`�F�� ܢ���t@>�s��/D�{�Fv�E�v��n�8!�tͪX�!!��&M^����L�8W<�pI�#��bi6��
Qh�B-�X�k2T��3�'�Q����$8F]y(�ۀ�1H1ͭ3���o�!�:�%X���Μ�+F�O.��*g����Oe����0�T��0�xM- A�5hk$��� ~�Q/>��e�2*�k ��[��(�����03TW��m��4�C���Q
]PNN}gO�$��q%�(�!B�X�$\n�y^���`�m!��	�Cy��?5N@Xn��$�� p�
�k��7O�I7�*fz|f`�?!h�}�p��N���J�(e�qTڳ�J���Y��DH��@�(K�����^1>20d����R��*�̱j' �rJw�c�X���!��\�<���Y��h^΄tm�0�[5�
�楗��ۃ�EoD�����֮�hcL\bv��殤���2�Ju���Y=��y ;�p��Nr�jMu��>u�g�Ie~��4�T��#�S�L�3G��os��)���:�}ew``f�u3@���kbU���-�(�m����v:�s�;'�
�K�p��v-��.^�G�݊����Fc��S��������(���yL'��oGX[Z�W�|t�B���ռ$2��5<�GW�S';����϶ū���'f�Z���J�ιI9_�,���fP��GH�s��9U��t����e� Zd�$VT,]����j�t��*�J�5�w�QE rԑ�k]��BX�K�vf����[%�W�9[?%|�>�B��!��q"���.g0B�qJ&98�s2]L=�O��(�i���=q�~W0��������6�����'vǻ����cz% �RZ�k�;��M�FU�P:�8V_�nj,o��w!&(����6�l�����IFˍ�8g�&S�u����ƴ$au]�E`���%��o�p�GU���H�m5�lz<�B���@�uJW5�i�┎_�Tbl�����]@r���Ϭ�����F?���׆Yo����N59Y��\��w�[��(�2O�Tx�_ơ̈̄��$&�ь&���ONZ�O�/mpC�:)�Y�Y�=&�ה�OҌ��:��ڍ]|h�1��)=E��ӳ�俇uf@��*�H�
0���(���D�A���I��cɬ�P�䊮W �	q�,OxVH����;��o�o�7it�y;ߙ1���mZܷ�D;�0��"%ǫ�U�&,�W� Bм��6*�3k�6������2�	�ɒ����٪�C��+���$�(�<:�oAm��I��8~#vG?=Fu<tzK�yP؟����Z�&҆F�RsX�ICf:��MOj�����Go�.�y�Mq�4D�x ���d�$<�vrGT6��X�:01UbY�=L��Dx�tCf�1��xĲ.ˌ�Vl=�`Um����?rw��(��vE��d�Lk�J1�A��pcbi�;�lّ����W�؁7��7��e�������7�~�k�_�t�����Oy��%��"���}Ph�k��T������F>;��M����נ^0"ȟ2�`ŗN�syW�&ho%hL�L�-�U��HUa>>n�D�LT6x�E�k�ߔ��3~�U~1C�`�� `�����;��j~yHl;L)�5R��o��"���˵��!!-G��{,,��y��颫�0N�j��sܾ�s���5�V������"�~����ԙ�,�Q(��J�$��G�ޕ5�h�驜�)r�1r�ؔ�pu�-���l�)G���䭺[Mv�1J[j�`t~r��#3�C:��w�g�>�۟��Lb�O�=��R#���`.��Ӯ�tN�EB�
'KV1F��5~��I$��z'�^��Y��	�x�"��y��"o%��Nn���#"����A�?fQ��c��eg�>���iV���?����.?�2�����TFV�-�T4�J-��	<���^i#	}�Q���_ڑCN������Xtj&�l\ƫsR�8Hn���_�l�罐�O�ήdψ�_��S5_���[�h��Z�ƹ��D�ц���zi����$��0q��'�W���P\�(�JE��N�������>���D��Bi!F^�>�h�/F�V&e�63C{f���ҁc��C�Y����?z���<LE�V}�����ap`���VŋtT����"]�#�U,��SGM�$r#J��KwM���4Ę���%Z�a^V1,���������K���bM�lq�OX�v�����_�↷�2��	����ρ1aؘ������'��9j�o_q�o�h�>ۑ��_�G�t����w$��ͧj��9����yf���6k-�h2��L�`��E�·nppK�kze�VyN�0�����	DrּE'�,Y��s����=V�n#wd�tH��ו��(���Ω}��S~����_���̴�@�"�[��+�}�R�D )��y@�u��؅\�*�WP��Z����߯l���wJ�lG��&4$[�!X��XR�"E�������L��H-��u����,��-���߃@�0&�9T؎8��������A���!Ln�Bd�0}�S/�4�8�N�&�AaX�P7Ű��U=�"�o���5��Y?��7�!;�Hi9�g��i�t�9/���:�0�Y�N�%��dy��rnlu�Bs��o����~�CXq��(�"��@�q��#j4t4��'��چ7�&$��ՈU:"�\&w���}���С܆�=N$l䜣�px�d�)�L]����W���F����ފ��P�D��������O�	���U��@"�>O�J�zL���v�KP�へ�� "�����}Y~f����g��U���G')���g�N]���E�M�\�"͵��c�G�CZk�"�_�B-��IJ�Z�0���G�<�"P���?��8Fi>z�K^�b�ˎ�����$(�2#��v�qlkt��_sy;V�-��Ɯ, �Ǌ�,���?�Uَ֋��w��;�,�Q����7�uQ�	�������iM���˓m;Q]؉S��*�ˣ��~������h%���"ʳ��5�C�V�Lv>�{.�P�#����I�0�[;:��Y�w�H�b�ch�ZeN�\�D&��Ip�ì ��4qh��I�G40�_�D�'*G�d��r��K ��S�]�T����d�� ������Y"���5�.>Vr�م��u���pN��j>2�"��ʷ8����-ذ�V�1���Bw��(�rN��Ok����d�[��� ��f�gSr۰Bw�Wo=Lg�
1���X�eP� a�=���a����!{����K��Hq��@P�-�c�YI�0�R���/�N��dG��HՊ�kcs�C���j!�V��H�-�v�?�?�5���e��8��e9���k�������AE&���1���74 6>�q4��8P�5��Ϡ#\�b��Zz-~v�#��� ��Ԫ�x�w0+V�O��u��@b����:��^���f���H�AUԈ�n�����R�[���v�]m!	<|?i�ew���$���SG�i��n���:�s6-%F�Y����.���
��/�`�	�8l����*����>�g��l2IasB�p����9iƿ=���������)K�E�-��f����.��_�XgB�LeZ00�^�����n�cf�48Xr)���E���}ݚ�\��?L}u\T��5��� � �%RCIKw7J7�RR��#0 C7����tI�t�Π������9�9;�^k�=�L�Y�¿����V^V�����T�&�'�*�-��g�j�}G��0tr�_4�����?�gM� ��7�9�ρt�صڮ��w�>*;��I�p��Ac0�E�p��7��ɐ��i����o`��E #�ƥ+삾�u b+o�2�v�����i�(}��z!�`���n�V�))����A�cl��1b�!���;��[kVЁ@��
\_�t�s*��,� Xo�T�6�X���9o�U]�gt����[j�����l۩��F���h��^�b��x�����HӴ8���H�(,�f���(� 8�1q�UBO-�S�O9�g;��F�a+��-�4�VTy��b.A���{��j����Y �b����������U�	�0Ɓ�n�e��s�8��)��C�U�l~�SQf�XuWU���r]�����F�TO#aU����Uۿ%NӞ�5&b@e�����y�۲M�L5����yY��7�������6�z�7l��	�n��ۮ���q	�)�I="S�7�C�Z����˸C���K��bi���۱ܥp ٺ��Q�Ք�~�ϽA�����2���L�B��]WǛ�ؾ�955����|�_�HO��8���/ɱA2B�z�ed�c���m�[j9Q�X�ۀ(A��w� "�S�ۜ�5m��A�y�T�G;�L�M��8~Y|Xn2h5՟���߫�8�nr�2�V~F�� tt7yt��讎�y�sc�>0!sa��f8�G���[͂A{�!�N��v͢��Ϣ_͈3��'@��a�`м�SR��/�[���=� #x�h��}�``��Q����<^��H��C��
C�*ejDE�Js����0�-��Kv�����^̃T���K��Ş�Aw�]�]�hR��]�R;C�v��c�赳�����V)�)-5��:v����e�r ���-@U���@z,�ic<��p|�ʿx7��utX���(�S���Ӥ��L�������&̍�(u��"�c�&13������J��˫E�˫��ur �O��������L��PR-��Qx>�N�����ڃǙ��;�ʙ�p�ʕ��l�Sy4Tqq���UV	(6U��+G�j����%L�+��K����m�x�,���)p�*�qw�;	��v+D(�i�/�H$o���a�£����[�����!ȭO#J�gNG;R�:�G���Mu70��}�0��� A����y��=��6n�|�0/fTIv�qtt]H��<?{����;J��k��qh�ڣp<��k�s;���j��i8�R�Vc�TۥD�l2�9�R�yؚ����B�:~d&}�K@���$P����d��?�D�m`��)�SRkJ��(��K�G.r+B&��U��vKkkϬ1�}2�S�l���؄qr�A8]�U�MX��6�3r��^TC#�K�@�;�!w��JF�զR�N�7�_��摜h�e��2���b�
!yw~|��!;��s��F��N9�O����!j
,)A�3�L  �DDŖ)7�M���#"�ꛍ]}$��6ͳ����3$��zSTa>���1e]� ��ɳ�����E�"��9�� \%ȱ#���|���.O�k~ވ͗��3O�H޾�2���р���d� dn;��q ���R!�;�sjW�`�X!��cm�"eo$9�O��Q�{�[4����ԣk����� o������#���G�d�~���~;
&C��Y<�!�����&�m"���&�@b�k��X�����	��A��^0����g+���]�7^̙C�o���P���)�n����[
���V�s����f��:��{1�����~�l��:%N����f�F���FڣYM�!�{g(����hg1DT�'1]��'�c0	ᦖ5a崻��gD����i����d'niU�5��Z�(�o�!�X�|ac�7rJq�������w>E"��g�,��Z\/tb6i��� r�k�H�Nn���B�{��X�&)1Ͽ�0 ןN콩�oT�����>����q�0�d����hO��fxM"
Gb��$�����ʲ�>ql��_�8����%���sF^�d�߂ET�?:~]1��:�k��.������z�٨��c�Sr*4����L�-ݨ0Hw5P|��VY�
&B�bv!$���6�(���٦��?�J���XU۽ڞ�/�Vh�E����ǪGA^�2&�$3������R�""5���p�ւ[�M�����3�X�i���s�" �a'�G���a,.�!g��u�<�b�9�^�U5�kLa�<@�`+�n(�)�*�!���?�;9������p����p��	m2�1D1@j��`���F�	I�n���<��/�y�H{�U�6:���FD�x��6Kl�n�?��Zi�z=��t_�\��!x���~1"��>�,|*�x4�68	��� ��� �3�J� x��^|���g=շ�d������g�͂�@�f��N�� ��X|��\���" ����;�Ly��}����-zl<5,�pH���f=v��Pm�_�wuf���$��S�7pD4��"{K���I��.YV-�s|��߱#�iW�#��Y$��~��>�{��I*b+��AѲZ6���2�]�f�[��X�;�y7l��x1ŧ�\�������	ȕ[��O'f��y28SE_�ˌ?xBDr�y�m'�K�=��oe�i�|eJPZ��9>��B���T���O}�����X�&E��(�M����J#�wG�AL����]��!�g �y~_��[}�oa���x�6so2@<2_@�� 	r�=��~|"b~�����ҩ̌N��k:@�!��kf��f�i���t}�Q�A�(���h����u�b!�o_.�5Tm�X��\�Q!~Ws=�g�v�fGզ���̢�6���Nfs�� �I0���̻�4��?O��XRG��2O��gU�u�QRYћ�-�ן5*����efv��c���:x��p�i�1#�i]���g���N�����jJ|��:W��e�M��9~U�ED���dHvm�I��+�X�E�J 
5��3
f��J4�����^	�J�-��%��� z���k�~��:�eo�9z@)`����������U�������b��%�*ULgV�F���B�g�@m��(f��@����~���a �i+���~�{%��c�O�`��){�����A�L��G�خ6aΊ�������z�Ӗ*��G�H�� �8���7���4�8ſ3�>�0�%��j�]�8�N�[rȮD�G�1����\��S�{�V�+s�L��TwŨ0 �3*;/,~q� �d�p�3�s�������:~�b�mAf������[	�Z!"�J^�(�Z�4���C��abz��?��*Z+*��C���LV��X<*�AL] �H������H��Ub�.�wBhj0k�̏���N�heC_�q��n-��F�;�N��e���c��ƗKz��Kq�`����o�eQh�ӡ!�[������l�l��
�c�����<���6�^��I��l�1��u>Cm\ֈ����~�(%$��5q)� �+[#f{J65�h���Ds�|�וV���B�b��@�P?�Z�_~�_ ݗH��l\��!�/#O��˝�5���s�ۍ�Z�ˁ��l��#ݾ��E&q�.�U�����2D:��ԗ4�EN,�Ê��	��� �u��P8�j!�Q8�Q��) ��4E,O��NQ��n��[Ъ�!R� �|*��^q������ز θ�ԅX���(���s���'Dl���I�2�"�Q��e:zy��>.V�l~��s]ca㒳v{��٠]�$�=ڂ�̙:�%T���l�0����^��wH/]�\he�5��\Ij�����y�����d����m?1���.Z�^6Vz#U,��S��ߨ��5t�|3������myq�ZZ$\f̑��qf���K��r+ͦ����Ѽ	_2���}�����۝�,5G�2.�/AtqwF�t�R�\k�QY�����EHPI;D���IS�Y��u{w���}D�eCkN�])kyTz�[s"�E�J[J��&��j�_���E���i�+@T��;����0_�d*s�E�f�)>nr+��v=*����A
�VtK[T��v���pe7�}k$�.C}ʜe ��( ��/)��0{9����� 0^�d�z��&�>{�"#>�я8�=Pm|-��+f�t��M�ל*�Ǌ��N�'�=���&�V�0l�A����en0`pZ (o�r�K���������?ij��XPN-V�J-
0�4ٿG�v	�q���SQX�P��.��J�.HPpų0vpP����(4�/L�h����vu��.2N5p�uv����]�q�o�@ *1*~}����X�ru�n��ѭ<C��@Aa�o� Qw^�������/���[�Y��G_��X�[�[7�y��(��NS|OϺ辴�"$\�B�&�`5�m��/7w=\�4r��1��X.��?E�*��5�k�?zq
1B0����ӱ3���{~�邙?# P�!Z��J�x9)�$�������G�e�:����j+#Q�j<8����W��6����\K������CC��Q "�Sİۑ��B|�Ύ(�[��C�e�F^,\g,G}�B
���^.��-�9-������G��	ng�Z<u��ܭ�F�y�������� l |��܏��yGf�f;q��G�ctL$?$��%�������Q�^�%��Z�U�r �|�$8xL8����ƨ�S���ye�����(F�wJ�)Y]bP�C��0�(:�e�b�h����'�:�
��|�O��_G�FI_�֕�W�� 8��T��ۜ���}ۄx�s��͜���M�`v�;���E@y;W�ځ-Kb9�Ap�o(b�����aOL�y������3����_{�[���Ց E]���$��d<M4:/��"mj8b��|�l^�w2����j���մS�s#���pv�[0j���ń�}	����k�%���Ʃ����<u�i�?~�t(�� ;���| Cl���RRf��(c%�V�|ķ[�53���k�N� ��q�e/k�$6��N�d��s:d�]a2v Y���8_�8O���GO]X?�� �Oޟ���.0������~RCnnB��׭�Ɂl+������h��T��;R�xŏ�b펠H���;�&��,�eK�m��g�3�Lj�Kh Q�h;R3N�	��E�8|��El�IP�jh�'@��������9>b�<D�KbW;��Ky b��;��U�9�w���(����y�&o5W���<��e0_�,F�-�
������{�`�3=(D{�����:1�6��NP��\��r�����3pX{�T��u�o��g�+��I'&��ۜ�qZ���;��MV��Ԣ�Mx��uT�N�VSN���ԨB��.sV���\#�S�I�ҠhK��1,�B�Bg��V�Se��!u�Ľ��}v��u5Fl�gui#qA[��Cg����DNԔ������c�����oo��>}�՛۪�3�p��0����-z�J<`-�"�ݠ�ܿ���1��O�2�AO��t
Ũ���?"��acX�����u�׬�=ۧq��keh|���p���M�_�2	=AL,�q�b��2�Q̯X猶\;�u�jݿN��W92�^���@}T�%�K���6����&+=@1h��5�)\�Ӓ|CK����U%�ٶ���6�y�&���o�ϕlҲl+k�������߾���$A�j����t�Uu�J��LܮnK���'vDH�7<�	�Z� )Y�y!����O���F����e�ZQ:b}�/_�ZZ�_��Ȟ�SPZ{HH�j/�e�3��B�" ������gU]x���wջ���.��?�1�%�!��� V�E���W̦�~I�L$=H'��}�c�'�^��e/�ܙ���k�(��*��'��V��}�bBA�C�=G���o	G3]�V.���+�f�Uژ��8^UĊ"�����@�o�(�g
p������u��ZG�t٥���c?uA,�f��hgǙ�[P�?)������������=4������oFx��\�4ʂ�{oc Rc��.�;ڑZ���Z� �0[�4���X*֥���5;�;~�"�j��g�l�9�^R�4 �����q��3�v���s�Ζ��^�d:�'�Q���A-���)�Y5�j��s�/���I ��׎���4�`��gg\��X�xe��1'����A!-7�;��T[������?oz��@�.hg��[�����Ji@ɗ��x��D�
��p^��zʌ����ᥚ4K����4���럏���Z��Qѕ�(}3�\'�z����#o�Ot�U���� m�~2��#>d�b��$�L���+�-�F�~y�s�B���B�����3��҂Rlu�ޥ��'��>�5�	m�\�7
/
 7wՓa�E��_�R��ߗo�(<i�bU�ܡ�m�T�I���uNۓ&�Ŋ��l��o1�Շ}.�Pp~'�H���zz����b܂�(�zf
&h�K�j�!Ӣ�E�,3H��a�J�� �����5��g8���2C�=���&r�j�$J����̑.[��v�.�7222DGKO��5��{���DBTC�5���q�2{�h;Vi&�я�8ͱ4�~�*4��7\�n���f�@��Ց�ݿ���+��a9N�bu��WVW
����o��A�O��:B�a*���޽�aX��	]��UfK+��fS�2�:��Yq��'��"��O>@��~�p��<���R�*�/QZZb7<�k���-#�Ό��䖘�1��gAuufPT��F5���Fɶ�����V�[�����Q�j�n�׹�\�'ԝ��)��8�57��x��|c{�"�=�����kr_;��\1���PNB&�����:�t�w�Ȝ�	�UAJ��8b��=[��C������� vU�r2�ܿ;���D��P�3���<��*HE;ǎ�%&�f�c�h�w�X~���O&��-����c��v�jn� �l`�>xj'�+I��/�S�1��X��
�?�5F���}���U����c)|o�_�(�A����ZS>w�(o9�۠�]z���B���%@�Y�澠Nir��+�jF�}�G�1�R�鴂~�?��?�����4��#��嵰#��=���2���>���:�nHj�Sp�g?e��Ja��28,]E#_���y���tz|D���Y��/朊=��t���tR�4g����2��m����/w�W�R�>1v*h�h��&�k�����g�����^S��)P�f�ZHhsc,��ʖ͘�������	���F	���l'�66��eW �0A�ЗFZp�wb�T�����5��4�?\�-#��.���Ym���C��j���J�4������pZPT����0'�3~0�M�(�O�u��J>>Dr,�؀�]��[ �,�h G=���U��~��\G�E��^�\r�$N���T���C,�+�W�a޺��Ei1�W�K�&��g�Ǿ���#k_����k���+���Yvqѷ��Í�!�\w7�+��-�-h}��^���Ev8}�Ǻ�pfTѸt�x&�|�N��!���U��\x�cm��	>��垭�f�C�T'&.1�Rx4`8�3,�!QP(�Zf�"#Ɇ�[Zb�O `���g-���~���w�~S�A}�u���<�z#,��/ �����x�j�1�C����h�ܒL<��$�s�ݠoq�Z��e��~z�����xT���/�R7�da/e�g�5�\���$��1��o��V�;�E'�j�2̅IC���b��'�H�ZJ���
qt'���ͯ0D��^>��>c�M�n�����~.�%�9��\��B���Tm�U�h�t|����7y�h�Q\([*�ėg���&j�)g=��^���#j�Չ|�ڎ�EK��HB�4��;�{�Ebh�lyRj������ڛ����?,�*�\�AT�T4 Vnَ/Q�]��5R�#������o?{���0��jD>�����R��2��0��	��I�`���DKF9��1�D�N���k��$Ό�s6�oB߶�hW���2��((�*��$��mN�>��x��!j�W��YS��M�S�-ٲUdXy_��O��5ϦB�SFD�__�f�!ɫ~��,r�.�V�@����`;��(�8����({ N�nO��_�
<;�}�%\�gQ�}��J��?kډ"V���3L�(���PQ{�Q�P� ��K�:������bR3'a&���ߓ@���Tί��Zj��G�Tڃ������v��n}��k�?>s(��r�s��# ���@z��MH�I�d�Dꔌ̧;;k��u�7����d�����R6�j��}�U�O�׶[���{ETړ�^f�i�ث���>C���R}�M�^�g��!(T�*��{���^��������*Z��
���?�ۅx��i���|��+�۠b��$�9-�I�6 �7u��&z�m���e ���8��h����=O ��)cg��x`��.CB�2ڿPOm���?ў5����9�vrNo��W�-�^kr�>�����ؖ��-ݖ9{j̬����k��~X�3�nm&X����.__�O�7���+C�͛�5��<�.? ^�O�\e�O\<��%�:�߳�+�V�W�/|��%�9{�T]�IOO�ʜ��^�Wu�{�E��{�O�s�}���{?�@�E���s�ߨ'P�z��)"+��cBa1j� ���[7�JJ��H
~��yn��?�aD�B�~�%S�6��8�N~�?��ډ����r~��UO0[8$�g�G5\Ե�`s!�]%ך���.�H��κ3�HH]�^,2�n�ZU�AW\q@[�_Iۏy@��4w:�~^Svs\�L�.�-a���U-�8��wR�����1����ԚO����u����l�@�K��u��� �j�Y��쫁�NM8�ܳ:��u�ˈVA��l���s5����l�c?�т@��R+\�aȽ���)R`����A�`r?S����y��bą�ͦ,��ҫ�1�+r���ʔm��.+�� ��U�u�SG��p�J8��!Iv�����	s�g�O�u�cS��ol����*���@_�U�ۉ���e:�|��Ǆ􄷨�h������I�1���Ns�N�I�6E^U�Li�$�)X�9v)��Ȳ�oŌ��>����D��O<�[p�*/Zu��`?�%DN$���-�oLWq �)_cͩ����� x~��3oP���P����}��IZq�֥���h�����~qY�E��o�f'F5�o�v5y�979rlKv���]6i�`�b0�y��`��u�D�$�d.R5?̞�v�,���������n��'�c��AC�h��p��]M�pޞ`�5���̶�e���w�K���Ť����A�k}��@���E��N��c�ƭ�?�Ďl� ��A�0TJ��'�s/&�����C�jPv��'��Att6l���L˗���Z�И�qn��o���a�N�<h7.5UlƕI�.�Y\0���`��G��U�K/��9����K*�:�%.��R��-�[YoI�8>�Y�qǚ�?��;S\��us|��7'�oM���7
�\䁽NYo�찗E��^~�����w��MmS�R�,**%�v���c�hg�q���z����pW�;������2uУIQCrѣ�2q�2:T�?�]��v�Wdi˵�e&n�po�Uy�2�[0���uu���&�H���Z���ڷ�KÞ�ӡ���e�ٰ����I�kk�/���z��i��hk�49`�����A�����'��<�w�aw�;��t=�g�n6�+��,����G��[����u��l��d���ҧ�d6��!��������3꼍��>?��Ɣ@�j�NyN��r�I�p�Z�uK�)5^���>�:N*}f�ޔ+��jԠЧ���+�p������?�$��1J���l�aP�	����P�ד�a46j�&��� �1<s�REBx����Qt��D*�v�	�_���� *����rN�"�����t�����L��:��i܅����LwL�6���c�.�R'sZ�~�v�}�a�	��ޛ��+���d~�ȓ²������}$�v��V�%	��>OH�cf�|���o�@Y�?�9�{�i��6b��I��K�bw!�Â�Tz���86Q��Ds,�l�0�#����j3ԭ��p��'.MNE~�}ݝzu��O7M@��|�� �}T�M�.��Jt!���`�;,�!ț�O_�@��T<0�R/�P�/*���qϒd��~�c���?#J�6:���{p'_����m���tw0x+Ȟ��H�H��GvTC�t)pG��Y��c=�PN����EX΃_n3tU��q�B�JC���.��=�����eD�9�Gɔ>��T�F�D9L���|�ȡ���6.8�.L���,'��+�0?Л�m��"�G�폺�2��#�MDI�:N�f���i��oz'�|�B� �K�;y����F}2�Oo��}��X�X 0UCK$�����P�7��<��/>����G@�$5�7b����Ɖ�5�)�A�#O>O
74��y��E�M>Qw&��\��㬢�&g	����&O©h-���Ȼ[3��3�xF��	���d�S�͖���$�o�c��\6o$�LlX���^��&o1��?B�2��Zj*J��J�]�F�]h�j�����ש�I���u7��Dco�+�٫�Bo��Qw"�,X��R����æ�,K�h@@��-_cV"u�l�~?�s&�
����F��}��N$6_��c���E��ʍz��5E0�����ّQ���1j��-�&̭�G"�U��$�+#��w{J�?}=��o'�k{�c�+h��H���wV�C	��)�� �5'C����󳾸�&����kv��"K���/y4xΰF�C.F�G8���~����s.o�t�Q����<� ���x�)�f��6�@� ���QE�>h��@� t�����_z��I�L s�1�鸓��5IK�Mt�T�Q���� ocFz���]�i��䑶A �� D.�Y'C wQ�sg�\�J=3�T�$Wwe�t�"�7t���oڐ[A\����&K���++<#�Хs2)�r"h|ݡ�O��C����~[����ꮄR�A�p�PZ�P�\�'�r�:2�zw��<N����9P�S�֌�[ܿ_���D9}S�O�Ҏ+�[�X�6@���� �Y���WC�s�+�\�{':�W�N�e����2~�.��qz ZC6�A"�]�k��!���v$�5�7X��9� ;Ocg.ܲ��9��VC �}gp��B��{��ΐ��Z� |�=��oW}����?�V�拏u�e�W���� �p��bZK��hg�uR@����f��4���-�C���;Yb�~zE?!�R|������>!�0�-?(N���01������.�=��V��ƺ�R�<�E�偺�xx�T���#mm  )�Š���PE{���6�^��~�0��
������N����d�3���D�[X�!B�< ��߻9pՔe��X��N�M��������'�tW������[η(�)���=�|7�`j(�i4�-���cX�����.;	���O�ӫe���8�-%b7�͞_�$�vt�ּH_��5���Q]�����?�FP���9�e�m>%����Q�����h��1 �!x+�s"�����ط�?#i���L��r0��
~����H�s'�R���I]�g�N�5e��D�k��$ $/���Uw��M _5Ϙx�N�M�����\�fMK1GH���l�Y�����S���p����e_0c�����Z2RM�FR��򲃃���^ W9�u��/��n�8,R�q�q
s���E�Y;���oJ�:�t�a,��9���PL�Cm��5_Y�1�lx�u�r尽��1�)��6s#���'J�A�iU��u_���ꂍ|�����nyŦ��C�4 �ݿ���,���rQ������������#m6�G�F}I^}x�.8c�����*e��-�T �TM��si+P�!Xx:�	cn.�:L�ﮍ�'w��J7��+���c��v����%@"];�A��Y(ڭ��_q1U��l�(�NB��6��^cX�=dp6���L�N"��E�7U�4��*.��<i__�x�x����t2�~�"A���]�6�,�ל
"�������4d����]�0F~`d`�
�Y��Oİ�X4�_�W��M~�;;�}�o��-_�\�P^o����a�YșN��٘�����$E�&��S�7K��`J�W�=��}��O������$g��i^/OH�z {��A��ĵ�ʟ�?;jrM� wɕ��]OR@��t�4�Nl���֡���� �4��l�� &��QQ#z�W�6ܢm��h�?
�+�?��
4�B@&���N4~d��"�����r�r�MF��5G�X�'��M�[�h8	Sd� ��|��y2��`������4]g~C�;l'u�Lb��/vT�����'3�Úx���J�hF��J�U� 2q�S�3�<���L`�gHR�w�A��,>�:܎�.�t�������Z
����IO�H�]�g��F�j|q Ѵ&����@�����ߙ 'F��6`J͜ ��4��� �Q�H�1P�\rԠ;kb�;_Y��y�W��F�o?�h츜��T���Y�����ˣ@��f�<�5���11��Ps��`�΀��"�,!?�g)}2���X[���xpX�1�AL[�R��=��?@kQ��m�)�O��̶��O>F�'���k.a��ֿV�4��B���yJ�v���W��SF�"���K��*&n��P~�K$��]_2Nl���f�/-{�uE�8�ǥ��1��k�rAB%�mP`�DH ��'�y��y��?N3�E��{;�pv��	�_�� d��/�t��I����<�1��g�^��Q�+�2�b4�$r	��m�9c�[��b0yjȩe����14�A�	rXB��RU��E���:�Z$R��1�����G�۹�q �G"8
��#���B50�r(�C��0�E�TT<���$�j���fM��ɮ�y ��sR(�|�8��JA!�L-�	�9�(��K����I�b�T =�� y{'S����'�c����<��\��{?n�$�+HT�lNTM�I6��qV�5ۤKc�������<"�lLU�9���+�W�[!���t�@�Κ������$�@P�M�#?Qt~7y[����H��k�~��ޜrP�
��"]����������併��}������LoǣL���׶�JQ��)�[MF��cz��/Q�:��F�_Aw��{��wK� ǄO%G��!�'��,�ڨ���9A�c��3��1s���ihA����o��M�e]��7(��ˆ�h�[���䑡���"q��@��@B���^��N�]0��f��iҡ;�����?咶hّ�����5
)x4�YA���J|�_C�{�N�]%��rਗ਼�v�K��JO���C,Z)qNc���89�T�Q9/�����.�7�0*��'l��Vi���B�x�%��@�#�����z�qO6�-v��ʬ�<���y_ZS,w=��Z0��m�!=0����sG���'/Ɛ�E��Q��C�3�F�ssz'G;Hqs�s��2�y�U%�.Mv�PJK�d��ݭ�
���^kƮ�f6�&yD[�:1������s�㡒�յ��ŚM��T�Э�tAb��瘌G�����m�Uz�?�0�K���3s<�g���q�$�ֿ�3�n�Eoqԯ��5R��3�j!����Nn�]\rQ����Q��n��#�� �2\#�z�œ:��F����q���i��i�~�a'�*�&�@�	�c)+@Ĥ�Qݛܮopĕ� RC�P'�??�J8p�<��N���F1QL�tЁ4By����KI^�T��{�Jg���Yak��"���ۏo\Fߙ���^�����	.S�E���(����aEϱ�Jc.6a�_-��8~�ûT7���qa"��Գ!�cA�� "7F����k������ �$J-Nr���dҩ��-� 2/l�p���]��j�N#O���[)Q��q7��O��b7r���#��,;�����c��B��̧;r/K�5�h�Z���Ԓ9I���ef�1���|I�D�h��Ӳq�\�7�;s}8٤J�*dߚ݀�>�v�촭>�v�g 6/X�`]C���oL�{aT<gxiP?N�@m���;�72�<,�(b�6�-��(��r,a䝴�N}�$�g  �1P��T���R��`�Bl0L2���/ʏj�%�%��������޸����?w��=�x���e�ܟ�v�4E�aj��b�[3��Gܚ�#cu������>��|��h��N}���9���y�R��H��V��l-:Txc�*��M3�q-t~`	*-b��}mN2�ЕQ�l�"'��Z�����)��(�^m�_:x�}��åEE�r	�p�/����;���� �֮ߏkG �� �3	��e�G�{�_$p���=l�]��m�>Y_c��˪���`5$Qv�
绎�R5{_'W����w������5T�Y�����0��ⱞ{3B	v���d4!�;V��'#W`|��M��v,�R�zX�<p��6M�7w�|�m&sz5��1�q�h�LT�m��s'�\����w��K���D�:�n�F�v3#�4�+�@M�Z�ܚ/�j��{(=�j<����}�����{+=�������ӣ��sԱ�ML&�O!�Ov�sNи���h7�h_Z���4��F(�V�I�������:{�(2�Ip�~���%��ze�ԡuq��b����c��r�&���FFn���<�_x�c�3�o��b�ʕeZt�Ɖ��QAG���"��R'�D���uep!�)n��8���1@���kT���(��?�?4ЗH���t��=7�]�FJ�X�)3����k��򞓄l����U�u���~|"�=�[Բ*�6,\����W.N�Q/�\�11��� P��{BXZ*=qS�z+������,�
��ZP�v����z�^�7���b�.�����8�R,���I��o�d=,�A_[}�m��>tpȶt����ɜ���)���/��s��<ٽVӈ��i<'���ViN9���#�rx����<���]����B��(�ҩ�KM�
�����_zh��h��/�@:7P��o�с�e����4�M��i��ā}��H�m��q�so'۷���P�Q�&'�!�Q09��N��G��#u�
����:��\���������C-��ޘ#�c܀ț���z<7 q!�1��Ҝi8��i��f<ƛ�l�I�$v\�m`�3y�Τv��V?P�'>˖�{����y�+��%�1�!^%AZ`��pIE���}�^'H�1������7�I��X�&�%�SS��v[ +�F���B^q��%��7�v�!wjq=k�봓��+|~��+1�����힒J{Xg-9u��8�$l�zk)���F��
���W�]�"�*��+*Xu'��Q+m�`�=q�E�5G(��p�g��9�gK�b'X�������3 ���b��O��.�{���V� {�Έ�C��Q��;��˔�Q
�H��:��@s��Ԉ"|�#�C0����PV)�"���M�N�Ej�E��u����!v�a9*�m3�|�s'g�1��p�U;�@���SB����o�<w����[���(���c�	�cnPw&<���~�� "M��� :�'��|�ה��"u'�NploN{*�z����J6�jw�A��n�)�4�S��4,�9���ɣ<���cNo��&�����!֡�����t�jC�6��^�cc�#l�{Hw��Go~�����q����8}(�F�gW�y����{wj1C|�(�A�B���^�~�+,F����>�!�	}�҃�=͘c�T�Hg�v��a��i�x;c��H�-)rݑq�{&�?%��Yh	�܎�Å,kX|f�&�ϭ���s.�A�R�Î�Ņ�N x�Y�'�u��,�mk�We��L~A������?�\_�z{\/�&D%xc�˸����/���� e?L'B�����4W\g'��$��1�n8>?cյu,!�E��G4�KZ�E�b��:�v�*���Y1�P�&�9.N��P�Yc@�-ЉL��w�(%n�E�Cz;5g%o���Tv]���݁��\j�	7�����HUٙN+��_��ٚ
 �+]7(>2��% M2Twz�V��N�pz�Q�c�.i1/_�y2��A��^[�u�ih1¸���,Y{5��$�|���%Wޗ!� =h�;��m�y��l����(W�՛7~2�/r�/�����l�~<� 2Q@an>EF`��@G��x��lo@:p?'%�����p�<Y7�A	���R��R<~��%Ÿe�="��;j�HA�V.oC�Y�*�"^Qr;,�&e�xY�|�bW�@4�2.� �n��ˉ�>j���z}S�WZ�c?�?j+��zS�:T�ъ&u��%�O�]1ۏ��#�nZ�Ϊܧ�D��6v��g-B揫�@��*8�6}X&	Di�kD ���3��u(���9����Q��u��F�C���7�5G��G�o<�k��8�����o'W��#'�.�m$e��1*�<WF����� �9���	�|��3��)1��Ձ/��x�ۡ�eI�dwX`bO.������$^]e�Ũ�3�[�������'�+Iwh�m��7����m���F$�؍<��w�J�l\��P 9�̣��%���1{Y1����Z��usI��ќ{�����gV�4sOMM�`��IÆw���(��3��΍&���\2%(������V�kZ/O�Ȭ?��9[ѻ �ۇ�+���y"4r�r�j��xl�6�����0��ņ��>aw��I,�Ԙ��ͤ���� ��k� �t�tI
��R� �� �K��!���R��%� �t7�t�����~�ץ��z�<3w̙����+�/�G�}�_�z��u���ߎA��]�-��J���ǖ�G�l�og�ד3{�ǏՓ�J�E�l����R��>�����x3W�ۺ���}F�hc��.#n$�p�^�[�&��}�9u�r3�H�4�5=�<b�s���I�W�s�N<�̠X�d��l�˔%�y�.�7�1�e�XWg׬��z�X2�X���ڭPQ�����I7u�5���W�+�?"f�~)c��'�|a�g�)&�lH=5'�	���ȟ9 ��a0=���r>��nx�觺F����r���<l�Vt�LS�l�\�Eߏ�������s�)b�bXL/.ל���碩������X��mq�Y�H�x���e<-�����������zV��zA�R8q��p�m\x8��oLL��+`�'omXU��L�!W"��w[�ͭ�R[Q/?;�<�=�
F�ό�d��*/�Ӝ��A�\���D��``�u�(����,y��%w��Q��u�?7:C8��ZIRp��	���FFD�|����r����7�����ވ� �����P���w��9sq���O�h��sG��e��V�!�R�%�#�P.o�t�_Niu��w��G�'�@E�C)���?��tu�LX�o���u�l&'x�HVj�C|eE�7�)�|��0�����H�w]2޴i�SDNm5�C��yB��/� �\?f��"���Tz$�"���Rgʹ�L������vC�ֿ��v�D��=;X�����c�%p.�g\lj�x�Z�g����b�#�I�R�)߇�V@|���L�MO�Pښ�S��h�H��s��u|�)q ۦ�k��Mؿ����|_�J�0���m�C��~�%�
8�f�;%|k["�	߮J܌Z\�𫃎������@��&�~��0#�����S ���kwg؛r8C���Ԯ�J���F��g6�%°�K���KϛZ!C�T�0��hf��Z��j|���O�V7C�w52@�\����{� �0���W���S�P��g�;�=�Ѷd:[���d�K��6hE8X���,��ܹQ	a<���>5���R�Ss��x� ̍ �빑Z>rBv4��q��߬���)�z~)���� �a���h9j���zش9��w�A>!}�����3 v�����Q��' �	U�����r�9Xa��P6u�y0�G��7U�����a��Ӈ3]d�������î�أa<޵2�\�QW�x(�sj�=pAOGIv�),�����a�~Q��i��a���I�=C+�ɕH��3��`�'��ޅ*��=��v�7�甼���7�/)���s/�(�S��-�$x����^M�����+o���ʊ�����S��TDo�r��)�☚��TݽpZ+���f�E�L,<�.��2 ��7ң�j���D:�q,�:b���#��|S�/x�M�v7��`;��-���gcւҮ�b	?�!g���@�/!���5J�в6|p��mט+%9�O��>�Y��=�嶎|� ��}o��˒����5Y�l�t�5�*;Gy�_��w[�8�p%��/��CW��Z ��}U��ҿ�B傴���ځx����D�)٤�n����Oт��A��nPo7X�缨����e[����.���Ļ2�4+RI���"��è�Dsޫ��2:˲���u���Q2(g>�H!�f�yu�s���������<DnăKG�³5���QCq����O��bQ5�L�i"�������3�U��o� k%�P8'ɫ�����'��E�!�<�!��Ѫ ԶKR�{s���O积���/XNmg"���VA��=��s�8�1�.B�$b�.Q��29%�{��G����5f���n7����%�k��.+��}�}�`�����9}���k6��K�jH�2 Jb�X����	BF� "�� ������q��b��L*�>Dy��/��k��?�Sz$cq���E5I��m/�s�	�3�](g�֔ֆ�P�73�N;�m'f�3Ԍ��y<b���{�����A�?�F�-1�(���%J��;�%���j���\'WR��=$�;�AIz,�f���a>4x����̤�e�c�2��ynT�����$�GF�5'"e�'o|�d������'~񔳄!��O��=���.�f:�Clz���U��Ywm�Pl�v*�� \�N�ҥԘ^yu�m'�F�Y` V}�����U�#Y�:~�lI}�к������#�#��:N���$n��Xh��;/�kjY8d��w<�~c�����o_�ts>�>��Λw�9)xDS��я�P�
�W�A���Є�p�"�I����V�CD�H$�����X�Z���z�lc�3?&H�����s�],>W	^��{��|\���DRO�98Rn�xW���2Ѳ��@�t߶g�U4/?V� ʐ|m'��b�A��gy�nĈU#�
gr\�v#�nt�<|�z8�ƛ��$��NS�F�����;�0�
8�᧯�Ya��h�GP+L���@�N��\="| h�[`��P�����E��鸆L��t���l�7�	[JW� xT���ir�\w�,��^��T|`���"�N��%�7�����ݒ�����]f��C-�B9�t�7䊗�t��L�S�V^*m������������.�ۡ+p���x�uC��2�jZ�|�ڞd��w{�"�Vڸ�S�]?�������&ܝ�5f���n���-`�s!˲���|��o�uf3��I�T��&x��'H8/O�d��8{̊��P��φ���'��u*R�k��D���9#��.� 	����g"R_�^��)��>p��(Z�'�j!���9�r�=kvq1�����$i�O�V�7+~��M�H�X�l���WV��O��}yY���ۘF#�<9�)�跾< �`l6Pֈ��)��.;Ji�'$��PY��0@�e|B�P{ϓ6z���P��`$�f��p�����*���������C�\r�wdb9X{c�R$��]�|�SpH�P�w���a�c�h*�#F��z?�,��U�%�8�2�,���Z�/F�v��W�!�$��O���-3����ۧ��p�#xSh�*#����w@�1�$E�K2�**��|�FF��1��5�nJ�lM����rFCi}8�B��!��*P�w4�I�k����U�`�yad6���B!sq ����b�������˨B��=���f��	v�+_i�G��j�I�&�e��0O�����l[��Y�١:�Q!�~�����Қ��#1Ԇ#*34�r�,��5�����`X)������3?�WJ����d$�@5��<�R�(��KO1]�}�gh�
C����V��䷽~��-���ʆ�)�4,A�d��4,ϻ�f'�����Ջ
�R���ȲL�!�����>�#Md}7�hd�X����D%�^�D_��{:�xR�p��Q��4��*�v��hxK!�tEg�#?����!�>��w�ʆz�K����8�F�����&}��B��}������ٝ@�y}{���˷�C�iO���Ҿ��>|i��ǃ�Ԗ�6���ެ��c���!9�ǥRt��p�ecaG��T�{��p" ?6##*���Z�硚r{�ގ�=wJ/O4A,�9�欫GT���}ĭaǃ�m9�<�O��*����A�-�lI��ȴ������ <n�xH�|̡�J�ПY���zD����������t���pdcʵ!�I�&���Q3Y��bg�^���@��F\�#]����g�P�+(*|(Qj�x;���p���"�+� ${�l��;��E;�§�9�-'m��Q�j�Ñ횁ǖ�^X���'*.�Ü8��u�n	��D?|_�<���K1���v��̓b�g��b����p�����w"�l��Q��T@����=���;(�E������(�Z��;��|���[�O���E޳N��70���n�b?QI�[���]֭Gq͇4�w@��a��UՠܯY�PףM�ć��+�.ǯ$:������R� � ���vP  ݂ �L��Z����(�[� ���{�Lb��<U���\�����ȟ����l�̍/�,N��02&�:d����z�]��C���(}�C�իbU�<�|���4]s�}����Vk;�]��#��
p�P
jA�{��aGě�=6b(�Z�в�����?j��l���"I4@�����> n	f�><��isIp�V�*�?�WЂb�����S|"J����)�j�n�j�2������G�g��UC���`�������z鿡��|o�(��u��Y�
 ^��C��!�J�� ����"-�d�����-eۗc���H$K6rƿL�'��q叓�M9��/��((��+�ؑ�P����-�K��Q�l�_:�#��_�X ~����M���^ʐ�΁�E�y�K��5���R�k�T9��fE��1��� "��C �0�W&���/�g���Ն�i��C�Ym��2 ;��4��se�����#��|�m� ������ľ�D�{���l��������Py[.�?-��c�G�G��֘��?��Qc����2'Wo��x��ܲZ������Sq Ֆ���y���H~����"N�P��2���`�Y�p�Igh��3FQ��u��pv��E�#���R�4��Tm��dA���}֭����F�k\Jw�s�J�}�c���=s��8!-\#	���s�ԉ����?��4@ �C�v<�n#�2�ɑ��wT>���7�cr\[B45#>���,ԪD*���**�e(�����e!�>�l���>cC�}l���q�Uß��m+���?��Kpr<P��X�Lj��B��L�2�J�n�x~�_8a-�x�37�L#�4۳= 6P�_�#y���w���/?4�	)q?PzS���>
RT�g�i������c��'I/౰�j_�^��~�Ė�CZ��+���C����-���b[�s!\�F�̸�b����r�K��⑭`�ѻ�<��D5˃a���4�P�˨��u���7�[؝�r��`��#�]DM���ȁ�8#�`��s2m&��-�4\s��:��=�Ž�W��j=���.��9 j��멹��g���������N� �ՠ�4��K�]��.�vT��^�\f����/ܐawh4Ƥ5P�)��8�j����:�t�կ�>	�?�c,)���,&�%<Rx�.��X��[
BV����/�p_'�

�8������I
+	il��2��9,�N�}��1ȱjRҜ��e���n�Tt.��<���t�v!���=���ߑC�^"�!҄?A77~L�$����)����3��Ѯ��'r���y�`�x-�vy�z\����栾�������@��/�܆�1m&�r�|��Ы�i��4pA�e�)V��!r��% 8)���qƂI~�zX
K��̋����
p��#n�_�U�~6X%�'���
�5�I�٪0�v�R��O]�U��ۄ� ���)̓����T���~�w*����0	�$�����2��=%���8�i����/
�XH@����,���!�FNy���N�M��R�D�߉a��\���͑u� �5�̑z|_Im�Y�X�Ź���)�K�p������A7�}9
�Q�|���W�����B)<p�Д�4��c	?��<}Ӈb��l��h�~o
I�V�]��-(�J�N�|be�g�ǐ.{�JbS��t������\��(_[�U���{��E��_��i��ǈ��\�	]ܑ��k{�"�8_�E��Z��N[g	�ew�!]\D���$+7z�so�Do�����⠹5QMgJ��ꆑ��\I�?U��πE��)��rY���r3ۙ�FSJ����洼&�	�Wd�Gx���@�}�\Տx[쐣I�p�uj�2k��c!	I|x������	r�ی��Ƅ�G�����#F�0�Y���+E!^dr��iXU��gG�9@�o\1� ����S�o�Af�����-�� Q+��e��En ��vR4p�cȟ�1�,�b��s�{~����r���/R�d ��բ���/�Lg��6o��aJ�1�\rvƯ�>Q]8v|�f�Q�xIT��f�!qy�T�D�#���i�s�Kߜh�&������$��G�1+I�cD�Ib#t\��v����% �I�~�E��;>(�l���������N~��?�*�5p�&Z�t�>'��i�Z ����{�9ldKz6c;�`+ċ<��� ]q��}�m��WV3���X�q�
#j%�߾���s���=J�8ɫ0�>
%�A:��U�]��k�Y��U�+~�j�I���~T�*����1R8,:�|\�>�]�?i|Ɨ��̲��l�g�}c�!�R7�����6GT�Q��V�Y$��B�;S�ۑ37����l�c:Ŏ��p6�u9�f�8��R�{�>{�4��&F��˄ܜ�U^:B���3)e�V�0�3��I"�;iU�:T�B�]z���$�mԄU����E?ɂ*Osl#��h�늣��@��z�KB�}'��ȵ쮃i�'Òl�9X��RLwf�y��|u��,����g�i��Hݸo1Sȧ����A;���]{x�'�
�C������7"�$T�y���1E�u��9��RV�jhޥ"�j��y�y�t�jQ��W_��f<��u7���7q�ȝ������#C:�T &V���'���l|є�s���j�{!߾�o����g��,�P�I���/���G��i�9u�"kӆ� �˕U�$g�2P���J���5�,D���|.����u����uq�C�����c��y��N�ށoX��+1KIb
ޏifj_3��#[���c���/��^|�>o�p^̵�e��u��t`o�#V=�D�].
���gg���q.��P�e[�Y�I'�N�1�!``�A2����Q�~$ZNQv�~֞tch���g���ۥX�����c�w�6�m $�dqBZ�����h3D��޽��_X��D�7�Z��Y�_����ɂ��cq������l�D�S؆�̠Β���0q߶�0j|�؁��$�Á��\(��O �ſ�E��D)�5�}ڌ1n4���ʠd[Mi4t=�!^H���b�%�hV���N��G�^� �-�M�~�ZR}�ء�E�|�Xh���!�wm��z{H�����C6�,i�j�a�!Y�-��=������,:��7�jhəv��ʱ|�l��K£o�-X"�mD�s�	�\P�S���F��m��?3�
"t��,��Iǘ��̾p�����&@~��ZD�0���]L��M��=���l��Y����P�"��AD�+���T8Z6��� R��u,�r>3����w؆�������26}h)�g�pHd��z}2��+�R*��p�Ȗ2Σ��1@$B�mBO!�&�rɻ�r�K�աҾ�����~��YȌ��>�C�o������2B��7�Ή��	R�<��pz�>�:5y%�$|G�4����*�;��`���!)���S(f?���P��m�)�s_i^��:��2�#Y7��D�}9G��|n����&b)���G[}.<�ġx}G��|�g���������j(�-��Yqڮ#蓬W����^^�LY�N.��ʆv��
�l\�B�&z<�G�Ds�Ԧ� 9�/�N�'�Gn�#���Y��JI�W.��a����z�l;R����Χ���@۰.m.l�Dn�u�3$r���O4V��VG?���ӈ,�[�gU\�8��^W�������p�d�|^��4D����Z���
�1��t�J��q�Y��7Јbb;��U}��z��!�Z���}t��h�\�x(���,~�q�<R�٪z^J�M�(���uu5�y���.X\p�˹Δ�z/��H����X8��k���x{�� �+�����{D�u�c��4���w���S�M���+��t�����G�}�Y���YY��茔zF�ҝi.�a/��U2�Ly�IZ���t�O���Ò�d��˔�Ƿ귏�"�e�=�±#�X��i�TM�s��&�M!�.��{���Bh�ɩAJ���b�W�#��r7.`Ʒ���ڀɫqBV6u4�$.9���~�C��E���;��J����<�*��;*���=�u��R��a)��x���-��|��( ����wJ���#�,&�BS���M k�d�|�2p{i/��=So�#�]ߖL�4�Ǡ/��}�{�8�x![Xa�wz�
vz.l�=��YjV�Ռ�?���E��8x~�!_!̅��p������U�C(/�{dY]����NV��H���P�oZ�eO�ӱe
7>�#���� �E㴜P/��ϓ�u�Jn�tM���u���S�?����=�n�LecM ���Q��>��ld��&��̈́}�=�Q���*��C����c�tE�0�,P���U玌?Z�����'�1�1p�^��JZ�W��e���M��4�TGxU�c��K&_�Z�L��0������)@x����
�E�-��3��r4�+���4ZA5�
,�տΈC�\
�����}b�{�b���w�(��Y�v�岺��Є㾳�Hy�R��#����i����"�S�3��c��M ������3����
��A�,�Q>S�5St���~�
T���_<����w�~�+�NзR�|�y�Y�<�j˧�K�����4i�Z�mqƣ�tAW .��^��p��z̅>�h���<L�Q�)Y������C�ݱ�ki��JG�a+6(T)�>���;��G�|�Lmֿ���!�YT��s\���ѳ|�e�O�\�UU�+���1&������S�#])��������K/����.c$r%��jօ^�]��d�-�S17��i��vf��Fv'ZP��<qj������/U��\jB��-vN�0G�
�&D�xD7;(���êp�x#�puR8M�0[ZV_�seQ�M�}�"���͏R@�M �i���Z�l������־՛Z��m�[(3�o���Od��J6!)Gg�ۇ�|����T$��;+��N�7��=cF��ФƸ-�,�6�H�d#:��q�3=���,����ݞ���VY����P��g뺉�1ZG>@� vP���9�"��b�J��솓	ŁrL�o��!�ܞ��k��e�#־ۚ�ʀV�Ջ�nˌLJ�v��i� $�w�U��Y�Q����d��lb�<�e��/ih!ĸ(�UP��}�j�Hx����`��#�*OMg����(��{B��=e|���!��F'�n�h��X�^X�L~a�%����8T�&5�<�:RQ'm-�|���,�^$�}��x�.J@񖥩G/�/��'�Q�E�2�%u3�QH�ꀤ�H@I���ض��C�V�eѿ	d2��_Aj���x5�P�sc�ݙ����O�\�B������'����\��?^�=Ѯ�����/1�����j��(��m�clZbˤX|SZ����e?<����ʆ����km���Z�I����@I���כ�#6<�U'��%��U���M�$P��3�����C�Zzx��HG�GXA�mK�d��9��t�h�c �Q����lt�U��8E�=�q�����J
������ ��h_7�&K�ks.����ר��w�@��J��(�h�.���lVX�C,����R�pe���$n��3y�Kđ�'�l�VYp�bT���"�h
3\�"�\��B�HƜXv���vB�Xn�+-�֑ncI��Ф�#�o]�Ur2�n���[��^#]�l殜�m�wa��ůJ�3A�f�q.Y�	����[��:�R�~.�_)>o0˶o��U�eS�X͑;�F������k�8���hA�g��k�m%�T��(i�(�z\��r-��^Ǒ�a�6��VN���߾��?q��v-a�C+^>�@�AjPHK���)T�8�3B�G��C���T	�c��"��mw�����F����[|�≳*�o��u��P��oy��@�A)iܺD���݊mk�7�S=2�d�rE�B�����k_Q�� j2����LtR����"������~G��X��V4"D�e;�y����4��4��K�Z�E����X���CÌ��1��v���_!�N�3�֚�"G��*��'���s&�F�jaI��F�O~臬�B��-���)/-�ۈ�B
� �J%��P��z�\�7X�^�Վ׼�_��N=�/�7!v
Qc�^����|'�}�<�յx�S7:A-���,Gr*U#�W��-����:��cw;���F�XK� ��H�ȩ��m[�K+N�q���}�#�C��27����6��͌R����?��7�TMV���4 ��a�9���kc�r�z�L�0�aT{ν��8�UY��e���8PH8�1P(��d`�iyM@�+��5r1��&�&�ݯp��"}q?R��� Ӊ��8�ƿ#a�\?⠣�*&4��	�2� �JG�r��j����;���I���>��ֲ�Z�X�
����I�t�~��n�
�Xb'�I`jH��[=�8��tCTɣU�Y�'��pp�wj&�s#�o)��y�Ó��p�#Ȝ�'+O���(]ޢKl�!0�"�d~	=|oe�R�75���p��i'?�������őh	A�j!�E��������2r����-���5q��/衫�3q��F�-K��`���6����eL�6�dafp�� ���da<�/�٫�s��Z�(Q�
%���Y�ɚAg4���hV=��%��6������sӹ,t�^��g�]�����;��R\�a�+,p^�����IA����Tß�Y.��8.�OJB��GJ<?��&HZ�5D `�=��&Y����N�G�N�F��h��;!8}�u�<+����3�Hb�-���p�n�7�rK�k>]�=Ω+Q����$�,�}�͞��j�2ॕK;b�#�MR���S��Ֆ�j-:�r�J�+��l; ;w�L/���������4�1��y�X;�1��T^� �����2$)�(ڶ�D��ma �j��:���^�^//��lI���~�19��04�����8C����{��[1j��"B��r����V�z�	�V�����C�=�����5��}��$j�j��!G*�J:��#�aۉ}���~��/�q���Z��P[�9��df�۔���%�(�&z����o�� ;�C*+�&g\�(i_�a�Դ)U���<4��J)����� C��8���q�p�YPcŚWɄq�:��R��n7�	{�K=YDw�ͨ��>��J7cu�_3��Sk�����y�3l��۴�f�1�r(}HܺL%
��0�:������$Ьt���YHF��lM���;�K����M��8���6��`��ON�o����~w%�+we={x�)џ���a
�<ip%�+U�dv����a��2.j��l��8b̐�z*Qw�E�D���!��_~�!�L����x���'���PG�����o�T���c��W��z[>B|�\����,g�1X�R��ߪ@?�9_���v�K����8X쮎*�+	�ڢ2l���s,��S����� <���)q�����Il��!kR�1B�]m��A5��豽�߉�G� �Bt�d��QN�Z�=��n}���8��I��6f.�����z'6�RM˔��@�!E@�4���>c�XX�C�Z��M!����q�uu
���l��&���HՁ�̈́��S�b%>F��Dҫ��)�[Y��0*�W`�_X� �4����\�7Z�C�G�m����;���|��;l�Eǰ�,� \�\_g�9�0O�V���������	4Ķq:`t<�����t/[���n���0�S	�) �H8+W����M��@�l����-87�Cl��,�|>x�e��:����h�C��ٸI��8�o���Sr�/O72�N ��%Z��Y�UM�Y�;�"=S��A��ąz0)�|~ZA�?=��e	�act���n7���;�8�󙟃ru����#�D %��?ꧪ�g����y;�¾�as�o4��)QزB�ps�I�au�VR�MC�7�]t�W���`������G��Sϰ��$Z�To��+v�:��e��&�C�q>D���p�U켂�	�ȣ�oG̟��Т%�}�L\�o``�C���vo:��>q����\����d��=1����U��o�ly����z�2��t�+�7��%Zrw/�|��ᠠH�{�Zަ!�'��IR�J��x�y�x)�P��J����"M�j�"c�@�b�����W���`�#-w�K�r�;�=��Ͽ0 9"�@GWh�;�9����U؛4��+6�?5c�WG~�<�Ռ�'���M�
�o�-�O}��l}���eFAb���"�I!#��_=��w7�ߕ_e�J���&#R-ȯ����d�P�xi���E��=ɕ�#	n���i�l�Q�BW���~?�Η9Z0�y>�{��v���󺜞������K�Xp��J"��C�@�����&@t]6��#	̊i�X�yC�48E����݄��h�n����?o(�,���]O���׼I��xCz���/�����׿�O~ �Q�Jޒ:k�i�<�D���L�|�P2���RW��v��țkC'��3�s�*}o*�~~���K�[g��y<�}X��;!���ŭ����n��3�>$�t����S�Bq�F��4Q*��X�U�od���@����W��Aċ>��(y����[b`���)�9�b���
[�V�J�
�]M"�:ET��Y���5�$ѻdr��Q���(��#�� ���5��@0��U�jIMV��E�:�E��Ws�	0	i�Ǿ��� ���S���L. �ib���h��?<d�P�
�?�y������x�;���_�+�:@]���������θz�2>�a��G���c��o�`k$�O�����);.��\�B��_؛�b��#8>e�ی����L~�^IoJ���4�0�>�RϠ���"�}�Rn/j��T������X�����D���1�^b��I�k�!�Ǖ�������*?;�*9�$	~���֜əUG�ڙ�O׆��Q��d�Q'� >�Pґ*=V�c�I2���}���HQ��*��Ux�3F5N/|�"��(��nc�ٚL'�8�����o�u��H�,c�����1�7C�D��3]�>|[�=�)�Z����"�[�vh���Ԍ͠l�T��$����\��.}�2L);�7K`u+Oz�K^H~�Gv�S(��1��ϧ��9<Z$� �2�^jn���i��p�ɩ�^�o�� ����	F�����u��؛ĵ���OZ�5�$O��&)��Y{�E=b���$9)[]�0�S*$��o���޼{��%~}E��5PR ��#{5m*�S���n ܼI畦���g$H|#�a��\0���/��_�D|S>p.7m��ᔤ 4�'[�8�Y����3��U��v�D/ɼ��cq��;�"���-�E}=.��F����ng�4�8�I@)�gh�=�r*;({�)ə~y�f��dhv��������ԋ�=�Lw�?��9uTy�>0����4zQ��1��P��*1W|�a���d[��{.+=�Ip�=zGׯ?^m�'���q�T�c�	�l��X)k�,k~e��l�l�H[�l�bc��t]��h��9�h!F)T���ە͔�Ǜm�6ƿ�"�T"��F�Q<�x��6|��U����Q^e�J��6�b��XMs�z����/_�z��=��*�I���X����=.����@F�P��J��=��YQQ4�OU"CS�t�S[��k�TG������E� ^�e�VBZ�LTϻ��+���͚+���Ë����DD�j���� Q�����K���
�5	K��Qְ�I��������o!�~X��Ԁ�14�'0���2�~�r%�7x��`c��Ȭ+�����\�K���L�<�����J��Q��p��(�k�J_J˗h�4����h�p���#䅬zX��V�㹱uS�s��mU���c1�YY�n#����yS����������*G�w��5���ݗаj\�H2�{�N��+��R�ya�J�r�q*X�	#�l�M��j}�a�d�U��S��[�w�*��Y	����oCDh���zoyU&�b1/����l�!�9�Ǹ�4g��)��f3�������OO5��+x�[�% �=�ѸbR)�֙w����S%/ƃ�څ8�xU�����_%P�|I5��g��?�|�W�⹭�;�k���$BN�O@�;��(q�����D�o��~�QzM�_�-�)��24t��]�`��m�_�흎5�V�Kg�J���2�Ci�xn\n�f�G�2��ʇ�D��_�F���J_�:fU�qm�f�2G��FeO������DHu���\*|f��g�ݻgt�Y=<�h���K���"�U�4<�ܮȽ��5Y
QJ����+k���1�ybh�9��qxe3W���Tr/?���J�x�[�␺i�MEm���j&E��`X�/l��S�Ä��;�V�1�����Ξн'�{��+?�j6���:�_��c�5�7����9Uʁ{���s9����T��Aƺ
>c'���jT��e�RCƦ����Y!Y��p���?7l��?��DI�����\���Z'���-�I�>�I�UnR�7\��5g�����d�=�sZj�R�7�W�#{�@�lׅ�p:�7�e�7��j�S��*v� ��F������y(�Dōz�gesɩ�����Q##$�n�钴TO�Ms�2li��>I+�9{�ED��~�-g�$S2�OS̤�
䍉��d��e�?�Z�A����	���}.g�2������X������o��s���U<k�8�'�q.������&~bv��ўc�'E��|��^b,<��0�ՠ�ޕ�׼ �2�!�#�4�v���3Hn��:.���^�p�h�(Z���ܷ��%`Kl�Z�s�O	���~�z�Z�M׎�p������S9� ZY�U���J>�C.�#zb$|	9��5��R?�l�
���]��	/�ٟ���`I6��^��r��<����mX@����B*4	��fQ��hs�C�D�f��Ww߾����Gg)i�au�<sr��*�;1���#�&$�
�6����?�������+�j�XIM5�x��<B^�CJa?[d[��ںF����^�-K��J�4�l�S����k�P�\�[��R����#�.&ƳV�Oú���Ui,�(Μ	���,f�#��ʀA	@�������;,5��CrAq�%�^����JWU��6�]��/}K�s���^��C��}�V�N�nI��k���f�d�X{�&>���_� 0�4��mX�Uϗ�~�J��nYĻ~���O��л���w�*4�e9�>g	4�?��H$��ym湧0v^�f���&-P�LY�\�췱�����&U�x�,��EJ�N�P������|����/39�
J��������s�x�q�C��hm:(���A��Sw���BuQ�y�D�LwL�O���UE*��}[�ż�E�p���b�V�G��m.�X3pܫ>�y>�%/Á$C�������W&S�����/ԝw���0]O������D�o_f:Ŏ��P�=^P����Q��o�Ȯ�Ѵ)rkkX��^�4 @� �F'j�>Wz�9h�����߶�該Q�캬�I[�=!�l�����_�ƮM8j�xL��Jՠ+_3���r�ܹ��-K�Y:q��(H����r��2�j���5?+�%G>��� d8��qI����-����"k�g���}C R�`�z����oƮ��_®�� j�[��w�+j|�n�@�d�Q��pLF��g�4DG�߶��犚��+�Q$jn��ؼ�,yMt��FX���N�jz�o#�H� e��ٶ����[V٧T$�ܱ+lU��?��A� �����ߎo?9���g�}!v�c\z�i���qq=��&�n�F����y�&]�v'�H�:�1-��Pi�9%�
�o���,֨(r�s�V+��{�~Js���/1�=U>�E�W��&?�9R�&|I�V�/֬��R� ;�/�hEYʋJ�~������j(b�*F�C�uKRk�b�/��s�qn������w׸P���d*<O�1m�_�$���b�
D����$���(
�����ˆ%��8��_���J�y���U=��+F��x5D�V���wi�?k�R)�Zq��y���������-ZNZ0����ܬ�h~AJ �'._b�;9�7��p�Mo�y	��#�rtū��:6������	�S�j�._�~�MkGP^��w������uEd�r(*0�B���)^L�BVP9�0��i��=�uz��)~�v�f�ZJy�`��L��}������!]t��U��5�	LR�o�Rh0�((��V����wF�?$<�2K w|�5��x��:$P�dZ��{1�0�im�dR�M�����p�0�1 7��WJK��o��*	i���j ]�k9}��}q�ֱf���M������%,յ�u�Z/������N�a�[��
��HŢ�3=�x��6�:�o�E&&I�����j�}���UϘK^v��kG��hn��m�Ӓ�h�X�8�;Q����߃/NEW7��)��i:��C�y�|���$Eq�L�WaOm�4jYT,� ���_����BX��Ң�[���`����<?(T�!��vOcĺ&��n$?���ְ~���PC�)ďE�?{$�~�KS^���_�=)�"��� ����������^����h�d��*kZ,b�s@bӃj���:(�����[�?C��܈�C�A�����v�:i8�3�@��!?{��︅�챻�1ä�x��_�&lK#���W_���=����������R2�R�ݩH7��R�C��HI����ЍH�t�����f-��0����O����7o�'{DJG뻰Ф�`xVVYȮ�?�	��W�����k��H��ϑ����k��N�(�;�a-6�H� ݜ��TT�Q9`xIdӊ�I`�RшH���@@(�N\�w�LK���:&�T�L�&�c�S��0���z	��<����[U)}�w����<U�y��Z�L�t���<lܛ��|h{J(�k]lp�}��V�;M��*�'@�e����ڀ�gM�gF�Ly�j!>I>�����V�����2�U`��r��e	�~�:�TX�{�U~W�`�հ�Z=4Ht�h%���*g��Ap����鄝�O{�}\�A^Pt�+"�凵*�f�v%�HW����j�y�� ��������K�y/%��ޅ�پ~8���fO���&��É�M��D�B0��k��h��qf�I^n����[����'�
�ж?y���5Uwx��������y[�H9|��Zwjp��H�]�����(Î���׫�i/�U.	��[��С�`U��y[ۖ7)hGn͝�Ue��S={2�)���K{���F�?r[W�����2�����YK���<V��x�>6\Iot�Mq9�yN]���ܰeB�/��$��Gp虄���0����+����4"[.8�*�V`�Z�B���Ք�е.a���|�)�a,)��:6Ф����]��C�w��e�OP�� f����{)쌳�bS�^4�R��ER�;Q�m�3N�#\���垞ܻ�7�Օ��3��D�_�����G��*��7�!�4�=���=���h}�a���Aj�o����Q<�GBeg�P$��J�2��0�P�?����m��K��:C������]}�m�C����e������u�?7z��h����<p��ݪp��l�F�}���1�}�g]�3
�'ɞ��wh+�p�0
B�衸5���N��H������:�%9�6O6iY~늪�R�,��D7���~]\ݟ����<������@;������&��vVt�R҈����S�T�n�<^{��A����ׅK��!��?��J�%M����6f�U@���Y�^{f�4Qg��@\����}���dg��"��qI�^$p��I�F�Ȏ߸^N�����悁>%7�o�+'��h����g���W���dE�����eݷ
�R��Ō',���w�@�.��\�	12��r!2�a�f�������)�ƒ�=��d84{T"�T��([�z8��5�L����Q���ګ��I�	R$����&���gӐbYM���������#��
�U�A"�/�q��&"�ݑ�Ί�f5CK��2�\V��	�
t���
,l��W��P.��4����6�T֪�GDKB�/h�I�A��D��w���;KWk�uJ�:�t�i�Y;�� ��6�S�#�Ǩ��NiH�sz�F���N���s�Gu��i{�u�@.L����UEx���u�6|���0.3�ԫiD��E��HR��W��,�K��ZP��[��L q�Z��T�l�L��oB�z��
R�" 2�2\'O�V�.��H��L��4�M~��L8�g%ET���
c��Z#�'��� ��p�v��9�oЃ�H�������z�}YjH#z�x��`ά�Xj;j/��Ϧ�Ҽհ�YBvT$���B�5$طV�T�Nտ+aԙdL8{��� #��?-\X!A}��ٰ��r��;��$w�	�L �;ۋ<=�t_Pn��֒u^@�������	~�R5��-?�p�C���7�v,б5mJ�7�J8����8Y�+�ܐ�#6��Եn�5�?���uҼ #��Zϯi6wk?�̥�� �3������֔N�w�$�h��k�36�����հ�: ~��fO��� ,(�}�<��w�mN���ԜA��,��� �ExG1q����P�^|���zDt�ly�R����h-���p�^�*B������C�(���
�UF*��[3���(�6���* ߩ{������)K��	Rh�C����� �}o�F������@����{��2�B^��z:k��Nn�3,��_��ʴ�^�h���*��N3��яt�rY�l��Hn�G��x���V	$`Wy�<_�EzT��]��Ԧs?0 �:�QOw�4,�i���r�0qȔ=A�%�y�p�(J9�r��,���I�d�+��l,��,��B����A�T.A�A��p�֦#O0�9n����x;zZ�_޼����!a�	͵g��oi�)�����+~�r�O�����YU�k�>��浩�C���7��7��W+�ޑ�a.�HA}
���s�0�V��%[�W�|hݲޚ�߸�NfFp����F�=��	t�&q9���f���	��}�e�1|�
.~hW�I����8��x`����-R��&'A�3$���ݬ�W��/�*��%����~�p-�\`�
꒿�}w��~���(�ڞ�lԂ�!)D �9�JE�o���b�0��!�w=�$e�ܞ���aP� �;�vnߗ�����.��j��}�5ݯ�C�Sg[� ~i-!0!%�{%|�Y�q�_�z����r�wCN�3v��n'�Ɲ��G	����Q�-���'A���\NnB6;ڴ�	O� i<@fн:��sPP�t�0'<'�j8x����':]7�s���٨�rKiH%� t�i�6�׏�;�r��A���"�(s�D�B�d��2D�Ѱ2}x,fH����0'�	��>��-D�&�i��������ɐrY��ϥ�ł��e��j�(��d��e� 	oᲣ��[�dg������Bݠ������d|Q0�p��C���Gp�����Jcn��нݯ&�{���ȼ�
�*;�Z�2ip���x�p ��J�����o��ܖMJ�OjEy.L؋[�Q�tg��KE>��y���9�mT_f��V�,Xm1EG
�����䛽/@�\����s�&�2մo��h���*��fr��;�C�!�x�酌�ĖahR���M_BY�MHѝУҒ$����d�
�/���n8�&�H��H�f��wJHx#��C$��t���k�(H�6�#�z���W��3�p��%d�@M-�Wٸ�
Q��v8�1n�ژ��8��v���3Slؐ����m�gR��{�I�G�����;��@�~�<i^E(c\��BS��v�\�)�;�:b�GW����LL���s�v[u�־��U.�pB����!PO�ϖ����(`���MΆ��)���Q=������D%�a�w�j�V�J�̋�p�S6�D2�-E_���*HE��{A9�`Is�	�����~���S�S؉_�sv�� �f�顭�G!YLpQ2_ٰ�N^��Hr�n1��[8�߅t��;eǔy�xo��	��.$�i���\ae�_���֗H���$_��~;N�,K�8l��S��y������&��ؙ����ggRٶM#��CD��F멾u���C��A-��7�Z���.��04��A
��r�6��	Yd�̌q��I���S����~PY��\��uƃ�缙�����72֩G}���QƂ>t�_�/xE�e����=�ρG�/�w���;�����DIU�+�/�k֜Ï�������a�\]�i T$/�B�����wࢄ\k�:�����{�޼����V�G��W%�q�y�;A�@Ho��Y�$[V<=+�Ok6��й�w���h���Bl�d?k�,x����"X1Lq���YL�*�\�X�Dpg��/~<�����TQ�Ζ�(�碢�3Q!�Ĺ���,C�~Wo	]���&�A(�٢��A��~Z��I��%�ݪJ�	{��A[�p�y�W1|�<����ҟ2�!Ð(�S�x�.��1��1Y��(�G�iO]�&�~���妀�������˟�`��Nj=��k1x��}/���L*���d(M�Վo��4�g�k�ZL�]k�����*kA��f���Mz�E��	��0���0�H͔�Ϧ�Q���Ad�a6���p�ZH��QﭺOQ>���0��~�OG�	��Ő���*6kl�76GpN:M|���Kh���Y������F�҄���Ӊ7��[gi��A3��ϐ�F���+k��eD�C˴i%!Y��j��eT1��������c�j����L�9,����������]C�w��ƫ2wK������5,a-y����S�qs|>��������i� Vy��`�<�����p,�fD�h/�g��Ղdw������o(��{����#^�"w�'�-l��U����&�[wM��]3�~�p�����<�K��8I"���a�t$��u����	��IH*�E:��y^���9�6n?|�&O`=�(_��e�/�y��_��x��5�`���l�7UA}͊��CQp�4c������Z,���7?�<2�&2Iy9�
������n���Acc�Ew�,�}حVo^o-�\�.d���۶� 	�v�G�raXc1u���T��F���^�Ԟ~s7�=��j31��Ǯ˞��wOە	���� ��,�h�]���*�3���+#���O�[�ܵ=d&�{�KP�=$ �ʕ|��k9X��W(a&�.����?ڕ]�=TB؏��'i����Y�>��, 6&��R��{Ԓo63�i�����las6���ʭ꾌ƟZG$�a�x�W(��o�be�Q��*o<O2�a�B�T$7�7�\���k�Utz�B0��Y��WcN���Ԋ�,\���'�<û��Q�Ƌ?9f��C�����,/Oy1��KskyI	�e�_7�j��Ek��5�^6�_�v�2�)��zV+o�t�M�o��ߟ���������I/}�h��|M��I�[d�f�Ŗ��{ѓ�Ajbk�3�1��n�"˥�r��u�@^�.���R�1��`g\��L�=?c�b
c�d@y���Q�M���FI��b�\ 	���%&Š���
�c�.҇��2�����.��f;R��e�����$�*��MLM�r�koz�Bg���~)Z���Z�5q�'t��7�>�9�z�W�4�H�fc@�,�bl�	�܊���Ak�-^LGY����� Qb)bE�TP���Š�Qh���a�n����D�ނP�z�-���i��s�~�<���}�;&d��Wf5˶�
X,�\��b݆��$�㣣�#%�u�:���b�8���7�ނ���?�P^�<`��;���f�G�&`�p�(v���&��&��apU�Z�g##M��ex<���=�&���b�G0+?�4�<B�^���i��[���	�Z.�o�1J�<�x��M��q�G�c��<�HBʻ q��	�G���^J��q���l�]W�_<���RK�������%Xy�h��%�A�}ٱ��׵���?������im�vN�+s�����c�Tꌐ%��Y�ρWR[�#�>n�w�>�^ɲ4y{ŏ��O�	dH������93�g��$�j���aC˫�W���ӂ�;��K�/���݊W�G��b��lI ^�X-�mL� �p��m��ͥa�ʓ���+aYq"�&�v�����@�.&ܳ�7�^��V�bӑ)7��?&��W���u�#���ؾ!$���4��
]HuKϯ�T�ZI������Jw�4�=eip�A���ɱV�I��0�4��S1v64�S1�|R���Qa�MG�ʶ�fɠ,G�FU��\��K���Nn�7���Y��u��j�/����2<�[AB��d/8t�Ύ�e�"ܸ�p�b}����q�~R��m �.SiL�+�=e\𧔤��;O�|�g��*R�eM\�Z{�����34����Ino����H(�-^�����e��ۇ�Bc�u@����������[�pRʅZ��>�=dG^�^��T1���De�-��1�;�Y�Ծ.�f�򗏋r�`�	2��.� k�ɜ�� N�Q8ʹٲQ�ޮ��ħz:�ܶY���UD ���`��,��:��u}�hP �3��&���u4�QA�zo�^���F���5�����O����u�=bV5�*�7��x�f��8���!M�*Լ�_��Z�.�*�F9ps��q��My���%Tq��퓖j�r�"��Y�ȴ��q��A;�쁉�T��A��G��FT�薼��Mzh��i?�����c7v��EV���K��y����(��,��,���R�I#�xE�ˮs٣2���=�eg� +�5�記�7�2��e�p�A3�8
�R��T>�늕� ]lY��jƱ�ˈ^̮5A�a�_A����Ƞ�@-���J���]G�w{�[�=nLtE��L](�}��Z2"���ݲ��h,({�-V��u{Xc�u $+K���G����a.���I��z���@DO:���j�+`gC��D~R�4���R1��8�%C\0e��㣕�Pel=���ΰ��ٍҩ��Y�����f��f�OzJ��bg�O]��T���T5"#�R~�բ�:Q]������I�6mƖd��P?�����^�
'r��&V�2_�ܡ���W��I�\s>= I}*�C��;U�]��Tf�;R������cZ1A�����[4�y�kκw/<xAv��"+�w�9~������!�sw(�˷e��O�8�ؙ��s���v���VV�����`����	�x����-�����)���|�3|D�'�����@�N$���-?j@�O�LnH�(Ś60wo�*�.s�]���`����<+�:6�w�S@#X���)ͣjq]�_Ҿ����a����m�T� ��v�ʄ�t�W�͊^����ʺ�m3�����Y���Ƌ�����>�g� �j89��ڢH_��U��)9��E���.f����#/$Q����p;Q�Ûf8�rQ�3J h�Q���	���dr���q߱�;���0d��J�*����}N�V����Dk��_�7I�/��jAl�N0���F\*x�R���=n���c���e�]0y���^muɄ�u�Sp�{U�gQ�����+�=��|xj��Z#յ���M��k���:=���z�Yd_��h�C�Uw���qQIW���<Y���d�&����{0�M	)��W"8�1����r\���I��{������ dZڏ���J���U���(��]Cs�<4qF/өi(n�5;�(�;����-ߴ����XRrǌf�Wn6��gP��vطfԎA l}�M��
�D3�au�ؗ�ԋ����d��p]���+ �	��,:O�
��Ļ���B��Cf�`~E�lIS��ؠ�>��t�e�Sl}(���JF��HpPvn��M��̕����Q�J���#��I4^��\��f1=����q�2^,b�����^Ѩ��O$�۶��]/m�*]הS`�t;[�s)[��ۭ���M8�ʿ-k^k��Ę��|�Ԧ�� �Y��nn�dF
Ȣ����pG�DN�0.�������5��c@��^��B0 Xr~z�^��
j��"�#�X5Aq���:��t!�aSa��iĎ�X��]1��S�U�Q1��|�'G��+k)H.��� ��V9��V'9	@@��R]\^Jo�$����W���v�������R�����?[��/�DW-;�� ����g�/������Ї[�<2N��N��v"��_�o�yC��6�o���TH�^χ��XdM���ˠ���S"�C����b��gx;M!	��A[���X�[H���bW�!��Wq~<��۲[�Q��'����nض���y�"��# Y����h�*�2'D)��3��MsBeW�"J�f�L5���X�L�ca��|أ��1m�> ��t���-���p�3�(��C��N�ȳ���ӁF��H�X �P�[�+Nƫ�#}��
'�P0�J�� ��`o�3������Vj���r��)���0�r�Sg7��\�&���iz�X�R��a]�+PG�v���Ԛ�����X����<��Q�2���c��D�·D�u�M�Ĥ�.�E'{m׎���^�?��c�B0py�Y�k.�zR��x����rS�~�����0^�WqT���K�].���K�Ql݈��
�J��Ե�-�gl92v��ܶ�
j��������\2�RD��]��\���)�or<�Ԭ�.��`@ś����2O�PF��e���n�;����"�h|�\�o7D�f�0����+s�uf\w���]a�(tAf�2%�T�l�Y�O#�l\�}�����W���30�=�E\���m:��&��0�c�D��B�nG�t��^
��Atr�q�x�6w�|2��C2�����As���t`�� +JRVb�%�z1zt�a8��z,T)23�K}���MO�-_�!�Qb/�^�Z)R�W�矰�|����Z� "��:1�ꙛ׺�����M��Ȳ�Eיj�x�<~��};C�Ev#��� �>�BS�G�?�#,�L���U����}�-���|�����h�4��2{�u�6���������`����k�s��?��H��& [ya�8�|�c�f�l�������$��E��TF6�$����#�4��8�jw-�0*Vi�?5?�j1�e�O���*F7O�5�8��o�*�]h�h�2w���zY�_Wl�1*�sׅ;�"���a�nF��1�ݟ�z4!.b?[1�$���I�y�wjV�P�2n
Os�ȉ%|G���1X��Y��<>���y���nX�,pGъ:jme�/��`/�p�D`�������F��Ā۾xߠ�QU�����<�N�w��*`}�:\���9�`�$Y��=׀y�1:O��������|�\�OG��m.�JS��0�Ѹ�u�Y���9!+\/�uO�ܝG���,k��=$u�&�0��_¯����4�'�?<�,�@Zՙ�&�ʼEN/�\\�lxtM�E��V���+|��5BHD���$��\Ȍ����V�^��v6�E��V��N��`���uE8��C�'z'Օ�&����^�3�`�ș��4^:����΅��L���m���5��Io l�/V-(�M'�a//*�D�z�D8yTfr_;�s�����Դ\eac����*`3����H9�����V�F_{����,�PE�w�u�˞���]	���hG�R!,- M�)~(�B<Jn�kk$���]4C}��Ëj��;�Y����%��6fƟ��i5�Y�΍/X���ZDe���<A��F��m:����./
%$g���z�Ab>����%Q��q]�FH�+M�f�$|� 0��,��	��\K�?���Lf���u=,:g۪�q�\�?���^�۷_��K=Q�{qW���2OF��&��4�_Py�Ŵu\S�>X�A*:���Wke�0PNޭ׶6Kv��t�(kj$�b�(w��ٯ�{�_/V6��I��ڙ��ȧqѩ�9^Z��Ti-.9��lH�?2�_Z�񐁩?�����bT<́i{��G�Į7qA�A�WR�M�}��L�S�y���Q���	�l�>��D\���# ���HK�i<^���P�
�4������ݘC�a~��.ƒ�p�w>G3D�ik���	��:�#p@8��	u���b{��w��E�e�
sI�7���O%E���"�9���Xm2}��X�ށ�bo�N��6�E�O�����;��aƮ8h�!�(켧l�9SJF����8�I⹑�+4w��jd��`x&�����Щĥry���&w���� ��"Kk=���hfQ�L���03 !�u��H�oϓ�}pj�4���M��	�������o�[jC�2$��4�w�CZ�t2�,���9~R]��Э�|!]�T�f�1=��&�e�Asw�jQ�.C�콷n�Ym[�K4��>���9 ꃅ�:��ck�)0�˳�?����/�1��ߋ�)�Ч�ǭ�����茎������q�>����KJ{1S뮤�K��j�����ji�-�1x����D���1��f�D�{�lQ��� WD�f�zS[��y�^��w�����p��F�|�^�]��Ph*�^�bs:���A�OZq��?��L|�ѥ� ]AQg�1Q$�c�#��=}�Ӈʋّ��J��@K��s�|��f�F�R;=}�:;s�Ͱ��i��$��+�r]1�~��"3,�L1�ZAe�ﰞ��%\Sb=�:��P�v@0��o��f�uZ/��/��TA} 
%ҶǊ�
�e��ԕK�@ >[J�RǭW�,r�5�77+�7�'���	Ϗ.��[������M �-�����gI;�Ϸ.���w���Sb!{}��b���� $�`ڵ�ڜ�6�W6рs�zh���Uun5����K�SZC���|�4ߍ����^l;��a?s$� >��z��	1N��y�ݓ�R7��F��[p�[cG���<7�Ƀ��Z�c�<���5�(GRۖ���A���A�9�K�*�:岞Y=�ؼ�'̜ݧ����(��Z����K��Z�uM#rV̷�w8+KzD]��P:�n�[d����;�\g��cK�}W@��x%�6@�Y!l� ��_Ug����<5ȳ�׍C�D;�Y?�6�MS��U�_�{���� 6Q�ǲ\s�p]e�v7Q��ֵ�������~�{�t��!� ��z���B}P����z�?k[|��
�y���F�z��ŧ&�̻�ZWz��X�X���lX��%��e֫��9e���������h�����搚�ž�r7�Ý:��Pr��CM,� �yV�VPt�Ie�/��|ne�h�"�����ڮ\��4�z��OJ`I��f;f�Y���,��_Jؾr@�`ꃟ�-���4
�D e+=�_�{������)Ո;"�d���ҥ{���qі��3���2Z;/[+�+ӑR�i�42\�x�����'wo�'��"˕��Isb�(���	�Rk�	[��r���/<������5��,�C�EN�
d���=r�22T|62I�A+F�!zه�yd�����T`|�l�75���a�w�&*�xKVׯC:7��cڄ�H�z������w���]D�!cR;R+6����)��ʌ�ɞ�O��uO�ZW������%oܹ�%�`��>�0q�o���3"c8�70�� �ij3��{�I�.�cZ���d-���}��خg<����V�x:b롖��`hD��bD՟�MzԎEp7eN`�,b�.$<nq.�v ���l���P*���5#�\4㩝Yn s@�^z��,5�nU'��8�1�Qz�,��;���A�*�x&H�TUTͶv��?�ʳv:��}Ɩm$,�P�X����6� ��XN������S�{�>Gs�kg�:]��Jw�9$�o�_C��\
\�!(8����S�� iUX324���2���~	zm�����m�d�� 
��/b�t\��OPs#q���R��r��O]A_����E6�h`ϗ��ˢ��a2D�&:�;\���� p��:���f�.����2�|c�g��y������je�Ͷ���3�D=@��ɇ�����3�e�#n���D��x�p-�
�L>kq���g��-n��
n��"�:ԛ7(c�c)�̋ƙ o`����lr͆�m3�b@����D�^hL���y�-j|kzA��UN�E���/Ǉ�5�_T��<��ܟ�4����sV�R�/��zB}4��:m_M��T�O����\�J`M���wg�u5�~A��U�0����s���?�R]s�d����{��p!�/�$E_�c���{�E��C-d�����N�e�$ap	�5T��Q�r��P"g�ZA�4ç�0�Qڛ<��z�臐��)��k���]�����f���T�z�92�p��ub����
�/�+��G���׹�b.~������o閅!���<kN�>0]�sKU:u&_���sF��|)��T��L�sV�Kj@�J�_`!��Σ�����G�,�>F�
.�~I��|v�â~���O�ʜ�?������1��7�TV�*+�� �)hj��Y����?�>)a�E: ��ܛ�'�h~u��ˀ�)�o��T���AՇ�/�5{��p3� u���L)'�z��$�4�4���R]���Hۆ�X>})F�R��]oR��/�d��T�׏�zs��k~�'����L}]��Jq,�3�N$d|�л��a�������@�8p��
�������j�P����Y/Ә��9��V��EP�����r� �R��R�@��[CTD��N^E.��!���㕡�����pJ;��;[:ў~i;S
%���/i�4���t���(�yI�/b��r����E@�,�CbTK�IT{��Ɔ�'{pz��:���p���g�h�^�٩�y�*�������!���X�K�Wؐ�^W����K��!�����:ӟb�&�$����� ���a�⻌(�n���{F�s+�elW2��]��4��u�����Ұ��<�P�����  �Z٣Hs-������A���]�x�����J�Y���n��`���iQ[}�]*��z�7��2�Qp�ķ��=�q�t�Ht��9�/��v������(e�X
JA��P��fj�u�\j��/���g���H+AuT3dk/�L�t�4'u���������"��л��'g_}����M8)�pe�F5�����#ֱ:V;3�KGK?ٶO�g���9cs9���	�膎�3\ՕȮn�Թٍ��˶?�ȴ��g̲$�SA����-^`���j��U���@�����KԢ�g�p�q�w��h��ɿJx�_ہ�to�j�%�!H֐5���E����{�.�٥�f��^��T|� (�)��U����"FA�8i$��:�d�{%���f�P�("��2/����$����p�8�^��4m�v9R���檪��j�[_�~��Г�~ؾl�'�Z>f.463GӁy1)��o���p�ch�����?#�ō�#?G�w�=B�h��~S�UH.µ�T�Nj���u��^J*{crN��
#���=��&j�����	�T-��^	�~"S.|��?�S"�5)l5hsȻ��n�LV�"B�9�^���w��0�p@X�L����L�������S�x��w�ºY2v�<G��i�^ñ�H��(K��~G�d���a��W򽲺���Xֲ�ؤ�.P1տ'���Vuf�y�+��s>y(}ơɀ�I/O���e������承��Ѕz�}�U�`ܹ��{�����/�|ַ'�j�"���K�� �BI��
C�j�*>pf�P�9d����@�oOR��=��v%�s";@ٔua�4�_T�G�%d����iٳ��;;�$SK�2kwi���o6���^��s���_PT)��la��Dȥsd����}R�-++%�+ޘK�7�I�VnQϞ���>bP}&�5;�	9v�h�wO�d�$~��xg$� ��������I��*^=�Mw�v�T�ex�?�d�4rL�iǂ��I��?
�2G��#|�d���S$�ki�r�!�Bs��2�1J[#�O�/�'8hbx�|K%O�23K�����_U������(+^����Z�U��S�Hn�-Gl6�^<>�1��W5�}p�ރ��K������"�WhA������9C���0��/v�h��X
po�U�p-��j7a6��z�=����?!Xy��ivyV3c��P����H�L��.�)���[�Y������L�W:���h1��-t�e���O؏9k��lp�6I�g[�_R\�G5�ն&����Ż�9�Ӆ����t�ٶ� �V������7>b��%=Dܑ)g���븬�iޢqʓ��kӜ}��J�r��H��$���[��-+Ks�ތV#�o�����|#]���?q{��������E�r�,-�M�vv� r`_2���ƩQ+I$n\����4��{1=K�Ԃ���D��\�7�����(m��ܝ>X�7u�����^��.|�,���#x�v-�)���&x���8;�t�B�ɮ?�=s���:�`�qV����T�\}���V����VvG��BMO����}h�R'�-+}9n@�R�lY8��]	Vh�3#f�0����aż���vY�JJ@�C�
u�Q�p����֭��
��wS�[1�������b ޢđQ&ë��v͒zhjH�N�t^ִ�Қ�x�;"2�E�jP+Dg�4"lܪ�';pZԉ9/פ4���;�HE/� "8�oݭjf��1�cP0�l����-�3|5Wit��Aܟ1��\���y���P�Ѕ2����1�r{"X��Ľ��D�=ZҶ����&UD�nQ���;C�6"V��UY��ۓ�L���4y���_<����~�H��U��;s��6�@�*s[����l�����"�? ��rO]x�	�{�����.�s�E|�,x�f�M�K��Hzӹ�w��7����V�x@ic�f���$�4�2��-�=ۭp�6���@׹��V�g��?�-p?����q��ƚXMkrE��_kC����p␫�4:�˛W�P�݇�8��0(�w�P �����=���-rd�����=.����dpfr���toř@҅�(�l�~���-�X`��9�ࣾ�Q���G��3�}��-�S��W��EHu��u< ��6�-���m�Q��}��z�4p9XyP`�&S�w�b�2�e��^YQ��T5�����Ҿ�C�X(4D;�o���/��Wq{������:�x�?��d���t�ے+�L�9���=P��*�X�hmH�Zq��M���{�A��e�א�����\���R�p�<�48�M%O�aN��ļ$H\��&��ɟ�L��h�F:,F�a44��?Q�Wb�}/8��+�P�G_B���e�F������L�N�	����fc���������ל
N�g�/<�t����:he����Kǹh������bf�Y80�4��<Yu,.zJ�qy�q��H��~f���8v�ѓ~|I��#�6������<��+u�/�����)�=[G���,`0]�Є�U��XنS� U��3`�v6X��]��?�fk���L
<��z��t��E-+�7^��~�i�r�~��W~�3^U;Y�;��[0�s��8"�3c��Y��8�|T7����X.�E+4O����r���SK��Y�����_�й,=h��@�Ы�9�n�uP�21>�*�65+�6ׄW��e��K��Vx����� �W�+�m:�����[,c�g%4q{�l:�P��
ټ1�<����2�R��璫N|o"j�/H�7��x1�U��$ȉ4` �B�;^9uo�@6@�����__Q�m��"ʬh_�7��|	c-L��l���v}�*����i��j��^�0G~�\Dkm�O�\_m�q����jjR5�L!��5(C�{�Af�~��}FGerҒ�+�)t^�\�`E�XCһ Q����y�,ԣ/v����h�yǴ�Z�׹;�p���2�sv�^�������trԠ-�����<;��|�-�S�3g�#�E���y[İYć���۽_��r�9TSo��O�ׂ&zQZ��"�"ժ4�6�	�;�ރ�f!ìe+'�/��Y�#�[3�w��������qG��Lu�5�4$�!���,��~4��{�L�Ҋ�`
� kO5������aE 7���w��G���م�}]J�?k�Aƥ��\ԬN��3��!��JB�6�I��,a��!rDݍ
������Vm��(I*Ì�c����j�V�η��%�ΣC�0B��������o��.�n�*c�F����g2>MU��1��9z)�ڷ^��yT���"�vG]tS�Խ�|�#��'��{�"�~{K�S���l�����J�� L1ш
�T%���W�j��9�#��������%&��)(�f���{��ƅ��(
b~�@3�f�)d4����Tl�w9X�ຏb��H����ԓi|r�UgtGq�҂�ow�)���+�2i��[�����AMbʐ#�8V@��Aq�36��}H����Gx�,m¶jא�2����A�]���uv�0�Ո%����:5�F9�oų�����9�JG�R�+ۙr��/��e�� Xp���\��J���k��	��Q�a`<��䢹*�a���mM y܀���jGC���}�X� i�
��E��? b,V6��Tc`�X#:���O;��_�c��j�e����:!IuK�c�'�M,��\��,,0qǺ?� e$_��Tt¢�{;*����LG��~w�&�!oR��z�W�*r�+Tk���]�s.���OJ���!�_�΍TX�E
������j����+?���Q���P����/3-3mhY#�*�Pb�ڪGy)�����`|��y�\|3��V��Ɋ�ߨm��x�sz�P)���I/���<�3�W؟;RZ3Kz�}��J�@�`�R��_��V�I��P]6���a.4y?�� �G괍�;9xu/��g?M�����k�XWB���}�Mh��c���[a�ͥK��n�˗ҫU�����6���O~���{�,E�tٺ��z���V��M��I�P[�ֽ��1]������i��y-�p>���qYp���o+9ڻ]*i�oe�M<�����������Z%�Ə�R%[;Y��d~(S�ʊ��L$86�cߊ�	]�D�D�����r��/�u~q KE����!#��6p�u��C�xM,����X��~ְ�T����e9�3>-��Yi��ȷ}�1�m�f�pNu^�ߌ��6@��c��E�>��?D �ͳ~�a�Ѭ{��qN�ښ��yЍ�8��^=ew��m�����r}�^8�~��ʷ���g���U�vyl���z�×+,1ձ4.�k�y����n�4e4�hcWd|�Q]ͅ����2�S.��%�xy�rk�p!/�hk�H�ե:v���ݫ��/�����r]��yn1��ͺ;k���/A��.�n����H��>u�	����da�T�Tf.��A�D�l"7�0 nW�}w�ا"g3�W�h�5�YXC��;f@=bC��.�����%ғ#���p辨�Cgs�Jy�;ccZk>�ݹ���������0��Ϥ�� 9�r�:~=~���ș�۲�P�<�G��F.K�%l����;6*��X�n�<��ӼDq2�q�%��ma]���/N1�˸�����tFh��- 4���v	���n�h�ڡj�*@ J�iO�������y�uwFΣ�!=V�"�i����V�c�:9tT��3�fu Ze�s��o8����1rf@1����	���]�!������M2֚d�%O����ؽp%�������I���+���j>��A2~aǥ;k�d����s[]H�eB��S��2T��#��O���2��ʠ�%R���՛���06��e���ڼ	��gW�"4�A�)�L�>���GнD�_F�����m�~܄����\>ggE5R�b�g�׶|��,�Q��ó��[�6���'K2���;���dP�}���n���&�=����Ͽx*<��f�j���C���DW�kV&��&�������V#�Ŝ�Ƨ�ߓ�j�������?4�D�
%���i�:�H��ͱwI��̌��}��(��<86�qp�=��z�������yy�s����������Ih����؜�5Ts7��+�ag�5tg?�DN����z�:;��;�\��p���pg�G5NAA�[5�/c�Z�_10<�u������Y��7O�~�d�����1��e���A���kK�[�]�c����g.���B34�xa�3��j���!2b�����t޽EG��}w�L�z�׻]�#-�r)�����.k����r�ůN,�������;���>�-I^} S��5��x��9��ڴW:@sv
Ch�w}�b�D ����x�Ǎ��a��\�n^���	�Q)\r�cx���2DAǾ^����g{Gw8*�����Wsv,'�r:[��zw�����Р����t��� a��ƞ����?�[��V�Ӹ��S.$Qs�1�벍�U�UA"G_0��8��+Y���������xB���/Ϟ��+�ˍ��:��>w������Ċ�D��ٝ����˥|����6�K5|=��v��Y&e�����?o�J��͟��s��\�q�ፗ���X�R���n0V	��srr��~����/��( ��ttha�M)s���.�ݻ�)��s&%��)!$L���|�䮴�j�Z��3"n<R����$������E��`�f��t�����o�x쎛o��Z�'��>㶱�'��C�b`�������6/d�F�1�53m&A��y�L��k>S3�\�g��յqV��I�9}`&��_]�. CDz��e%�w~r(e��L����?��� Z����s�o�Pf���)&
����.�4E��������H{��v$��I�M��;�1{}3�����De��k5��F9�\h�e�r��H$�d�\V�C��صۤ�<��|g��Ե��ū��,���
�=)�����=L"��b~`�r���Eh;=!�������8'5sʕa�0�1.�%�_����d�H_ji�~�`qRs��ʚ�8���}	q�+uU|��W�����Ş��E��e-�E1�]-���#J���R�'�6o�/�����ŝ6^��K���$�_V7��P�ѣƈ�uО3���ԑlu��I|^��N��7X[���HR��!��t�2m�^�������F~��]Ж���g��~Z�M����5�����~" 5'V/w��ݟ1��\l;	I8� Ia������a�I��k]6ET?�lm>0�ҡ[%�|Ԉ��.�q�^[N��R��F5��U����H"E��<���Փt��O�]�f0���{�%���>���/{�u�0�Kq&(HƢ`�o#�!FX�L���tV���F�Z`��H������9~�hSb9o}Tv���8DA��진����:a���>*���>�E8R�����w �5}��l�U�P;+�1d�;-�wњ<#�'�t׺;vI16��4�F�y��.`���Ţ�����Y��h�7B���7��(Q�d�u}e��e��R�1�ˑ��Sn�f^���u�~}����^���le�Ϻ+�VR����ɣ��%�s�]i)�Ӧ�J0���d���or`� ��ӌ6�#��޶�pk�����cآzx?��K����*uG�{�^0L�F5=^#~�g����%�%���RO{�=�����6�g^�z���țg:zӮ4�|�'>�\���|#�@~��G���y����z���t�� ����+��U�ʾ����,�}_^hI��fAw*���d���L����^>Y������=�J����;{BJC�S��M������Vo��ˬ�k�"�#�$?6�c߈l.%Es�ю-�	�<����3Ō�i��OX�� �b̦�k�6m��΄�+كA��������yp�/�R�Č\�.u�+�������W�ޙ��7:/��3�������J��)�/�-���PP Z'W,ǫ)6Z�?!
�y��I����7XX71���1���_�,�j�ۺf�"뷓$	��=	6�s/�ow�^��Խ{%kV�93%�#�dA�QN���$.n{$��+��Y�X�BD����bؖ?6�X{'׌ٝ�@�8���Ɏ��GU% ��r���*���2Tִ��-���5��n����=��K��dϝp��[N-�	f,�YG�d����f\GyY�|��}Z����[�	�A��E~�a��m�O}����3�*����d]՜� ��;V��nɸ�IFe��C��݂\&� @�E5�}VE6{!M�'�����/v�40ޣy��[���E+�_�~P��E����L�}��1ڲ������Zڸ}ݍ��n���3 DZ�9^ƽ=k���VK��]��J�,f1Kđ�;��;��h�&��'��q��d ����9v�%���
�pj����?4G�~��#���������K�&H9P��y�,y�*��Kd��}�U)�z��7�2k%!Df���Wc�{�Y|���ͫ��G��F�b�]�����Ri�4g��]^�I	�j@��-3J���)FΙ�Y2�E�1�K;�M����:�Y�W涘�ؑmCO\;���zeu��X��?pLs�~�H��{�-{^T �s��z����j%# �&�;�����!��l78����L\b�B��B�M�g�_��J,[~Y=���̢U�S6p)K����K��_Ӷ�eX��O�ןii���-���7������&2}��K���Y.���p�$9�/��Ϯ%��E��qfC^��K���T�@�I|������_ ��y�C�rk��`X������Zե��L�k��y��HW���Bv��������fh^�ĥ�BRg�	�#ll�F;����w��֍i�F�7����^�
���jq�[��7��륙v*Q́<��ka�/ɐ�'r��=�p�l=k����*� /r��ŶÞ�,2�� ���e���U@��^�k����)̣ ���{G�|Um��]�
��
=�m��R�i8�����H���Y~��c
�H��.e�5o�$���f���*��0l��(�Y�_IH��,�i!�A��Ė�(ՀΣ�PV{>�uGe.t�.�p�e�� ��;J���$#lY������3 l����">˂�z�ێ��曟G&x�#I�N����I���G�N����#��D}3q�B���X��{/�G��VGb���ϛ�Q�u݂���w<;Av��
 ��z�V<3�� 8&j���^xV�Sf\�ڐ�����zJ6����;��+���� ��X�!^} J�;�4xy	[��Ks)�k��<��� #-`ׯ���3`�cvD��/ܗ�]~��*��X�8ſ�*aT�=6 �
�:gn�cDc*2�T������l�]Z�"�$�e����i���e����nBTnod�߀����: @����\�s���?�4�D�Lu�*�ML���v82�?��R�C;���O����Bj���hۿ��HK['�2�σBv;�m����W�A?P⒒��r>�a�k�?��9p
�6�UK���h�t�����TzM&�{a�/\_0�����%�����H�x��P�&��OM���Yne1�X��9��Ul2vCC|I.�r�n��^�7��4N6�Q
�Xo	`����m��@\Q�5�5[�U��j?�zc�"�[���V�A�Ǣ,Ⱥ^}��������L���1�.�o1[�K)~��°I���e>�9�F��Y�3���)= +u}�b�fW�cw?l�6_ ����/ӿ� �
"�]�?�R�v������	^�
��	�9�^4.�B�l���X�~;��\�N���x%������B�Q�b�m	�#�9�X��[D��֞��S�C]�6�[����}F��7�
^�~o�m��6���/�`�ce�%�oȳ*։����~�����Qp?JL�Ϗ�V�x'-r �W�xU�?^�~��D8Qp&`)'O��1}��ȷ6*r�J�����yB�P���ݎ��g*�d�4��\�����Ù���B���]F_}P��N�/.����6��
��K�f��j�
ܵ$��tzͲ����@J�fvX��Y��hYT�t_��Qu�� k�L���ӣ��	g<�JIBա���O�II�{tb�؞̜��[���4�Bo¿Z�'{*2&�A�ǐB5��P�z��ͭV�H^RakN*�I�F�<Z�CY�M��t��W�~�Onk~�|�~.���|n��Ni�6��5d�cu��v��|���VL;1	Q{��fz"H����\F�Q�P6�����Q��/��������u�?�9�L$\{�Aʢ�<$�\�=M��tk�Spd�0G���	�.����[�LՒ��8������Q˙;��?y�0�m�|��4��B�3��qgG���'����Ŷ�,�$Z̽)FYVf�/��dg�D�q8@�kn���KRB�T=�Ӟ�}���Qn|N���~��2F1b�)@�o���+��{2o�H��4Oka�)��ҷ�:!��ڄկL�b�@�8%�� ��}��+>��m�$Һ��S�H��p�Xw#�
h� ���o<���u,�`7�Ze�m���q�{��;]m>H���A4���~�0����BMy1���U95��knU�R�]L�O��������V�)��)����������̠b�"�_���-�_
U��I��P��EP��ʹ�er 	1��C��sv�����-Uk��Mk���d��ۙW�oק�[祀��Qd=���GbR@8�uZ�P�4���+�qV��Vv���lP�A&O���9}F�%j����'A|Q+�.�	�;Z�rDBc���F��SI[��I�r�^mL��^8���sw4��7�����(a���"יF��\��b�+W;�w�"���e-wF��3��0D��f�g9W�a]�y����9\uv�O����Z�Ք ����{�t+�A>�T ��J�46'��.X�[���12���g��DW�,q�Y�OI�qVh���:�������㎔ ����d_�;�'�v7�m�4����y�����M>�x|����~��������
��F`cr'M(�*+��ŷQ��!�K n���N�D�Ԣ.�'��������JA��T�G�$Aܞj(�� "�*����n�>�����l��-r`�����HGl���OƯw�6��{yG���ҋ����^B�����g����ۡ�3��h�7�R$8y�K�*K�il�����A�д�,����`�jM)@�|�K��z
��В���B�Q�������sk����n޽�k�3�
��Dep����cb��}]o��^����Y�x~5�a�ViIH�Z�\��^2��3{�t�>�fU[��^˱�b����{��a_��U�b����ʘ-�)�84��a4�����Sde��Lqw��S{=d?s=�ͳ���U��S��P]��k%�Au­�:\�ˬ;6R�l���I����.P�ة�L������cI����FF��'Ԗ������*�vܢ;P��3j�M��B��F ��I�mOq?���0�A߹WП3j�#QF�n���(ն�l�q�E���s]��!��<��6�I��$eU�l����D	�'�{win6�ao�H]o�X��]H���"#uN3���X`?6��
��9:�ڹ����1��(B��~��M�d�^�R��������%��B�d��2����3��@��Ȃ>�V݃JJ��v���8fV~���Gv"��'��O<�_8�P�ҫ9��;�u^H>�N��I+��ꂎ滬��3˱���V~	��p�h:%�|�����N?�2�5����鍊Ur.�]	͐>�I��3��j�y��s���{�3�/�V�����z���Em��m��H��o��B�)��s���KY��d>��"�d��u�����cS�(�0K�*|k�\����t*]�Kg�x�����7����7�4�v1�4Q	B�����H��|>x؂�)~���	.7�?��,�{��e��ކ7��]�u�PF�b����G۪uK9�S����)Q���ن\]g��O�2�;h ����ǘ���7�����v� ދ�])ǋ%v�
�]"Z�ΰx��f� ��� �g�Պ:-��rYa�E�,��>������'���j�I�~��Em�w��)��Ÿk
EC^���������F /Ȁ:&���h�r�CinŐ?� �����)��j
����SO�+�-�����'	=�� s����q����r�U�)�n	;��ƠH�
�a|2 Pa����-���AϬZ�N&܈[[��?�bTb�i*x�~\ga� T��Y/|�zc$��C��g����������������2tK�3l�W� W0�]pS�K(��T�!I�)�������Qs�l��<G����5b�d�`��yB;)�NM: �7}������^�6Syq.FGJB魌�%�?,����F�vT�F��0���=�a3���<Xqb��DR�� ����pl�q�ٱR�~�m�T[2-�l�)��D7[6���B�Op��v�"Vs.�6��ڽ�N<������^��K2�⋢�GJ{��e���@�pZג�
�-ʗ#�8����d��r���@q�]�}BgOq���!�r -�pu<��< ��z���#�N�.�ur�p���Z[�~a3�;3r�X��L��:W�U#��I[��ל�uW��7����{��;'���zN�闕�6s3~��WG��v���p��Wb��`�V籾ѣ�p�L��xx��` 6��A`L�/r��X�*���RJ�b��������)?=p�6�������gM�G�\MσS3����#l|[k�~���.z8 �?��-Q�'m��_	4>�/�s�Z� � ��u6n~ݱ�z����i�iq�0��{�t�lb(�ނ�E�&��;��Z�XkɌxuEV�h	e&<M,�CMm9[F	8�r�Ri��H�Vk�Xa� �YPj-(!+M_��S7�u%�@5�`��Yz�̕��=3�si26������g����d����u�b	��Reyu��7�+ZXV�Tu�фs�m!�f��0O]��7�L���������Cq��_��>���4�8*�3v�-ɮFE1+�/R���[ꐆ2�i�m�m(�
��ߑÞa���yc��&��o�K&C��-*:&1%��@�,���ʥCsݻ��q=
x:�نo��/�\�!�?�ĭ��H+N�KӃ�Rz� ����E�!��l����s�v�q��Z5�.ٴ�?s����F$��N�7�-�HM�p�T�*�^�����xp���.�/O9G[ڴ�XP���IIT��s���X����䱒u�f\	��o��أ�W'�2�S��H��v��f]�t�,7R��	x���E0�9��_��[������PK��;Q[F����n�<-g`���!,����U�w�����E���E3D�NmS�{S��[�P;%u$:::3Љ@��VV��J5���+=�]v���։�J~	��a���{�ݳ��g�d�b��P��dO�X�~�p�SP���#�&��LF�_���=ܣʑ?�Ԕ|�[�'�})%�_�V�KY����D�����{C5nm�+��X���	R��@���ݮ	~d�U^�s�?�>{K�v!��0����%����	��k�mlŤ������n{�g9?�$||��r�����/A��(�s\!��K����#c�v�P��Z��(o-{��V�5��*1�������!o�(�I�T������W�8�&=_c&P��)<u�J�ݍ����� �05	������$a��Uq��� y�Ι�c�g�M�
:=7;��6CgJ	�C ��U{�U����%]��W�D)`��>�|^�F��(�k� |m�(����:�<5mpa^m��ă�1�n��ۊ�R��bS�}0'W��fZ��{������:�����O��2�	���-i���=|&RL|�����k0r'桲^���{�b����|ANe�際��|��A��<q� ��.���1
x�t�-�v}6���6wУ}���=3{���%S�ly��  |��҃U�%�bߢ��%�7'*����umlA��~t�� ��	�-�R*w��ݤ��g�}�iv��u���7ze�������y<���ڀ���֚ٲ�&�^>��I4�чN-� ޑ����YI��ұ�5�hAe���T�����P5�>�e���j���3+�>Z��4��>���oQNO�$�bG���%�/j���ÿ��	Ö�QN��X?8������*�}tj]Tv�"��;L�Uf����/?\>u����C���%-f3����^���ove��`7���o����3z����E����h���E��}�&))��m�lREm�}Է�3wx�X2�Pf��7=Ϸk?d]�H�	���;#���Sb=�ռ���?�A@��Yd��^��JM�8��Ҁ�^TD|�s����1�� ߏ���M�۝؟���K���ހ��v��}��/.���Ư썯��b�qVU�����3�T����7�h"�깂Ȓm�V���WdHZ�0��;C���u���x�%64�o�'���m��Ύ�x$Y�����q؅q }���8-�F��$6����'�<�j�l��}"OK�EM���;��ڢe�����ռJR���5��9�&q{ռ��=�E�c�!�  ���Z�ZQw���A�n�7	X@	����9PK/�;��QȻm�0��K)\3����W���A|2�	�";��p��_g�	THS����_o� ⍢k�.t�eV}M�����n��}|��^X�OM%n���KdM2c���>��t�ީT�]L�g���r��5�|��zk��D�p��<��(f�N4Qi,b'Z���J����,����(;�Mhq��ȑ�$h+�0�G�'��k���["5�l:��`{R��ۯ��X��y�7�����S�P�c�I͉��-4�b���ƹ�ȉs2"�o�څ�y����
 ��[UBM~���wO�@{)͆άG���Tx�����xN
��������_���I�C��]�
�~=d��A�[m]����]Qh�������w��,�'����t�@�t���H�j#{�ٯ�k��[�ڒ �2�h"�e�a��PG�qD�l��(�����zN)c?�:��|�T;��H3;�R,T�(g3�w[{��?^\hU��ɒ�]���ݾ��Q �z���b7��F����|5���{� l���q������~�L]��<���.	�t�/L���gj��۹�jTt6��^f��,�_�x�M�_��wXO��vx��= ����;���w��P����aP���+��:0JۑC�}t�a��h�h���Wmվ��s��{�-�{�n/����c��6Va+��E>���3$-�C��>U��p��ܠ��0#!�c��o�4iq�2MBlO#a7j��D��ɋ��!
?P���U��ޓ'JX��%��NA�B�<���#u6ǧU-mSܪu�K��ǂ|�
6�?kt�������*鬒�}W�o��uxz�����2)g�5fi�*	 ?���fK5��E��Y=��k�Tg|�*̬�</��I@!�lzch��zE�)�M�v_T�4X�
�"C�}�D6��q�dBʹ��7D�{W~	B� q���G�E~�>/ľUk��}yƊ�xBQ
B�a���n}����s����}�l\P@�䟻\q@�خ9�ފ@!=�l��=�F2����Q/2�;����p����4]}�d��To��ο��r���yɧ)��7��,w�n���?�/n �.�k0��,@��i��kkqF��t�@\.v+AE~�
�F�:R�9,��0��~"�	8{��+��!�����_$�{�`]"�#�
��Pio�]��a�+��Gߑ�󍲍�E�>>��	xjo�Z��|�@@XU�P��Iׄ,0�����߽��d,�d��Z%(I���E���$�!�� �p��@�Ŷg=����Vi���H��mv�>�N�lE���_��X��?4(�����_���$��2����S��gǽ�4�:�d�X�ъ�7B�g��r8�(�	�}�GF(�e=�F�h���_�/�s���)m��"~Sz�|�$�<�?%2@<�����e�b,=��ae:��d�q���zY<7�����=|��WK�X��{��~�jSa�L6a/����a�N�Ժi���d\��^�'�����iJ���80�����}[�H�a3p���3fȮ���8c�8�7�},���'"u��V�d9�Z�o��^^{u.��^�ӖP��Q%��������6λSR�Kr�/��E��Q|��ْ:���g_/��^����?���3�5b�K"q��$���lU�7���w	`��k�wcǤ14���]���3�+1 r�t�xQƿ�q~Z�[P���?�K�ah��6`զ-���}�O�Ό����4"��UW:�!f�Z���z�j�&�wQu�r�Q	�ƣ���&.�%��,8��Й�_�&�e�|�ִk1=lμ@�x&/�_Os������8�T�BČ:��cn�{��\d�:M�	ʕ�uj��̅ v~&_N��g�����)"��QP�x<x!k9���<Q^�w��$22B�+Yeyj�E��n�~*�D�
��S�M�1�4ҷ�I3����U��Xɾ�c-^Z����������2���8���T�V��Im\.��S�m��!��}��!yO�(v-����z|��*F����T�{W�����H�_��
7�}�Z"�v��+�ry>�H����Ǚ��/Z؜vD.Kw�~��}kP"��� ����b���t��R���0��B�$�܌X�J�&\����]Ș��@�X��z���}��:1O�$a ��Û�����7K�-��[a+������nnIj�~����N;��xȱ�~�{p?�:w�a�����5�`_	ܙ~ܱ�}�J�����ј��df�4ѹ5d�mÌ��7t�0�;�謹�%�2l�YN;��|��J��N�T�u���!������s���/��������mw���iݗ�����b�a?!x�w��p:�r^j�3ߑ�'8�1:�e@���y��������a�s�_K���*̟����x]Y�F��#}�a�݇���]��צ�Ȯ#Yڝ�m\��&r�-ܿ8�e�m	��Y*�$��Y��-W*{�d�y	��_��2`��su���>�/}F�� 6�V5 G��ݛ �8�3�Bs�#v��	j ~Z�1xC&�?�������-K����V&��+''O�!4���b⪪�R�*?5��#FFF�R'�)����]V���[��\t�
����χ�v��	RT�Aܓ��ư�H}�L�:?X@��_�_���t ܊�����~�/S8�l�Fz-�{ߞW�P��3�F�ib����p�v��Þ��6��A�WE�<Ӽ�=��C��!�ã�Ͻ���|�����|�ɜ,�{5O�%T�j��5M�z4V,$��/,�.D��3�.$G�Z,ʣ�sg���)����n��H�p�%��������hF��p_���n�Ec�R�AJ`�HF3�`�Vt_]=2x̧�+�e�U�JZ�>�o����W`<��]� ��Eʿȓ�0�QvTECu~C-Qb�DE���v�@���9�<-��2��/���Xө?PJN6S_>�F���+}����TsՂJ��]�ꖏ�Ph��CJi�����v���Wd���"+�	-�GX
���ƦyQ�v�;9�]v�	��nr���b�Ž�C����Vt��W�$�gk�UR�Ap�>�;�K�[���{?���?Ò�n+���vQ93�����:�J���s�姶Ս���4��>��'����~�jȽ�	��Ʒ�9ʚ�����F��������g8�_��~GQ%�Nm!I l	N�B�D�Y����/h|l���e����۱�X��8�`��W��8z��]��PO�xo��A^�o;F���]��8o��{�M��r" ��
�^��j(i7ij�x��.ד,����Uj(�Ĺ��������3�P�y�_CV�5=|�YqKP���+�B�4����-�J��V~�] u�ȖAd�,q�C<��#`SWBD9~�`L?8Ǫ�V��%��'=LW�|�M@�M�꾴v�M�l�͛A2���|��][����(�f
�hLЀ�5���{6"�����1��F��t#��+n
�f���̓E���{[�`0�W9�ʌ] =��4�%�<���d�L����ƃ��2�ܹ6��<� R�e��x�B��[�4�a�E����o��j����:�h��%��枤$<��)��=�=���)�~;��O5*U	r��kwP4�$?��"m�'i]��.��������B�4_�hau�Ab6�a ���3(1Ќ�X&�Z�����w;a<z����H\� �6,Sk�m��φ竷��`�Ó��#���V�*�����yt����V��e��'�0P�\	�������F��u]m*��2R��
}ΐ{�z���t��UuB�Y/���!��5I4k	����
�-�Ɩ��J���/���d�N��yA��:68l��,��ǋvWԝ�a�-��K����������|�j�}��<X��R�H3���O?��-̲���Jޣ��xW��v�hy�k�K�o=�Շ9�}����)�*�1�&l�Ÿ�����"�a�|�X<&��%�G9���s�+ 6�-�E@��gaoZ��j0��/�����5��E�����)9�Hɖ�e��\j��V�9�� E���ۑ�ܽ�6n<�ê߂�70�V��ȶ�A�Wr�V.���%f����]�U��tV���/{�+�Sa\�7�VE����� �$��y��c����A�xL�v��q�yD��J�h@Ր�&]A�`�HeR�(��#��<��R��Yϗ��>����"H�Yֺ�/`�0/�QZ!!5-����jBO>��%w�ZD��K�(��r��dJ�}d'ڣ�f�pg�~E�o�o	H-�|ض�����=S�̦��B[,���u����k��g�>�G8��.t@�l���� �C|��i.=&�����������IW*����!O�U.���E^�)�G��2��߷2RcITy��f�`��)tΫ:�W0+[���zxV��)����廊=H�U�C.3J
��i����)m(�04����g { rY͉���ڂ�u'@v��)��ğ¿�I>>x�k��ڮ�N/*�k�+���n�YQ���i��� ���#h`�Ek����>���N�r�J��F��������b0�<y[��
H|���(ַ�D��
Uݗt�G]� �厪�7OBઞ��,��	��z
�K.�\B8��
��b^��|M�Hj=n���>FC��l�!D�!��#��0"��?��O1Qa^����|V솫����#�ă]��>�������J�"'�e�{` �#̇���"�S83S|�d7%�����kwP�L�1�Uyd姖�/�9���\�1�<;�H�ϋ2z�]��gx(=����Ί>A��!�9-.9�>�$khht�"�vd�-�W9�W�E�</�g���m5�w��c���SS(=�agof0�=�|��G�4l��z>��%: {�1ꖝe�G��T�P|��	~�/��
հ'F�h耈v� ����k���4��W[c�g�(eΎ��o��On>T�8�"�W��k6���V�/50-':�t��U��>�O�����M�y���?̟+�l��oO7�J��0�2:����SN_e����fx��	�kN�P K�w�0j\�-���2�O�Y��#�X�d����}�^��ЯIC;sʶ���E������)�� Ff\O�g|���,Ԯ��f��=����zqT>��W�����-�5/�ڴ/>-��cg�%dx��4+��J��e+���[^a!��4׭�����(���s�{�����Ty䥖
ڱ�h���"����2RLm˗�4�[�~M:��;˧JZ_�`�a�H͔e�:��>��F21�[ah:U�Hj�Čn���*����ۚ7w�Ha�6�YqY6K|(��CL��r1���r�9�$�`k8����i�ûMx�<��o�@L;sl�	�T�_v������=<'4��j�)Ty�����Ɋ�-��ydg:	�^����-?:�h�z���0ju =f���jf��7v����0~��5��t��XZl��t	kQ����F���w�ʷ�9����헢���^x��s�|
v�b�O�N@�N�Z�<�������f���?H�]!���ZZA���9v�����,�Gs��ƞ+��t��Q�>|�v��}�u�y�R�PJ_'1�l9Le����BWx)Br�~-v��6���im-9,@�������Ūs�ڼr���/O��>�{�{��x[��hxL�aw���_���ƽ��, ��㕄$��L���T�3\�YO���/9��ڗc�*%���������;)ԡ�!��K���q) ��Ln$�50ā�?���u(bԋFٰ8q�r(��B�����#4�Ǝ�U��Oz!��Q��'e���慣��a�������5��.�
T?�v|�t��S+(��Ī1H��T3���s<�ۏ���|QkU� �N�a+��c�M���^0��w��n�y?���N��m},ڲ+1�/�u�@��H��
)Ap݁#ӑ��l�<��ph��U��{
����R z�x���]{�'=���&�8�X\tW�V\;�X2x1����]d�d9���I%U�9��a�[�M����[�.B��_9����h7�
�����+����J�{�A�͆q\��(��k�_�U\c�$�/0@��ͬ�c�:q����7��ܢr�����4�z�a�P���?�]�ɳ����,�3�	�|=-4���q����V�� ֭��*����7p���74by�_�+����{r�}|+�:���H�������=�aU¡�[s]������ʂ�{y?�F�B��]�w��5P3R?ɷI5O�/%���jnuV� q�u��ݝ�b�.a�M�"9��_����֧>v]�#�?�X{A�|�E�����7��RJ"E��WC�-_�*B��F��K��������N04P�	y��d����}�u�ڿ��^Um�x�U�2Z���4�}��\�t�	���JT��>O� ��ܔ(�f�y�>b�U@Im.�!�+����b�����Ч������n(}L�z��]i�D��}��A���2��5�>�PQc"���
����/Qt1���	,�t4O:�6OG6?u��噸5c�'���3=�k(�P����i�~����K�i��$�k�Q��&_H(��>�1�/����w/ m�,�$���k�Pm�|�����T�;БJ��=�G�*C7���	Z[?��|[�g2���+����3Li���P��p��_���4-��|�Wq�r�� ��G��IQ��5�^n�є��5��Sd`��)���\��h��^r�$�0���q1�z(O��L}·�$7���6�0G��r�_o��3Q�=Z�󢈎v#�"���4M��A%���z��aJ�*-�u���ˉn0Rۗ�v��#�j���_6N9V2��H�8�ܟhK�.�G��Xq���?}�K�,�h��0?���4/R��c��p6��)m󏘔ЏkM��5KD������gE�EKþ4��y��ۮ��=b:7v���2�[��'֒Z" ���c���E[G��9n�=�;�}��nb��d��]�f�A�f�f���^�O��:�~6����a����P���	D��_L��_�H<�i;(
{o�U���{�vm�4׋]�?��veg�����	kkY�GWﲖݚ!�{�n=��YO�W���Se�׳�?����A��S�#�R+E���WA���C�5)��+��q�����[��>�us����ɚ�0�K[iqZV�i�"��E_饯�V���e��-+}�N蘯���mz�Ū�ܜ�s� ������D�}S�K�?5c~Ʋ#y~�G-W�q��Hv�j�&c2j�����`2�h51��I�#��&?��;Y�yH.f[��g�8�h���1���w=��'�n��Fpz���� f��[��G{�o�����]ܫ���7�_#�n��_������m�iTӥ��6ґ��]V���%���n�#/,I�CQ���t6��XN�织�0���������q��!'i����گ��PN��R��Nv��.�\�ş�q<K7�z�ͨ�\��Al��y��<:^�6욈G|u�S�4[�i����ȗ��<�������z쉙���[K���d9���9���ْ�p�J&��
��#�]�SS����g泸���&�i��_����^lEY���g���Tz� ����Q���	���ZC������L����I��N�.�m׹��<�I����)�tT���(r��W8���c��Q��Z���A[���lDS�<�& S��M*p�9�s�[�t!�:�6���5���Z����xJj;�����>� ;�l3���,Ola��:⹘QBٓ�oU����]P�}օ�j������qI<�\S]�3*)9+�΍�S��2�[Ss���A��"�1���Ʊ.�,�ԙP1��^���b�''�HsOFѬ\y ��ӵ:wZ~����.�Ӆ��Y���ad�����x��5�̟���|)�[�HaF̬d(&�'�Δ~�؝B/�C<���
��1X%&ى����s�Pjj��^�6�-������a��}���+�i����{FÜ����)gc�d�Yj�c�_驪�� b�JOI�ů�Xq�Ƽ�����~s�G�+-\��>u�>��v�(NPjO xW.5,�K�@a�5+��G�$�����>k����1�ջԚ���͋�c�{�������U�����Z�5�NꮴJ��:O�2���)�'<�iɡ���Ւ �U����a����~�.���y�`���Pg`ۯ�}�Z��v����5�B1%��Z�ym�q���s3ݓ1�I6/�����FI^��,u#�v㫋|Qn���;$�Ǣ;Tsa�e×��e��C�y����O�hL��h���Q�	�V�U��>ٛ:�9sug*;� ��T�bD�O	��e�-}���
ȅk�����Sj+���5�D~0�?UIU�����mo�y(�s��*	�94@�X�e������	�=$ �u�?���0Zf���6�>�YH	S�(�NJ�W���n��� ^���"8e$�`�p�j�|�n�d���+�_�v�f٣�G���A�C�ȗ>�s����:'*��1���t��T�ߟT>��T��WȼVY!TY��5��+Y!$d\{˾���Y�ko�����|���T��=��9�y���:��MK�����5�ڹ,�rGj�[VS�+ђCX`t��i�V�JZi��d�
�G��g��B<�{d�G�
R��UmU�D�v�]���??ml�5�X8�9�J���KU�No�=���1��K�ڴ���l�W�d
ͬ��Qe�P0��4��\h��h���B6�Y"��'�8�����r�V	�uG�������E��8>�p�a��l�����΋�����=83R/��4�c��Kg�~Ԟ
?���ct(w�:�+����x�Y*�����"���	�T_ث���Gk.���;S��RS�j��ͷ��ɴyB��_[����#�{��e�!��k��1f�9o��N2:��Ǝ���V���=�36�`WO���5�ӣLw^�A���0#�w_�䋦c������[7�����f-3�}&;z��� 漹���V_ ��%��}T�5��^�ug�	2��|�I�/(�| ��k�)4��П�ÿ�(Q���f)Z�40��v��]���i(�)�Ùd�q�ɻ�Q������E�+Ɉ|���x!�yR�w�5_���j��b��</r8"~	���2��Ɋ&|�O�9aُ~9oۓHN��F>�Qh+"���h�ph��_H����=��(�qs�G�Z�i<����t��$����䊝I������2�y8YeY7-�~����B����ڋ{N��?=�}dk���mu^�y
����ф��e,y�=Q0�y���*!��USF�����T1���A��I������i�j������Mb|x�RMH���l5x���*[�n<�&7�a�ug%��R��Si�'��������z�ŝ�F������`.RǼ��{-6��;W�Ō���F#�0ES���u���b��ퟣ�*�.�3\�\Ħ�=�PB���s�z"f�蝕�[���O�I�O��~=W֦Y��?W5O<��ru	8�H�#�P��?��8������(V�mv�c��׹0���\�{I=��� ���/ ���"�r�4͠�2�����;OD����0@(?��J���9��S�3l�G�Ms��%[ܟ�������g�5�~hp*ƺBU}Dɧl�0�4����tK��EY�z<��y�q�d�N��L+_�Se��fs��[=Ȕ���_03����R�'�eS�g't&!�t�al��H�ji�h�a�$oq����=�md��e<#c���D��B�I��ħ���P�}�h�1�"ן�]"?w�8���e������������9)E��K`z"�����#(:�J|�}#�Oׅ�Al��G�����I�K$�<t���j�I��7�Y:\��E��h�"%39�]#V������- �P��_�e%K���=�5e���2���P�Hi>�/���"=bi�*od�!��?��6'1o��kl�M�A�"��Z�LpB>om(���,�),��wN�.:�"�fa�]��w�`���nQH���m��$g�NӮuҢ�+_[=B�8�6�'<S5p]�KE%]��.U�LaH�ϤQRČ�'T8�W>چ~a�Җ�1Nǥ�"�֛����vt�8\qy++
2^"�]:N@��O[�pVz�<W�^w]�=�&�E̼;jzm��׻i
�����ؠ�񰠒��ɽ��n������b�X].M۵�^��>�+�N��:b��U�.![�8�:��|g��w)!�y�jr��H�a����|-5y��*O~�ݯ��[����n�K�(�����x�a��bP��dN�ɐ/�"mt�V�ޖ��
K����`��*S�������fk�#��1�{<H�'dT0�	d1o;��R�S~.�P.a	�D$Q�N�v����AT{t��~�vt0K������9y���gʼ�n͗�ev�w�8�uQ,�U����Le��I�bP���>e�����>�O�3�S[8��_�*r�ļ<�p����+��H�1j��t�jη�=���p��x���TjAQn���}���.7�����p�E�v��c���^�kI��t�Xu]nr�m�&�2tY
��SB	���<�qɾOr�w��?�c�J�2{��x���Fϥ��x�u�$�jv�-ŧ%��L %�t�N�r{4�1�L�t*���KX>����g ��ǲ�}��j;�K�CK�Ī���N���g �oYB���jZ-7)�2unF��1�zV��ݼ�Ƹ�N�ju"9��W�@^ᔶS��q�8��B�ȼ�5!�cJ�.߹�x�(Br(��ϋ�MI�b�hr���7@�E%����I�G@HK_�E�9���?s��X����-�7�4�0�d'Fh��k�(�j�����<���W ;�X��S�V� ��)�*tV#��dz2cɧkJ��4=��m��\PK��t$>��]{&�/|�C��dMA�d��V�x�>���ny��� ��i[����<"o_�G���w�0�cCNMTOK������oӷ�Z�O�S�׼$��v��$���S7U����ti�QKO(�� 5��]`P{,�
4���}{-�:�R��z��Cs�w�����ӣ����9=pK�Z�i���Ku[��;!�9h�-q��U��W[�r�ѽNSŎ�iP ��/�̸C��X�뾷���S�1�����,;��3ױ�Զ�s�FޝɍU�yt���Q�z����Z@J�&�ɬ祋Ǐa��x~�(j�~,����~�c�'���w;�"zޏž��juL��m���f������:yp��^�����Q���"��ږ��:��sJ�������	p��bp����@��>��V��Z+WS
�E�>�]����ϯp�$�m:�տ��U�Y.I��
H�89w��b��q���S�t�����"�qb�po{s�->��{i�8�+i������Ё̈�0��7�����L�-���i5��Ҫb܏���_2�ū��*2�ThѝJD�N.�N�>hJ낲Ҽ! "G���CGR�ZǤ��䢦LB@����!1�� �z2�ӭ��^@���;���X�����S:m櫶;p�b�Փ�{}y�I���P��F�p�����c������IWg��v3�e�F��? �y��&�޸OU~�y�=Җ��S�"�o��a�m����i&|�m��˝�J�_��]<����N)su��zc4����8�}�W�C���
�F�-ݽ�NG�7�m��j��K��A� �|��`Ϡʛ�3Iq��,�x<�0�1&V_�q�ܻ���=mc{X;�x���Y��φEY#8�w�sT�v�F���Si�0VS��t�M姼������	�����f� L8Ċߑ��|��Y�bb���2$W��/=�����2_v���`��$F�j]�s�N�p��ým��������P���H]�~ƽ�(�(���х���j��1I��>�J.�FIÆ`��8�����e
\��Ď��T͑<�htb�D��o���	i�JA�al�b/����&2��r�-!�����E�"�M�X��D�7�oW�ߡ��H#�-[�NN����1�n%ĉd�
�L`�X��8l�ȹ�>k{�����@-�:=�����I�5j��<��R�d��u"�]k>����#�w�f�ũ��v�υa�_�pl��G�u|���lcP�{� �-�2E"'���,����� ��U���=�6K�I��5�&$�GFR��DG����O$Y�꫖��~��WMv�?]�p�>h.8�E�l��%]	#�F�kg]�e^�E����q'i�y���p��j��:��U�t�(��c-�M�"��Z^4�0)�E-Y:�X��)o�I k�M����wj^>��'Ax��M	ʷݧ�S¿�k!4M+�����o٣�F|dc!�M�s��!�_L^f��k[���-���G�g{6:����&Ri��n����ΰ)`E���OCY�69����4z�P0ݳ�]�N]�h��҅8pI�J�iH�l۽]�Η�����\�ú7��T�v�Ƶl��#:��e��M������牯ٸG.m��{v.����zћ�!�1���
��a�y=#z���y��Q����],���ۼ:�:	�rK	�y��ڠJ�'��A�-m�;;+C�VF��K_r΀��`s��]�쾳oV6:t�+�1�+�E��/KΑ�->��t2.+m���v�;��:��w�)��T?0�y��W�^�Iu&�ʕP͸��s¦�?P��ꠘt��wɼ�����Č�F$�&E=4a��� J	�9��$�̭��u4R5�6�.}-����q��0Gu�9E��U�}���F��aҪ3��J�Zۛ�"���{�@�74T�0�Dl�9�qV]���/<�����Z�P�:�>��r�D'!�Q}�Z�x�Q�P�ꤠ�jf��eR[;ü�h6+3J6xj�7�}غS����A$�mT'�t�:M)|}p�N�,�G8�+A[�aL�����Fnв�+������wP2�5���1�a�x�G���r�\�Տ�vŻ�Z�ޢsj��L)���J1Q��N�B+gZK�h����B�*�%�w�\�j�4��Ntz`��t��;�։DIH���t�˗�G��.�ݿ�8Ig�h�\c���6��q[J��_�[��]�p!�?��|�T��#����Hr� .�w�#�#_xHA��7���T�p̬���5�
",�w���/��E�tV/~i_�%��C v��ne5���0�ʹ��:j`W���ޒK٩s�!�:g��dd?�`�T�5�9kQ�W�ʊ�Q-�� l%�S}��>�=��'����=�����G�(%�oex�K����!��:�U���������zH���yd_^�/\�(��{�M)^*@)��hw���?�I�sɘ(йy�kk�Q�m).eg�s^QV�l��@Ux�^��OaC~��֕�>s��o�n�T��T�%�y��qB��
��,�S���ۺ��vcN�_k����PT�	t��7���g`W���l���Dh�'��HI������_!��u�b�{0Y��}'��|_��O�J�����s%���N�eDh���ƫ�U2���Ϝ�!5+���\��3�9�է�P��e"����r�����}�$4V:�@�(k��漃�T��h�3�*;?=�_��j�G�Tpq��t�Z����2��'\��Cz�T+�4�>����!ɭ��7��Gv&,Z�2�c��[�
's_	��7���&"BK؈�J�����
~��We�މ�w~��a�L�^��G�L|����zGΏ��kx����`c��cؾ�+�i9;|���r?�`'����IF��A�k�>�fk�ʻO��Ə�G��DK4��r\��e<��(I��,���E4���,#�����p��X_ilG@V+$����� ��i���-nt��a[h��>C�Wv?����p9��0���f,u]tƆ�ә8�9뛘��ӊI�jO�a~q��e�#'��.�D��!g���!kO��n��s�0%�:9��!�r��G���wpӞ4>3nZAS�8�*�juS{!Ջ�0��f�^W�:��w���������t�9h_^\�iA�ۆ`��jSZ�7�݁ɂ���У�AB>��51,҉��sJ�����F]�<��t��q:q���W1ͨ�g��ө�
GB&`�H�!6 ��)�c�P�z[x)�ud|���!)ӗL�G���&��e���#��L��P�=i$?gnVz�k�g� �h�������@I��뿷yTr��ҍ������e�[r�N���1_B.1�-��D؜���6�鴎� ˵7��8��c�6�p{h���PdEevb)�c03�-���Ɇ�0����;��ҷ�z�{�#:�(�^�ud���7x��0����ΰ�f)	-�?b�e���2�A����lDXD��BjIǪ�=X^�e����ܩ��/^/OUC5c�ΕO:�Z}^�Antěa�a.i6(�<��ڙ|$K�}IB�(������=�/�ͯ5���U^T&��Pb�bq�'��F�$K����.�IC�9֌��#�1w'��۪�^��h�g�]���6��⛆QQ�3��9�u��4!��;�b�(}_L�dJ;��|;y8~���-�IД�XԖP�鐭���w��f�?�m+��!���7s�:�uC�m4��|��V�˯�?py@�S�q�_��?E#��W �s����M��P������O�2� �a�8u<������M �/Z~(#�9�!_OCo��������r�BSb����-��\ߡ.V�T�f��etQ>Q����J#Q����AX��%��c�!����(8�������'7:w��\��J1t��+�?L͢�z>�����	�"G��.��\w>F}��	�]l����=�S��o��~��p�e���	���/�J@x��T6��T�����7.G�G~v��j���g)�c���0P3_B������OZ�X�X�kL�bz*ͅ�����Y�:�5+JqDR�a�Ms�:�Z�(���+��.�m�|�r�e���梌~�)��u,���)=�!滅�[����P0BB�CT���0�@Iw�R�)�ٸo��z1^A�{ch!�Qy-ݚ�ɿ��t�W��	���Ȳ�k8��PM>n� ����n%��_�7'�C�yZ�v��a*��-c��GB���ES��[-5���'�5y|�n�e��C5�1*�C*e� ���	��`��PjJ�\�E������'�\��=�wԆЛ�!����C��Db������Fn�i�����ʣO�hm�K#)D�O;����cI��ME�Y�喖�����S"�u�:�ը��a��<9l	�4|���/�e�� .ް#H�X�����p��	oX�1Qg����Vz��`Qi�I��.K����L7�"��|g�Gi�g3({���p$�"�;؍��� ���x����O��;��K����:/Q��J�@����"�ϼP��Y���_�Ux��_�B�?�q��<�MB�}�o���{��Y��d�ԧ�p=�x�a�߆(��㐕���b]mW�gwAn(��Pohe羭�9EZ
��k�9���ޫ<��O�{��mE#���׼�PrH�&��g�V�K��dI�R=#��W�b?�5�&�(�GRZ��fYZ6��?��-ПWV���c�Tõ�0&�6ߏ�u�`-��A6�#%�� ʔe��i��ӻ��/�7�=���ŭ��3�G�~���Ȗu������#�w�I\��й��!������o|��;��:;���3��}��)�D�q������k��u�k^e����X�y���6����XW�뮇�>�$.@:�՘Řn�r�nR'�I�Z66���[j�'2��@�,�.���nHr�,>�|���B�$ v�	�%ï]�� b�N՘��`��T����Т�*ڢ�b�Q��y��р�xS�.���H�PB��ɓu[,�nנ���~�I��'#�="s�g�n��Ѱk� �:��Ӡ,�"���!��JJ�3Լ��,��/'�<�\�,���\�H����m��a�'�_�F�%s���
�
�A�D��n7�X��Q0��6��2J�^����|x
�ĸ�� a��y	$��ee.���RB��������4tp��گ�ash"!��}�	��$C<�g�v@��9&�:��+�9�D�o��}��/��c�$�Zw�8���?����Y�L�����L���tR�@���	pT��K�ߊו�gw6�w!X����@
�Bs
��OK��g$�r�<Ri�T.Rq :~�91��5$�U�i���QHW�m�4n��L���w�h���g �_= *���z�Jc��ԛ�N�C��=���|���< �uC0�d��`����M�F3x,��y��VѳE��ݜ� ֩8�"&��8�3���9֗�R�茅�2�3�jTS��/�N�ݯ�\��6�#�趔T�`�@p��=�$T��[��>����_:����pv����13�%:�2U�'c<'�~�ëݧ���pmB��� �=*�_�e4��L���ImP�bµ����7!�
�O ���e�3��dD�cV�yU`�������[G�<�*x�"fޱo��i���м ��U�Щ^��R���`�����l'�V��H������}�q���L��k1n�9'�>g��9�k�L[��`"B���C�e?N8�YR^H��>f�G̲�t��+��"-�s^�Es_:��1��ꎿ�{v�8�}�p¦�+`��WnX@��\�����Hi#9%8WWG���x
R��3�8�i�ug���ܜ���T�I��3�����/�Y#�����R�!�|�M���~��&�3��Kv��	��\t�t2��I�����t��d�H#L�¾��m�,== Af<!P������~���5d#ߤOF*.�Ó�5�	��wG��n73Zn��D�:���Ti8K��Lj�$-<H"!Ѧ������n�V�L/�fr��O�6�OE�!���|�M�j�B���@־yy� P7A��a4���[m?h�Jȋ�:f3�C��#,L������WP�P AR��<��s���ⅇ���/m�=O_�F���gY2�����pR01���ԯ-x�̿�s���~�-ĸ|��]Ȫڻ,D�!8���=�'�z�%j��r~�kR�[���%~�i�$���W�A�x
�w���$a�ŵbt�"�Z��N�������+�rXnV�|	�v� ���S��e����嗍K�Q=V�yr&���?��!�� y(�����J��ˋ�'�������U��<��1�
����>�R&���r�����7�O&����������(+��̈�Г�}fr����'ﶺ����g�v��<��"
~�h$F�:p��+�MԌu��R��%Ni2,_�"�_��G�#g�D?��P�����"E	��cZ�P��$�7C⼬�15���/_5���J�����B�=,�ѧ���_�؊A;��B��2[�`��;����]٥+�
�o?4��5�c����Pf2�I�_����4�b��N<����$��K\�ډ��a�5��~U�4�:0>��Y8�������kښ��)�,>6VK`���r��଼�� �e��15���(VH�s���I��TɈ�����E��ݶn�#�.�-7�c͔Y�n��� Q���?:��T!IC�z?[��a�b�\�z�/]�-V*4�؁؊��h �j�3/L������_�4L3�Si똎q�rIP�λ����Ó��\q.[�1s��l�Ӽ��Sd���ۻ4%�\�T�t�+ߍt8d�=���w'�h8�x�(���"@�O*7N����;�2L��B=gH�D�?�m�8���e��(�jtt^GC���Z��I!�v����mS46��O�
�������&��
9�j[���$�w��5��!��h5�� ��
Z^�al��.c����A� ��ˏ�u����V��r_�> �lԨ�MY��Q����*�C�}�Brz���1DG��� ��Hu�Bw��> [��=^.*��5+~�#u�&�ng�.��2P\�j_�f�t�zb�$�q�ON�����>#��c�]�Y��@��5 ��.ARtV; �s���2髋�/ۡZ߇�����Zbo��?���>ۼ���l�A��~ְv-���)��T2 z��v%XC�JpT���jE���@�$�M�x�Hէ����1����<x��P�f�zk|���`���0
@�au��e����ْ}O�hw%�Q�35�w��d/VC%��
MӶ�VpXI��T�c<O_9_�D��	�z��&�[;���a�Bxq�:}�Z+{���Y�W~���Gw�M8(�뾥�<NC�Y����<Q�)��JB�=8� �L�)���	D�	=���-ޭ�����&�V�S�P��+��q��H��A�2������?{�e$,��F��!���e�(��}�o���{���ॕ�~>��v �9�/�v��o4�kΟ�s���G4w�/Gd�s����_Lvyh	�}w���1�M1N�Uߣ��ⵛ���Dd�N����:IE��t����܃��ʵ
���~
��C�^Ay~�[�?G�����g��#Z�Ql�<s�E?d!��>�Fk�s`
"G�S����5���3�T�Z��7&y'��x� �e��{	x�Rl�[��<�h|4i����0�W��<�x��P���iiIk�S�pߜ�e�Wyb��`���L?�b���Y�a9�K�����`
$zMr�U�7X�4��0K{s�5Wl	��n��XD֡�'|��v�ߵ�۠3�
�B$��>	���.^gk"���H��b���'�<!��'lQSk�=�Ջ;��	 Z��	~Ά�x?b
��8���J���R�;�Q�0^A����[z�{��݉�g�V��QY�e*����y_�l�.G�bF�\��Si7Y�[���&	��J�����^��6Ɖ�ot|Д��V�G�;�Xjb���#�~I�}ٕR4��I��1ѩAF��N��W��B
�k_0@�T�dKQA�� ��w�~Xs�s��3�xg�I��a�*��m9U�׽�`�����V�ʝ	�*9`� ��� 2��*�0xN� �u>7��U�j91�Y>�D,��i9�����ݏBU��X�3�ʃ� ��I�-��J.��"Q�pbl��mVBn;��TlZ��2ej�Ѐ�;�/�X؅p
����͐�_ɡp���ʱ�R��Dh�� G�<�,)8�=S�����J �تZ�j����X�SԸ����z���\���|fL�����:܁�qH̑�{�[=[,��cA ��]����2.W�\�j��q�-$=����"� ���Ŭ�V�W��:��uà'�ۗy��o}�g�pȧ��}ͰZi� K|���A����;�3U�}�/'r�냁�fU��b�gT�i� �B���*@V���L�ӆ�|�/N:gy��ˇ� Y�#�$�Q���/I��+
���wz�:�sR�6�o���<���	�dt�6�}9�]#�d��	��o����-K �22}�Ӟ�e_��eLl��Né��2B `^|�ړ6�V�(�c��-�4��t6�~l�_kqP9���3� �RKy�bF�1��Ԯ����w0Q�>]J�}�HQ�����>uS{� SF�ܩ�<A+z��o?��E5����r��DX|�������9<}����F4�mh+�xyU�<��>]���L�o���|T���;\���x�>9?1�>$$Ç�{y�������_yc���`�.������x1����pH�WMZtQ@��-�Ñ��iY1-�}Ag��U�@�n$���I�K��=��(U��/�*��0����E�߻�h��ޕ�E���������+9I榨��le H[Cb�^"@�AU��v�/�8B��B��;�f�/9�CA,�z���=��"E�w�2��YҼ.:�sY&�e��13���⃱ſ���Mj�Po;�}elgrM����`h�������J��9},�n3"�����=���W����ʨ1��7�M���ѷD4�t����w�r�X���Xl���<Ts��^2�� f}􏿄��R������~ ���ԥ��2Øi?Q��U@8���l�Y�o�����¥�蓼$��%V ��z�  � ��zY~�nGU�z��W)��$3��;-`�U��Oe���w_�)��ȓ)�~Ѕӗ3'�%dg�����V���Q��z=�&�,�\�ֶ6��KӇ@��I8����Z��;Zd@b��y�4�dνl��ɴ�ه�4HCM��=��4 ظ߮�K~]q�9P]z �L�xm)��-�-$��{�=�̊W<]ꖮP��'�֤N�
 �eh���iqW6����4q`-�����H�or��@N岥��?yJ�T��HLo�Dш�,d��(�G���F �Mom{���)�~��E��oԏo{>�tɔe�)4�y<�h{�n��${�B �	P�\�Yz6&�BB�����0��	�=�i�Y�^Z�^����}c}����t������+�{_�,F��o`D�'�� �W�]U�j΂�������_�Φ�go�V)5�M�N�|�"�ad�&Q�(��'w�GwhI2A�.��8f ^�J����|,�{W��w��J�D��zq씂��n�؈?9�x��� ��w|��P@��ޘ���}�px���c"s�L���e��Vi�����o[,&�������U?��'�Ȏ�@?#�w�iQ�t��Jz�A&�8�5�՝�m�w�<o���w�f�P�����n���R�U�7�KA����;?Ȣ� ����Zн;	��}W%��������ؠ*a�ѧ+�����x�i|� ����p�j^�2��kKZ����Uc<0a�L�p��TpA��_�X��=��rи��ć	���9$$ak5M�v��GS	��k�%T˶��?Z�n�`a��[�u����Jv��� -g���%'|U��u������Y��^�ߴ]�|�2?\�7Ѓʘ�3�$�7�����9a� (��6�S�y��Py����	0)�Ou|'@h�����_��6�2�F��9>�_<��i�Z�Y�u%�?�2π
^e�J,���' �N��om�n���N�^�F<{!�"q����d=�NwߞOm]d:^1�P�ޠF{�d߂�9�aMR�?��C�#�zv����3��iO�ӥ��89ٽ8J�!Uw�,�� ��C�2uk��y��>�qC�7��G4UUbK`�Yw��$�PL�i�6[2�}:��tg��H牙jcv^���+^�ʐ��������]\�x���{�mO�^Kb�?��)~5���p���k�L%��m�[@ӴGDG�vv�t[}ʘ�����*��<\o ������wu?n���3�����|����H�3��/є"�:�ЏpJ}%B��U���gE���A�-Q%�BF2j<sX�����SIL����\�C������ꅔu���K�r(���3{S�ka��[
h�=�ۼl�;�6[S�{��w�[�0�j ����!>���|x��ǅ�,aB�f.��� q�����o�������f�3�yp"�����>� ����Z&_�<}�纳�壄�
��i<e٤��X������k�s W��3�_��-G7�aM2�t���T��/҉i3�OZk<���Ѳ���<�`3�����'n�5��
v��Z�����ۄH�_�X�? �=-8zg�v�hqo=�B[,�~�M�\},��z����s ��}��C��Lp�7N9��S�]�V hO�<V�1�!����!3?�zD�,�VR�=�wcN5�SQ�P�'���p��|�;�/��t�q���L$�_�ks�^����T��� �t���'t���..�W�G�@dܞ,��6i�J����lm���A�����q��ɀT�id�e���G"�[����8�u3Ev@��K��T��6[�)�<s�6�JT<�A�p��| lր�8��LeM��qT��#�(�$�4�E�%=�� ~	i|9���v��Cv�p�jb��tjP�&acJ��D�"�`,��b�I٫���Q!:ݢ����
���<��4 ��w:�?QR R�Γ��'b���q����Z�L�U��)�3�N�-k��̓��Z���[�
�����O����9:@��6����_0@vp��\'9�Ѡi��7�=���+^�m>�h��2qx�����W�xY�E���C,��%+1��V].3ѣtě7B�BG�&w���?E��!�v������זl��&��U�
π�5�'��~��� ��F��僘�@c/���JY>�)� ���@�uK�����<��(�)j7
끨Q7��T9��B*Ap��&�9'\�YZ���3�c<#P[�O���o!��P�m�~�>�O3�����h+f�P�CѦ<������� u!�:եj���>�M� E��n>E{��(�ОE���X�I�UYَ
R��d�Jjٮ����a��+v����<t�	��� ����]�z���zbI�F �H����ˊ�9K.���V�Ե�[t��9�({h�����(M�ō�X9���r("�mǻx����n��{���$��Sό��O �Ώ�@m���MHO��2%:��!	֗Q!&���1��7Z�F/!/d���P�kOz�SB�|͡x�I a�g�KE���I��o�셇�b�i\�Ep>]:x��V�t��ay����(�}�~s�ȱ�鏇���{h=�'�,net�'dZ�4s�"����n��T��/h�Z�j~�rD���H���a�[�)W���s�[��0:���4rb�ʳ"x��aQ���@�Ĝ�tMAf���ă�W\R�������J9��ap5i��fd$=q|G���ˡ�	�~bpr@��wm���M�K2�6۞ylI[:�vk�^(�n��z��mC���r���-�T�e~ӕF�K{�k��r�`e�=���������t](���(K��P7%������S*���No�"$e M�ˣR����u����F��f�<�\��v��8��L���>! �<ȥ�|�f~"!��a85�w�m��7x�^��囝��G'.�ȧE�<.�P�z�&����SyS���z�CX-i��Y�*�A˾'Pf�Gy@�>���wh�^�3��f,��f����V&�U�U	�u��v�b��[I���ǜ��p��p%�����7%���!`f�@�z��㐏�Q�UG忲��$�}?�݉��8�}�kb0���'��@���*��(	}�/7���U8I#LX��hC����k�~��\}��'���|�Z�6������;O��κ��MivޝS��|qq��c6�\�G"o|`-�[$?��Ju��2+,�G����[j�2�?����*Yu�)�����k��e"�OzU�#��yJ��bh��v�T���x���H��oi�fOQ��^������h����7L,����͈���[?δ#J��ֵXn<��l�0�;[$������'�)�ߟ�38R!�ۮ�^J��J��5q�d��~<�
�ʈ���� HxSLY���cl� er�3AY9yE3}��	�b�2����D/����5"�Q�7<��j:UmwM���9ڵ:&>�!>���J�ˮ��-ޘ�o9U�J}G7o�:F�B2�=�Q}z-�y^fO��Sx��ӷ�V̋����ķ;r{�����sz=�V.A$�-I99Y�A�o��d+t)�D�B���!ql&��l�2���>)�4~��e�.ߧ��<'�2�@���~@��ՋR)�J%_�m���zT�4p�{�Na
�g�mh�,o �\X6�1V�����G�,B��_U6FO|��-�8_w�9���.�5�5���u����z����v��;��������h���D��/�=�kVb)�^�ߪ�y�,���P�|��ⱱ`L����O`f���;-���53��~͙ަ�1_'��L�\z�٘r��3�?�_��m���������j�c�����h�!.S٨=1�q�H�~v��������=�46�U�V�}̽t;�qc���s�X������_��O��O��Or�o�B(I��i��sXΟ1(u��+`�;Ň1A�琶W�LVzB��t+D6r���ɇ�Ҝ��;�*�aw&����`J��NJ^�б�
�1�dG�v���13��]�ݭ;���!���e��7p�NB	x+$�F�[��˄r��M;��j7K��ϋ��@nM�S���i���JgKL��L�\�G�t4/?��I���:~٥��gN&h�ڣ�a���#�;a!n)x�I�ו[���K�<��'F8 <s�΂��G:"���jY�3Fܬ��/�J��O�*�J�!AJ��i���w��r��f�ݩ�	��[�R��>�|��qﵶ̳�&`��ZnM(��.j;%��=Ҁ�1 ?��n7g�
��˘؛ԩ�����%'D1�����}�����D���Yf����-Zn�U����v����+DQ��w�y�"�"z��<�L�oJ���qZ|�75�;r����k�+�����T����V��[�o<Z��ɫ)N�1S4��G��E�c2���������E�N��+Vh2�s�TH�\k�����5ؐyq��U�?Q�:�c!��O��~�z����Q��82��^�
�пSBW׹���n��g(Kb��:>�#�����6�Z(�O�mk���\IV�5m��KO�"p��PɌ|��>��7Ύ�ɚոHh$ҏ�I�\�4t�e�թ܋�ecIʧl3�vs䘭�-ҏ����N)S�q���C�S|�ʢ����5�l2e ��� �	���f�r�,�����YG��<5�,�:uk�R�V���*���y�0`9�ٖ|56�<F�� �A������*�&����^�]?x�͚��s�b�7��O�Q�
�E���{�������m���I�!t-@�����ˑ�E�.��n��h���%�����H����9��r��//8Zz�TYr��V~��?��_�� �*�uȬ'JI�)7b�衮 q�������e�tO܁��oA�y���_�V����[�����|�8� ��Y��#I[i�28�K��<�����#2@94ܾ�1��d�}�^*'y�Z�TH������,�1�����~7���A^^�
�E��_y�	��Gc"��;�����Su&0�Gl��I�7�=����&�Q/�����"�}��޼.*�����BIB�a��97�����r��`1/��g
_z�Qx�4@�g��搵�H�!�R�kg>�3��lOD��x ��v���WP���I(�����jya0���ฉ��B/i��.T���4�G߿VT:P�*�<�R�R,̫�|�Dsؔ�����:�aK��M������+F��`�+��Y�H����E�A�z����Y�'����f�b�Z��*Bˑaռ�ʪ�?,~W���mK��S���#��;��bbh���( ����9��l�h���/k6�}��#�'S�G6�n�֡��zA���P[�}�1���g�����Y�4>�nQq�|u���ܫ����{1|��-����:��Q�@Qw�� "(�]�J���R�%(�-"Ұtw�H,(�H�t����������>�w�u�qv���s>q��]� u؄�M��Bw�m���Y<k��W����3H^K�?���p�
��G��ꫩ�VW�%1̢$I�����mC�����~���PD#�4�Z<��l��5_M}q��5vM/?�y����Ym+���Ӻh�&C�z5�-b��V�=��L�񰅭A�* D��{�􌔌�c�y���*y:��hȅ�uaI�tX�8�1��^�|(�Dԓ
�K^D�{��J+��U?��>��-��A���o��c2�qq]^-x�o��Y@{��rR(V�>�R�0nKj~W��pu�[ma*�W���2����Ų`8�5���!��?��l���[����/��O����� x�T���A��h�ϗ��� �B<3�c�y��s����;��E��r�ҫ��3O�~T��Nj�E��hJ��L'��W�>48-�GB�y~s�����o�S ��E6]�.��nk����w�_  ��W{����I�<�g�D���bܡ�h6�*���G�>�˱~�M��ydg�iʭ;�¡Κ�g���A� ؊g1t��V����(�g����dS��4G���l@�4��/yEmd�^@��]T�* ����+�fm�i��K�u��Dfg��&v�'oE�D]FQ�l:��m�(
"X�g}��Z~k���FD�ħ��P̚�l��&���3��4���t�d�D��8����2~�y6�C6�Nfi.�7c��� i�8�СE��l�������|���/��� @��"4~V���/�_����:�:���2��$6� E���g@�lq@PA���\��j�ʮ��1��xƏB"+��[!�@�S��Tۖ傍hw�:)˗4�5!�C3��FМ�*v���_�����N�-����Oo����k�'|�
��nŐ'q�A��+����8����n(&��fϘ����e� ��ۍ,� ���ac�"�s��9
�<�{��In��>9�	"����"��Mt��D��	��r[#�����ڂ$��դ��������b�P��AK�V	��i�q��`/Ɛ�2���.z�����������Y�Z��\2;ƥv{��ܺ+4��L�Q~M7KȩK�f-�~��&�	t�o|�%����`��E'� (C�٪�LJ��gy��pq�7��O�ǿⴿF(����4��?+�Uգ=~���֣$a�� �n���@P©ϒ����O����9�e��gˉi�z
�U|�mھ�h��eй�dN�E+�������Z. ��秅�ƸČP�D�q�il=���Z��v�a��PG�!8�32ܟ��A�	'j�K�|�˭��ϳ���I����/[����8K8˳�ᘘ<)�V593N궷�a����q�}}���+�o-m����`�ot#l�b��YgP胋��p�0��]�+�$,H���J�f֤�qH ���������GL���$�:"�0�}���C���?��I����5�[��m��" ɶ�6�Z�>p�D*�aqJ?|vȒ�ߵK�pt�݆��
�E�5x�E'��R^�9<c߃B���'�.�7낔�f�% ���C����̇�����7�dr�����Znt�	�T��a�Y�F>��E�p��vǎ�_m�W	���^i����	��\��f\U���tJG&f��"������J*>�9x��\��nRQ���k��<��U�����/e�*�/����oUޤ�hŧ�E]}��FT �0=;�\jE�o��'��7�-������V�e8���X�"� H��7o�y��}'�65�hq@Ő�Į�A�|o�R��E�p3�Q����X���r} ��{��������B�Ъ`�c��{_ʖs��vf�ټ_�xV�s'�� O��?�����;������+��_�x=���-�;-�&�O�ƨ�!BD�qnYP�w��T[7U+�5��=+ؽ���n
�5vu�ۢn!z2p+���:���]�O��������(9f�4�E<�W,�.d�>ϫ�)K�5x̭�Ƴz�R��Q&�3C�%ǌxS8K��#-&��u\J&�wu����ͳM��	��*�ć��=A��bI��o˅�6�!6`�:�<�~!�/�?�nS^�q�z��8nN�TB�)G�kL��2i����"�t�Γ")l<�H��cV׽�H�L�z)g����6)������$͌O�6��z�3R#"�"��9�y��wg��lP�dpֱb�����#�8p��)�c|Z�Lփ��P����D�@�4�Y�ѸͰ��{ZW��t5��Y���i���(UȌܗL$�'%��[��Q����9�����(���1[7��mPo-�N�$,����|��)�v7*$x.�����I?��3���_��䨗 2=^<m׿+��	~ʹy��F�,� ���ӧ�x�wA��`��:
��t��"�!�����[��-@~fA�Og�9虂Sg�fN�T*�tC��;%D%P��b=vg��z`�'A�uLnaY�
W�1�#�*�~ȫ*��k�h�f���6-ȴ62Xh����5��G����	֜u?�ʽ��? �)<30sn/�b�)!j(���u�׵^�LI��5��>?�8�q�K(�a9���Pm����Vg)���c�Ą���a��&E���~;z��L��p�Υ�%f���â�6[�c���8�����h*@��+
�Wiu�P	Iɇ��ݨ�^���$�݄��z�?�,٪B��6���X_�0r�6�Gy�k	��!F���G���Y��ر���5����Y����V+/�XÙl�V).L��h�����GHL�f> 2��r����@DK��i�����&LPS9ţ�������$��8�sI\�12e��p6I�����e!'������?�]��#;�?�E�2f;?��.��}:W�������-��DS���i�/��X�ƹ�N��h1��H>;3=�,6�FCl�z&�wxa8��ӌ@ek��<>ٍP�<���ۧ�4s/!�Y��|���%�.sfd��n�{3��>�)�'n��V�Nkqt����D�@��2hk��� YG�P:0�8(OiW���t>%�{��+JcE��@}������@7��H/
ݕ��+g��/`�%��ė��ex�C�J��� \	ܱ���"�l�Uc��zk�Y�b4(�W�:�;���^j�K���G��:@�Y���4�=��wK��;;e;kS��_i���ȴ���z�Gx�����tw��G�^t����Ond{�љ�W�A���益�ln��ɛ8�h3{?��Gu��Z�7Qע^xz|`X/�ƪW��oج0�����r�	�+�@����ʦ�B �3S��M�|̻�)�@�z��V��l6���=p�
�UC�@���z6��f��s�&p{�Z0�����5t��}�o��J^���\O�s�r���&Չ`�
1��M�a��I���K8��-����,.��_�������y3�+
�o����'b�a,�����T3Gq�w]�D��b"��*`��\)����?�yy���Wd�����
^J�Ӽ��q��/���J�3��$��y�����V��Ё0���_�N������We����/E�\�v3-�*�@�p��W��	�q�*��� 
-(f���v�z���LO�� �Weuw*�4����;E�@F1�:���Ŋ��!z�F����j$��sXk�qyA»��xɘ��S�)[���t�4�fu��?ɂ�C����cv.�{�m�K�4���`�S'`��"�IłZ�_R���*����-�Q�eb��(�?Q���k����SR�Uo.�P�����h�f��Q
�R�����L/����|m�a?�P�a�o�o'�����`�t��l�s��6��0��A�nQ�ł�K�+��B�o
�R� .FT�U��_�������~p�2�^D��G�7�� nM׫��\kʙ�u�v�V��=,y�L4Q��c�P��^e>/�/Џ�1rTC��^��$.��7�B��&DzYbk�́�Ke�s���r�ϡ��1֮88�^����Z�0�/����9ب�:�f"1��C;�@Y��d�B�}�k�?�9��������;��D&�Es�#�윂��U%6���!|��W�J��Ex_�ߵV���W�JMp�U����ݡ��<�5)�]I��NB��Ꟊ&�/6�|�x�"��R(��66d	�i�ǔ�y(N�.�����mI<�� ]�l�Y��T���
�^���]&�!o�^�H�1x��;H��&3��0�D,G��:ug4�q�
�$rM����#��{�0H� ,TC��iK�;�:�p���"��� 6��<��G2�i�w3G���p�l�t�|����Nv��p�����2<��Wm�!8�iH��4rN��L����!M�Y�r��e~w��K��`-)�)�I��J��Y�TH�j�]>D3d�S@\Y���!��|	aM��t3��O.���G�QgW���1���C�Oy]Ϭ7Ͱ/T �W?W�<jhG~J�{J�ߌ�TE�E�����AŒ�^/Z�D:��
���k���d�߿�9j�� �Q%А���^ܾ�.@Iz3NY8ш�a��SW����yǯ�gq
���������.n��<Rʇ��G��� ��V�lD}8���J19h���?O|Q��:�/�!����άVKH�n����c��a�Q�>�ʬ\�X�I5)-����:����;�;q�Dz�dgd�\�Y��wۀS�g7è���uc�g�o����4�k��o�b.T��B�$���d��o7�K7��aV�%�԰f-%�=��?ح�]XE�y���(u,��2&�+����jM���Q���K�����|��[*��\���8�� .XR�~��]���b�=y��Y	���� ��=��zkZ)�h�(sq{7�����Ku���ޘ��vl�T ����z=&9���>d���lB���o8��+z���� G�
�S������D|���"�:�C�e�74�Ɯ��j���D��4N"�R4i��y��p߮���M��G�n��*��
�/���D↭ޱ�Jca��eey8r���о24m�gi��ȍ��yѝK>�sz��.�0�iWQ*n�Y�i%��D�9�Ky'4�s0�8�&��in�w̧��#?����%�9�?O��b��`����6&�hc�Ÿ���|W�;�$G�'q<�J!]�6((
�������/N�u�ng5.�҉b�b(���J;4��2?_暆�+��5w�l+��t3#��J;�$i�N.5=T|��!����1�fD��i��� GR*��j�j!�]W��1HG3# ҕl���B�l�Z�Ǹ�}�5܅x�iL74�c~����C��-u���J�~݅]��m�1<_��1�X?Vv��,j���q�� &�W����C⣶�������X�/M�󯌝�3�73�1��M��`)�3i�WɄcF��>�]=�U�#��BY�D#�]ݿ灤<�8�:��S�� ��ǋ����9�ˑ8�;�����U/���;x1�*1��u���Z�V��PN(4��l��eJ)���@X��a�!;�<"%��<��[�1UK�Θ^k� l.�q�6�l��`j�%�K?����|��#%�|�P�43����?6%��:��e;�;�q./��;(8j���I�B���H ��gOQڔ0 �}�0l���J��͉�)5�ZM(du�Oê��b3�T�8$;�����+�}Or���o�a�a���߇gi,�]��O��?r����e��q.��g������+���y}�/��L�8\<�T9���K���|���U�;�Y���w�����ĀM"	�+�-�1A�3U�j,�jу�́���KNB�Nܺ�i3�n5���<<�#FZ ���c��3��j����f!0o�$ txF�a�Qх��������j9����d�c�N�\$�x2����_���u�ڤ����3_���PG"3�Uv"���̂��-�գu��pm/��ـ�_n�����
�����>��BNu�,*+�e�t�R���6 �<=-��^<��ƌP��M4�5��3	Jt8C"ud�}wH���W�!J6�/����H:��
�v�$�7s9~O��Rb��2��W����n�#6���5�G��Ks,���|6�|�5.$|�@PS� \!��?55�{j�XѲڸ�n��GzKP�۴����5�IA}�B_�Q��&빏G�Jw3�i� �\��~��]�8c.Ҳ�M���x�#����BKԛN�@��M�s���Th�2�v-�>M�*��Q�̓.�����4�	3TV3 A%m�a�v2G���A�k�I��U�g4"�����msw%qyq3"n�n9R�	��Ѣ���t�H���Ђ��l!�2S�T���X�e�@��Ć��Kʤ�h�*�p��e&Jy�(�Z2��x��$;������o5����4���=&��H駊�O�����g��:����V��874${��c��z�� ?m%P�n�?����8�LjE�M���r偦��].�O��t�tY�Y�|,`f�<�Tˏ�RM���H��d�ݘ���=򱥹t�^�<�IBb|��	|A��%�`��pj�(3�Ѫ����慖��w�r�	�!T�'K=������nV����l�O���s�3 ���"��u�=KL���qB�f�LJ�	
��5���g�[���/��ȵQ䣍]t2�����̻�/k��@��,NW%T���q@v��#B�+�1��jE|<��ҁ����Om]|�!R?*�hRC�	�zd���x۬��L �ʽ(AM4uu���'��&��$�2��� 'r4TW}II���5� ���xB�ߩ�������yJ�rJG�ԟ\�}:�[�*.��GS�m2����O��H��?ؽ��0�~+r��GU�����"OjC�i:�$y�3�a��߱^T��2��X���u-$|fd��&�KT�1�@F�N ZYٍ��A&���9e_2�)��\�@�'P�m3�].��1Nυ�2��P3��=�$�F{W~�a��
C!yg�u~���l�FA�JE酏TK�8���!]����eXcW�xxn`u����F�5C�C��D[�Q�pda5��5��W�2�l��޷���_8)]MV1g���|ȯJ[~D���N�����.��7����@*���]]1�̔�%\��%!��������lK�{�KP�ɷ�ٺc.��7�Iv��9��IϪ�?��7V����+1��$b��HG^E�A�/`qdN&F|ϙ�Њ��1�<�*��8��&7&�` �Q���p)�J��\i�w��r�cŰ����.���<�B��7IG�h.���b,�b�a1��-.]�����7�@X&�jb������DLPf;(&�lX�%m<N�p�,��4Hx��:Q���gH�I ���(Y�ٔܚ�>�{��2S�=��\Y#ݽ��O*<̯_p�V�-��'Կ�d빃�(5�MdWV�m0Nu��RF.բ푔�� ����� $Mz�'�i�L|���R懇 _ͷnNGQB2�By���_�7^��6�B���rrX�B�r].�8�?�x����C������-�3�{��Fk,�sI�,ޝ��D��i��D�L�M<Z��yM�L|����Y�!Q������� ���L�H_����yR�%=����:��z8n.�`��s��)>�@������xV�E B �V'�ah�)�j~f�@X5�b���/�k��Xu�0?�r�����J�nM�_�H�=3�;o��ž+��?��[��0_��т�O�k�^��@�+��fՊ�
Vj\X>V:��:�����I_y�����o6��\��A���7'2//s��mA�k[�b�����9�aBX�����5�s9�!"ƂȘ�6��f��p�s�Y3Li�D%{&�����I+pAj�nݮ���C&J�p����&��>���9��G>p���;|ֹ��-r짿 ��<�y
����gCX�-���W�����Y��B�����0$��!-oT|9,��+�Wˣ����k� Vy�w�H�Aȶ��h%�j��?���{�B�5x�QJ
^I��,xވzt�����|�I�X��7���-�d̴^�%ngCu���Ě�S�����i_��s�.�i5�ЀX����ĕ�s�g/ �F��߶�U_�rƙO��������w�	�5��<�q՛����<�D8E,V��Ǧd�S��{��YXl<aRh�����5I�^���K�f�`�ֳ���3�2W��.�?���8��_+P�1������M��f1j��B�?�UH��4����� s��S�~^���K4��=��Ѯ�1c�3��L���)���K����e�Aa���g��qZ�Ti��_�����̷)���������E��<�ȭ�K�2n�)��dĴ� _tUQ�� ����r�?���xh+��A5C��N���K�.���w|�����3�IM��^t|�F�^��WSs�q�홭����6q�i� ��Ĩ����N��sH�=��P�rD�h�����A h�2 �OӭgJ�d�MH>���j��e�Z"x���hz ��;DL����֚BC7�Y�9>���g%A��ͅf���:`'��p�\��9"
�E�]ic%K���j7�$j����Y�P�!���t��؟
�
��X-rA�o"��e <U��SHu+4�¼|�m��������n�ɣ�2���N �G��wT;����d6ku��uh9ܟ�WT�nv����L��� 
�L�u�8�U�E%Iv��||�iS�* ��E"v����v�6��j������R���; U���ܶ�pb�I� F(�����d�C�,g>�5���wݞ�,�8u~�>w�#":��L�b�Y$Ԥ<d8i�q$*D_�����h���M����1౛ICx��g^U��Q�,��8 ���̀�p��mg{|s�2��Yp �J	P�:���s_�E8��N��? ���a��0����e�4H�cz���a;~\�ϻmu�A���ݒ�g�1;P�K��B]K�͇[���՗�{���M�<{Hq3Xa�ۓ$7>���aTh��	߳3߂;�1?��٘ 
n��@4�6f��  �ө�	�������i�U�d6�M{��NMK%�}5���)ݯ�.uRk|U��yj1�j���-������˾mA��G%>d��`��k\��Bo�WY��)�9�y��fi��=��!���a5ː�?6��%u��n3��|��rf�����t�@�x�FF4�69�1�x�D�?���,��6�d3_Tl�*k5�m�g+�w}�\���K����j-��[M���{B)���M�L�V�L6���;��DP1%n�W�'� ����x��" =q�q�p�p�����B�c*z��'+:��Ϝ�d��&�;�:/=�tCI�1�I[�D��رw`E�>i�:��A Agz�K&&,���1�,99��)k�k�6�ӝF�v�Q�6<6����|��P�4td޷^�i1�Z��"`��r�ןػ�2�Ñ�8Br_B�⏷�)����T�S�X�{|�y+��zgL{�KƶE�>~�' |�65�����݋�b�����D��i�45)II�����4@a4�6���1C��#�Q�ҧ}�l�G!C��!9*�*�b#��cZM�mZ7�z�[���
.�b&������ D�#��-�\ڎF1:C�|*�P��:�x>��)�9o

���ih�����^-9"O�]Y�,Ii�'@)�W�8m�8g��f.țc���\j��0�:}�6�V��Aƞ]Q��D����;�
{�6�� q6ܹ��\à�iw�!��Ѝd�Ҹ���8��4��~��4ӽ�RJO�+$X���@1�����	�G�4��C� �P��X����4�b��>x�c�̤���y^6�ǃ:df.6?��h�6�|$�O����Pܿx���1�Yǈq��Hs�&	�䨗[�1�f�&�>���(��@y�9�ѾP�R`��Ί���%g$�G��;/�i��~Q�ڮ+<���8���,x�A�官u����PO���� �E�����́��/��ߠ�W��mY�`��΋��VU
Q�	 ��J�b����`��LFFf�V@0d�� �K8��֊��}��
���w7�y	�o���.�F��yf���'d ���E�p�6KFשYD�ڤab�,��0�/M���(�k��� �����]��^��;����D��R� �5�x��&�҅ ����Ż�8��I?>����E/�4��p�Xo}En�DȱB�݈LDMk��9�|U#���1�u9�PK�^�l0�tj���n'�07���|�`w(��{>�x.�1qy��`
��8s@�nxi�<HPD�ɠh����������E��Ia�n�y���I��P�lسSR��&�b��aW:�.bw"�1���JZ�dZf>$�$Y��	`hr���y`���gZ|�����P`G+�e~�8z�mK�'�z�Iܒ-���P�>mS��h���Y]G;:-���B,�%��+�� ~ �Yҝ@��S�ہ�H=Mb�d��(�$��+O\@��d	k�{*��D��$�3U!�λP�m��u^J��6������HcIu~c�^2��tﾈ?���FR҉mh&��) L'�4({d;�"rTy
|��?�R�C������=L�n��Y��T����� �zx�ηt�C-~�����<��z�5���6��d��׎?����G���� �˞�n��N��{�����(!%�>8�<r���."y\�H�쏰Z�/RJI9��5�h�ߦ��?����zD�k��{��<]�%4Sq9���Y��;d{���p����я>�h��oQ��i�q9kC&%\5R4x�|��,�e������Kϛ�߯DV��~�7�ܧ�/�����XB� K"� �S�=�DN���8����;�)'{n5u]<��+��٣t�Ͽ3����wa�Io���Z�
�ƻ'6����v9%���
�~V������5��ҫM���5����U&�ŤM4�U۝��y�M�Uh^�t�l 򥖀���&���*�[� o��L���O���R�//$%ٗ<���O#�\~-M������Px����N���TK jK=����-�Wr�؆����ΐ��i3!�{��|7펺i���N�\i���5�}�}�*�b1*��[	�r�{CI��W�%�,%,�*Ҭ�S������B�7�H,��@\����h +�:�oRnmA�`�/&�F�Q j  �}~M��w��Q-1�l����p�W����`�^P&y���^&r����Ԓ��$���^\�
��ƾ���o�]M����O���"��e\~���Y�^�\w�$9�y�����9(����{oe���@`� %ߣ��cW&ĴAi�9m��X1io�{����lV&��<�Hh�+򈎺"Ƚk%����o�3�����p�����V7��Z?���U� �p�8֡[�2b��ͮ���X�i�Ps��k2~�a��<��N ֣�w��L�_ш�6�qp&0�{U����A���~�mE����i�#�����!�����%�I�!#kç��mt�ٰ�-��I�1�#�ZfIt �����bگ6�L����GjQh��2�j>��$]s��P�G���P�����8S
Wm/��c��������>��o�Y�}0Ww#�KF������ Ŵ��K1@�l�a��72F\�R��'LH��<g4"���e�ǋEirʄa�����Ӗ<H�K�R��J <���c%3�������;{r}�p�5A�/�R����v%р�ڽ�x!Z,Uۨ����0󮙛�S_�d&��B����B�H���D�2�I+aL �3CA��C����<[������MJ��Ɠ(� +:ۋ�R��L�mr,H���p�n� �Ky!g��UNAݪ�e���f¤�ݎ/�>�״2�sx4dq;9�`%MT@A@��*�P�kg}��k(S�ߟJ!L�%D���3� �%1������ȹ�m�3�Jһ�N��S��%,`�υ���q�_�n�[C/c�e�c�FJ?=젥"�oˬ�B%_��Hu%�O&�k�;ւ������^���-E!�q_s7��O�.㟎�'�=ǒ�����_� ����G�����כy�V�5`y��2E6� <��h��&�R�)���C8 m�R��Ke4Yᢏq���NBbsZ�ӻ{����
�;	;E8��-��E�<q?]��2��J��UA��/��*���8��,衫�o���H�G�J?�\�af���}�lY�����A[���UB���I�r:٤������`�l_�vB���p� �-����>� «2��D��%}rO�~�%����U=Am���
��7�:vz��*��ޔ���'y\��8�����$7�jŴ�k��TjAD@B��d��S��ֵ>���������$b��ߎ�W���2K Rb�e��/�8������l�d �=�.�Sl�f>2#N�@L�1,	]������~Z��O���<�6!��.��y[wU�`$�[m_��1w�h���h3���"�T��0�h;�X�.
E����dՊ�a�O�ՍyS�ԤW�_��jC�hoPa|���o���(�=�S9P���� ,C�*�k��dj��2^-�A�����۷��l�F�q!���-�y�a/�J�;�٪[��y"ST�Zuw}TB c���w��j�&1���s�HԨ�S��:�W��j�r�: 4,u|�]?��D��@b/��o;�R(��_ׯ��7|����5���������nio�i�Y1=��f[�p\-�v��au/	�0�SL��>�+�z��tq���tw�29�|�˩�c��p�'o�Q��|�"h26#��R��1�T�����o�Au=哃�ʩ{%I�׿V����7��Է�Ќ���@7��X%{��y��D\� ��y_��aW��M���}��ݛ+�GE����c7�?���������
q��vs�0�A��F$���a��3��z�	�:n8��S��[Bj����u��ί�_[��w �烘�..X�����`h�;����8hf(\VIK!P9��Vr:11Ce��ԝ!ѕ=b���Z�#��GPs�T�I
 q)Y	��<㩫���s_���qI�3�K��ͮh�\�ĵ-�2���*"�/v���#�o�E�����O�S�g:f%rn^֭=�&/�t nl�p�  ޸"KF}��i�3TR2�]��L�&p� u��"T�P%p�4�� ���V�� d�� 8f��l��L�e��c
E����2b�I�?�/���D��?i?U˃�I>/�E�k�w Yۻ�~�C����h}|�Zt��|��O�n0�$GU�;��Z���=>?}'ۆ��� ���C�I�kZ�\궸S��Y�|U�U�b<����M�#�^ oL{waչכ!&-y6L��Ndk����:�׹���8^; �)��χ�9�Hr��3��������z¤Vl����>)��7��Aq�sa�\�L�xw����*:��/P'5�|��nߧ�~fo�@��Qɹ5[n�-5�aF������_Z<���rR��K��m��g�V�ڽU "?�(�����;6�S(F��/7ٕ�4�l�0�6>�͒헛ō���h<,�!��������MOT�mr�F�yNTÙ$_;�2PI|ک�D�g�k����
Mi������/�(���I:�P��X�W�=���4V���m��Hq2?�g�\]��%��$��#9� 5���┬Lm�p��| ��AT��zg4o�o�L	<j�~]��Hx{���w�!2�1&"Ι���䴭�nb��]:b>�O^)��x3S0p���x^�N�+%	�+����s3:�#����T�����#���;{ǔ����o3e�uо���%����4��^���#����wT;����7�����l<7Fhf;[�����A��=�9�k� ί�Ԯ2yEF��q#����I�&>rt�`a��̄���l��7"&���iE�q���y/iM�[��M�B�2��y
�VW��V�2�9a}h�Vl�wB�X�JN��s����������o�������ז�)�^[��.�7������dNbp�6A1��uW)z����r*�x)�4�\Y�^I��"a�L)���<�O$_�V��[a�-���]�.���z��������Ε�w��n�6���`�m�f	�7�'�Zʙ��!���4���'�%d����F����O�E��<����O5BZ��n!*5�,��繊 p�g�@����8���G��ę���W+��41�p���z�|~��l����M� Y	������-A�`ɟ�jjEc���^lP�V�l�">� ���me�.^����!p�R� :^�M	X�ߧ���7�Ƌ؁5&�
?����>�d���L `sl�Qox6���v���~u��=�w��a��M~��N�c���9A�6폄z�ƙr�%�>u�n������V��o�B�G��7I����m�Z���v�i.b(���ُ3��6D��˞�_��@>wٌ�!����e�<MX��� ��d��!b|����ӽ������i]Tʳ�z����4�J��Ze�R��cQ�l+��¯Xp�\�a"�h2�|�(T���q�/O��{��EΓ){��v�N��3�ym�C��_S�'c�����in�q��U������?�sO��e"�N��)T�C$�'���&9�i5)�Ե������h�\�a�s`�7�nGu7gg�k��� ��M�J;�:
=�����E����-�8uOP���~���DD���tn�~�i��;�5
�ҡ<�~����/xb�Y�m��U��Q@��v-��E�]����&�U�ٱ^}����F�L��y�񜺃=� �h7�h�+t��+���q�H�݅;�ZPHU����c�������������W2z_y�:�x��7yjex�P�u�`�>~�e#j�w�t�(x�{��!_�ׅ��T����a���G�cڷiCM��ޕ�V:V�e�8�8�$B"2��%ʆ'��B3�]��
GW4<;-?l�vlUf�}�9��bh��K��5��,�E��\.
""��b�
��!n1�$T^s���\1 �)}�'���D����ۖ�w=R�����v��MN����5)��[�����#hRH�)�F��O��(��xU�^�;������PZ@�i�5�hV���&�rs��F�O�R�F����|;�H��k�8�k-wK
6�RsJ�y��d=)���N�7��%wpk�� ���4ҏ��hM��o�u�d1P�w��O���t<�۩}ޠ�w����N4;�x��W)uDQ��zLO��6��=Y^�����q��&9l��0j ��,�-3��:��ahn[�2��:��8�`C'�eY/OsÝH��lp��p�YYHH�����}]�B��sq��I��O�Sq$��iIJ�53�T�1�Q0��	i�Ҩ�o�)���\r��q���B?���1��5�0^ETw S���FEg̉~vF~�opg��"���j1�����%$n���`�,8g||w�����߲@BB�ŜEFz��U9�Hrہ��GɄ��h�v�a��޽~�1<��U�����wQ�ɐ��0l�̺2̠K.%�N�|9���掤|�4�aH�=;g�wW�s���I�ZC�Kg,�"{�o3�!{= ����p�h3�]�8i
pD7�̒G/�d�k���<��U��̋�o\���ّ�F pi��?�	��i(~�E���w�7l�T;�顫��FŒ��\��'�ƭŕu��]�����XkO�$%��/G{��>�5qo؏W��5�w1��e�(�qil�K_�[z�YPŌ-��I�����Y6�;r�(WᱜyFC����y��m:#�����iA�`�<�)x��sk��;\;�9�K"��z80�S?�V��*��`N�|q�{��Vv
�=_���	h� �Ӂ������s�J�[��+DUr�l���_�!��&�}�!J��Ea�U�]Y�ܝy�z�B��8�9I�`����y��T>�����،w����e��neֱ-p,�8�0	,L~�j��͑��	$ύ���<1��w�+��束�dN\��)�������T��(D}�Wv�G�ukBe��V���e]v��/�t�p$�3�����x T z��JI�v{�8��پa�
�����&j�)�z�����~GE�a�8�	]��r�VR�Κ�w�%sݽ��������\�oeH&�7��^���n['7���O�f�ndu�m���9Q���x��3C�E�!��$u��{[A�����9ش�.q'Q����c��^|���a��]��������iܱ{� ���H&}
 O|T�Uc��_�䡘��@����.�����[����Qmt��;T��aS\+�I��Zm�~g8{�PTLE$E@�L+�Y_�R���S5i���������uP��U,R���_�8� q��X	�?=����r���uJ�(�:�2�If��#��Q �䡻}����w��*R��=���!UYٙ��Ƞ�i:9S?D�2O�����G�7#g������W ��G��	�����1��cַwA��ǵ��Uψ<Kw���8	��ͥ��?{ƫ�߽��m�N�O�d㭘8�;��Jt��Ib��? k)��`��U"we�TN�E������u8����$�[�5V��_7UJ��g�0結"���qg�tr���b3�O㡩��h�+Ӕ�j8 ���QẏZ�f���W@E�D}/��R(a"(�"���J���(,!%,]*
J��ҹt�"- ���R²t�7�����g�g�ν��3�tS��.[�(��V�j��G~�+Xak�F�<㙪���_Wg�&t�����4��O8�`{2�i,H�\��V_^�d��O�D�5��s oH�3;����d)[ �g��FH8��+�r�q������g9�n�����sC3��0O���)3��V%�Cv�v�a��&hE�󎎇�<����s�3�|RU��y�W��ϰК��{?|*� ����w��1Y�_ YQ_������4�\V���]�z�k�������Ťܛ
�����˗'>�)`�bL:T@���j�捸���H;�2��{W�crJ����j�9"i#�O��f�o�6�^�N��=#�;�I3d��B�+�H�ڽ�څ�q��u��0Km�r�<�x�M�Ө��b9`O��V�
�E�҂��L&�Y3��I`9PkK~�vy7qp⃩�А��`	�ڈ�ņ6���j�x !P�����e?>ݜ��}A $/nR��d)i~��b���8|o�pws���6j��t�,mӾ�������`����J�To�/�I������XѾ�R[�9��
m�R�2ml���.~���CdD �lf�83P��ų��EG��Mۛ��O��*|���O�B���{�L����l�\�~d�� �튔�d� �xjLEY!u׉�r7y�P]�j#I�45�i�*%�}�*�\�EhsH�_����䱽��
+cM�g�05��Qa�K�0�"��I�N�Z�^��5,�9e��sx &�}«z#�<d�,�zg�S��!�������sT�(�)�����:�T��w؛�5�\׾"iZ�����ZE��JnM[�@��)w��H�l���D�i::���F11�=C���l��{�6�*�`)��/�b�7�v�w3�;��8����Z����Nt�uW
���]a��y�qU;� ��PL�rM&�X�^l���s�5�-�'ؼ���g���~�ds/��rJ�X\��V�y�d!Iv��V�4F�^�0�f����q��kGu$7��D����~L�E�q+7�9�*ӹ�����t�C���� s\��0���O�5��ĵ��sqIqlF�.��zAƠt�v:=��uvz�خ�N��S�.=��3��D�7&��n�
��F�#�~l}�'i
o�B� �+H�L����.�&�5�ٌ���<ԓO_h��e2������F�u���],㪡���y"x����d�\`��/��~�u��&=�I{{!s�	irµy_Ĥ�M�0J�ub����K��E���rf����^DJJJd8%�0�M.���+����fo6�C�z�/!�ܥ�T,$�>pT���s����U��wS0�9��<Ѥ]w��n�a��ߓ���'䰌3[�ܿ~?�;s�V1��C�k�C�S�� ��$)��{6VȝF��n-~!c@��Y�Y���l�櫇�o�/��h6��橩+ �%��4�m�q	1�����|�~l?�n5Oh>�Z��x���՞D���_��[d@����ߔkkl�I~��ϢoW��4���Z&q|`�ϋVnH֖�$����yӄ��c,�û'�T���E��9��U�l�Hy>���F!��X\�C�g�@	��m�҂eI����c�jrʵ��ˮ��Aw {O6��^ql�U��^8s/��-Ȝ�+ȊQ�W
%����	*��=)�����J�B�x��y�հ&��Uӕ�c�_L>��E���^FLg���1I�i��n��G9��؇�g�dX��ԕ1�V3U�яٳ=s�b�c�`֫{�^�NF����KYʨ�ӭ6ey��i�)��=��'kG�����Qn���{����N�r�A(���s�@-ほ�+������[�솝:�d	L�BӜ�9�� ��\G��\9]�g���wn鍏����/�L�>�{�>��|4߫��j�!�,j���c��S%��M/h�}���;�6#��3�zhk�Ws��<UV�m��7�hb�"P�.��E��[��Tf�ӻ�P�<�} �*���MjfxB=���L �l���+�ȈPo�%����_:4����3H0^���c}�ڭal�_�հ��nP�ͼ���.������n�x�
?����/-a�c<���k�ks"uȫ;s�Y����:ȟ��p��Kt�u��>*p#�\�Z�p%_>)Ql����x���#ϳ%�W3��f��_�`�N�)Y{���.�(T��;m76�>�q����3`n=��m�
ڬ���|z���pc�C3�.[�d��I�HW�c�}]Yʑ5�\d(�� ���S�?28'6 ?��e�K�`=`k5�H�{v���f��M&�����ZE�balEaj*3_hX{�V�̌V(q����6n� �2Gv8#�4����W6]���lv�z ��R>N�
�b�ܗ����S��<U��ɻs���1���:ås~z�e�RfIM�cޜ��j��R�\�u�I�rr���,�!�kAP+0b�bι�������y9�R�t59ӏ2fr"(��E�W�tLؘ�쐮��WT-��lu�1U�y�<{��Tf��7���o��� ��������1�YFcƚ��C���r���w[h�X���U��n�n(��'�'�����f5f� U�q.�4{����:z��3��d�}��"�0mzpu�mO(���æDm_D\2 ���;�B� W�H���F.F����;�_\I{)���̪���˼O�]n�b����
H��:E7�˷[�X�# �
P}�N����<{�U�\�s?{y��ؒPC�<��,�&��UJ��@*%�8gv��uc�<�뗄*������a�g�j��\Qٱ��೙�����R�wF�m��40?�Cl))o�����`+6�f�6�L���cP�ic3^���Y|Λv�=��D��]���|&�Z8gc�B��F��s<����P@n
W�x.�hi���U	o3E�H��S	����SuRIA���6�=�΍�Sq����Ԫ�p�c�)���9��Q�Q.!8�]�v@_�refEj�M�3�>���*�6�l�:Ru$�r���*�!�����V��4��[\��ɐ��w�ә�N*����4�IF[���:٩�l^�F3�'�׿��	�*]��zN�ոnS��\�Cբ������:���4e��X���M%Bt����$*��n.���X�K�?��:s&��ӟ��R�K���k�e46A��zė�C#P�gu��j� a��_�����"鑒��(��þ�`��������$��_��Ԉ�7�B��X��w]W6]��e��� ;T$6�q1��l]sjC��&n�u=��צB� ���)�c�����4&��[6�g	ej܁�@ �X�ȘA!h�P|3翍hQ�n�G�xu��@��[��j2{��l9�W�?���P�L{����z�i7���Ź�H��5�
f��&؆��x
Jm��VI�+��N�����Y�����{=�}����Jٶ?�j��r,n�u9ص�#�A� ��2����t|F�T���y-�����V���{��V?+m�4NO�A?h$ L�p��U����>�m�^.�S�"�̇��LvW�Z�c�ֺ���\u�$
��6�%#K�Q dU'(~%���\����'��"��f�T�����O$kL�x�8�AUA0�v��>��u.�Zԇ�~_��D渜�X�쬼�q�]�cLeaGc�L��g�g�!�� u�e[���מ�7{d�nL-7��4�Ue�p����Z8�~�������w�� ���䜭�H���U�S�k5�T}�Vٟ����;P�Gv_�+Xa76�}�A����nD���CU-*�5Z��]"��9❁�/I�<T��>'�
���b�gYq�;��2�W�`9���&��I��C,Hثē~*�J<�JƿD�x��1��Y�{��붧�Θ�TCzu��Oo����ǘ$�j}������V�=; b�"�����kI6�V"��y��*F+������	&�� ��~��b_j�"�k����eʩ��V�ŷL.�\=(PZiHA/��?��s��nO]��R�]�R����B����)�8��;#��/�t���"}3~U��$��KcM�;�r,�Fo��5�-�ˎ:�A���A#� /d		Ji�6(�Б���N
��v��+	����^��S�5!g�VvWV2�)�Y��We`�<������:y��B[2��M����7y�����jV1v~��M^��n�^ �B�g�0�NASc
��Ӓ�M�T�ڲlj�?uڶ�z���hk>.�ڻ#�[ڨ���o�*5X�W_|�g���:u0�?_	é���v�!&"C����{�qx�A�����w'�N�FN
A�����H��#�cktwY�W0`��NBD]���0�8����顃�@�n�&����'��)=�$F�'`�Oӭ�+��ސ��i�P�� �����7�AS��m�n¯��H[������?�>4����Is�h���r�����D)���`{M�5j���N��fG�z�������\��ޅ��z��B4IA����}[�/�����K����6��U�@�f�g�
dN�\N�yߵҶx�o����΋I`��n=��r����6Y��ݱ&��<����R�{�j�
���j�����F "'bq�ރ^�(�-���H+��mS%�*�/D�����2Om�:��l�o ,aj��{�KL�[��+O9�O���'�:�Vo&ݔs2�ͣ����[���=�q �E��d��C�Z��25�k��Ƨ�{�2��� ���aH�/��� u�o�B��3�i~n�Vf+}�?�;��[�@�����ZW���#^���Pzv�>�=:z5_Vy��T�b�	qh�c�(o��.�YOX�b~4����˕��@�0w�&U��%��ά ����qj�ګ��		��q�_'d��ղ���W���p�Ũ��<7׽��>6����?�yS�+�#(��}8��7��(U7Ve�w��d�� L�L_��J������O)��6���#�[ͪ��T��V{���Mп�0��7u\g+f7
퀑��cԘgeӌΓr��F�r�e�?_:�4PE֛FΆ����K{�'���3�����m�P�ϦE�x�*�k�.a��C�Xŵ��� +�j`f�]���%�jp�)�:dc	�@��wЅ^�y������t�_G��g;�[ozj�f��U��_��G<���ϰ_��TA��59�'��� ��KJ�{���G�`��q{+��T��.vw;�ٱ
��3�0�II�HR՛>��S�V%�@�B'w���ȯYBV�g7Q��A8!P�!��q�L�K���Щ9�9m�Ӂ�5��壮��D�7���惒y�d���Զ �6�퍄E��X�J�;ee3�;뼛�S����<�P�?�Ʈ=4ͫZ԰8��N�jN[��J��Gz���o�Ō[����!
aY2�?�TD8���4]1	�����_:C�.��v�kP������K�_�Ģ����tb꣝�zFtS����H��s�җ�*+{����O�a�H��S��:���Nb����I�G��\r~�\٪j���}nW^Ch�M�jif�lɹ1a�p��i=�)^O�����'���.���W�BF� ��vk;:+�b�j׀�`P�E	a�R���Fv\ߺ$�[�|��2����N]y�Sf�rYb��C�[/7�q)������S��_�t�š���nB���lN�9��O�ĩ�~y[P��&������J���^	E������4	����ou�~/�V'����={ߝ݄�h���{��Ģsv�NǴ��$V}�%μ���J7Kw��6��a9`BRO�`��4�E�����瘖?�nOۖ�Y�ӿ��آԘ�$|���
KG��0z����5������N���c�Ϳ,�:����y8��,F-C��ԌT�5��%�������8�3g�`M=�M�G%�qu��!��T�����2uj��܋]j�6X�tb���}��x�c9_��#�FC���y~�_�U÷��te�$����pNi ��'=�m���T����J#����n����_����2�fڋ�;oPL��UmjX�ׄ�'�1җ&���w�ˋX��Іŋ��<��sخ��-�1q0f�:�E��Ǩ�Ldl����щ�1"�n�u�]v��aaU�NCI�?�9-B��S����WS@���3u+��k�L���4�b!���ի�j���S3R
��e�r�?��q �}�	������U�[X��&���BW�ܒ��� ���e��A|i��x`X��O8�Ar�D�T�#�����q4�q�w[��J�o+�x,�m�{����n�%d�Б�����Ā(��]�Z4��W���$�>��RP�K���R��G�z���i�"�Dl^���D¯�n���-5b�^�O�j��K=4�2��R���6�x�SU	C�h��̹ӋVd6�]��}�.��E8m���R&��엽 ����}���"3}�,�$�N��l�{�<�e��|�}X�PbP�/�ӛ�j৆x'��RƇ��U޷ｍ^P�Y��ɿ��uN(�!0�7N,�sF*�e6@�q�o@��÷b�<n�w�tו�Xȋ���d��������-X��R�&^�����iU��_S�p?���#��ј�)�7�%�jg�ɛPo:��e�،zD�@�*r����K����v��+�N=3�x�<� m��g��'Ei|��y1p����u�ݳg-�=K߹������h�X�����VW&�s�DGk�Vι��Ea/�l�V�U%�:��Ja��-@�OD�ϔsħo'���͡��}��gDG |�s�p<I�"�lˍ"V���1��?��G�;t�u��&�a�xao����O/�G�Wr#YP��W���$��|J�F�+�ȥ 5H�n�iE�8)ʬ�*B�I\�v)����K�<����=��jT]�t��X`r�@	d�t�*�j_ xd�DQ�cڛ�q~\3{.eTnl9���/r�p���k!7b�~��Q�#{�Y�5�G��Fߞ=��fK�� `8^p����J�}KYcO?�	��|�;�D����"=���f{�j��.����ט�����=B�P�glun(���S�|��U�YrZ_�j����KbS�o���K�A�R��.�Ɛ<��_�:#�vw��7P�$���O�}<� �7����EzMdBt�`�({u��E�%���}�&&�zV+�)kk�XƍsW#]���2['��aхnŨ���>�%<������Kǩz	��ƶ6�	��!Ju>,�_��;��O$PPup2"C�	:�0�^ ��C�].b���q1Kz�h��l��=S=����}��`�:Lx�����0��P�w8q�y�����%vz��w0��L`)`�~« ]���F@W� ��\$~=|˘�z�"qX̏���An��ű�'M��m��nm�9�y�� ���uR�ܪL��\�i���ߋ�{@��ҭσ�?.2ڣ2�	��C=in���Y��B$�q��1��6�F.�}�X���p�ϐ�~��ۧ[mvP�]�	�����aTG^�K;�c����X�B��`�`���-Ŕ�V8�*H	eC���<f6���F��@܈��wٖ�~q��G����f�4q�kw�������֎G�%O ح�d�Y%x�-�D�Q�|�P��~N����c&Ϻ�XL�����V����ɳ@���fS8�2t�~q������cs�U4��P�U�w��_j ���.C��hD����>\�\�T�Q;�z���npH|ƭ�R�^e�3 |��B�<��>��u�a�B��^ɏ�hv�G�W����n)"�QԮ/��8B-d$�����Fv/4�����J��~��LoCH;V�s����۳��$7Tq����<E�c��-���A;���hY\�)6k��C�� �8ؽ>s|�v�˓o�^�}c���*��ph��Z6c��&�-F�\����eϡC��{�ԑ�p�U@➢J -�o�"/#�)�46���}I�w�5m�,Y�1�����-���� <���v)�*���q�f�@��@z�� �J�ti;7fGȫi�U�xL�a�j*���a�Wa��5�3�5�gT����N�ԲCN~�g���t�c�a��m��]'��[�
:`�#e�
��m*/(kk�����ۑ���د_���y�bGh﹯^�k�y��<�H.�'&b���&W����H7Em�i ?���3�l:)-�Fg��	i��,ɇ!�k8
Ɏ���'�V��TSgg�t�b��]�ܯa�#�h'��z4��~�3K`~u<���"��2fa:6W�����Cl$a<��-!�z��5ם�l�[v{�4��)��������N��~C��
*0���	�g�x�%3�/+�Qf��N��G����PPU��������i�H6Q�����l��%����Y�і}�>o��S�� 91�q�4s�� ���XF���o��MVAq�kʜ@�z�܃ni�r�`�'{�@M@����4vTW{}���6FQ�Sߚ#�~�o
:����X4�e����<�=�G!�ȯ��b�e���HH���m��X�H���K�?���s M~A�����-Ó��@�t��O�0�n���W����ړm�7S��}|*%�W�g����/��G+5���̪���<�S]�7��K���`t�x�����u��|���F�.���&='߱�>�gO���!x'�`���g�/d4�:�����]�b��%�:&���#�;<	:��}ۑ��x�+"IL�����5�ǀD���^�,J;j=�nr�)��?v��Z�t��1��a�?��K�b�c��*�(�l�������v�6������{�`"b�ƌ( ��My�~�gh׼�i���%]�<��ڒ���it��_	G����_)�M5�
���JYɱ� "�շ_;1�U S�5�3�PzU��K��:��(����ͣ�(̻芩�'NiPg�s?^�I�`�MIá"���8|q��Ô�P� ��b�Ǚ��aY�"Y]�:�ٖ����a��}�y{T��S��1��L �]
�,���9Z;
m��ĺ��� T �4���֭_zD�L��(��K�D�q�G�?l��А�?���P\.T�U1E���l5�`��+�n�<�UfR�~�B'�g�9�Pci�E�/�Q�[��r���3�?���︌�����V�=�61��U�A{� h8O�?k�aZ�/�g�2�C��4k="Q���e���R�BG��Vk�x�D����}��%A���+�_��X��;��Ӽ<�ao%�i&v��T1w1��c�	�S=�:�����Q}�>����P�O���C��~.�R�t�6=�&{���^.o��z���G�@;�.d���z��xh��
�_��E@I�ɴӠN����حpm�n�*DP��'"9���Ϲ�~)���X	�	�7c/x�?.���Z9;p�Y't���i�֦��e�ũ>Q�DI7�AL�l,1vy+���U�K<e���i���6m�G�J~�ި��i̪7�>u� ��>'m�8,���k�]D�m�n׺UY���ÉӃ�޾�{9�����us��c�)�ͨт_�D�܎lʉ=��}�at~bf&��DM� L� Ŀ������s��������K����zn};�y�^��p^���D8}�ت:��� ��jⲥf�<�Y ��&�q���O�n�4�\:qɳ�����;�!��L]=n�޾O�A����]Z�®��u�����b=��4�ßSi����!�x/�`|d"��������ƌc�W�Sı䶠�����Ƴ`�9�Ӻ��i�s�S��`�+�¤z�8BGQ-����DzxX%ou��fR��G�dKeWa��������������!�I�XN����8|/p3f@#��' ��
C���n��7\L�i>�(g�M��IE58�ܭ
�:ni^^�w��E�_�}�ݛ������ȝ�h�n��2c3J��G�}�(E�e5EF��ـT�9���V3��������)X]�7Bb�u�3�⹧�$���C��� 0<����I/�~8=[vz4LE�^mpt|��z/����<�I��;���̩�wӱl���@�U�zߠ�����dP��bDM:G�H��V�2\`�٢+W7J0���R��-��.�*�����e��AFO�PP�ꌮȾ��J8���2�G_Ei�,���?ܽ{��TI�c8�+3\JZ���d�u)����Gh<i����P�G��7�ި�����ZG��>�O��C?�L�1�#�t }�r}�>�hC,/n��b��<�Y�����Q�I l�mU��ſvy��x��خ ��Vz-�/0x,���Vg�4�j|�]�r��������q�,=�#��m���i��(��.K�X���/!���l�n���~��3�p�Yo�G�����jk �IBٸGN���9��8~&�����_���y�C�ToX�,p�l%!�� ��r��C��מSi������)�=�3U����'�W����������"����Q���ܥ��D	(�n����1G��̀T����p����0��Mfx?O\�� ��K&�b��{*W��f�oD�3�܇��Z9<Y�9N�P�f{�XF���� ��W�����d/*�CْvMMA��ܽPO�������?^&^���C���m�o��T�9�N<��G����s�է���������'��z���ٷ��XF���SP���&�<��a�@œ���I&�&PQ���$-�]'#q,Q�N��A'��#�򊋽�'^��g*���n�r�K�H<'`x��j��r(�ˮ:Z����P'
A!@�~ߡ~^���s�����d��sxa��8����8�{r�Y�g�n��#w�R��+�U`�4�0���_�E���l�2g݇:r�u�_�$e��4�Ī���E��������H�Y1[ޚ�����<��y����i�/�y�(5���Y�D�Ϭ�z�1���j�P�	G��X6�o+�=��#���e�|�Ъ��R!���r���,�Tǌ�#"�?d2h�ٟ-n����1A~>u���u��z,hEAb�3�T~����T�U�Pp<o��oI`�<{�E�9�Ӫ������0U��D��c����r���n���K�B)h�tr/���Ka��G��h��xX�o[�,>�>�z0�?�����FC���T�뜪g�8yߩ��*n0�7A:��oZ:=�i�}쿉�"4n#Ԣ�r�%����bE��=�O�u'�D�? ��N�==�a�ݵvV�]T�)���
Q}h��M��֏�i�J�^sH`e鍽�]���ˁ�qeC���&0�2����.d��R#错b�t������xM��Ǌ\���b^�����_W�?[��j�sn4w�#3��;����9�1 �}8�4�.g�L�'����8���6^J����W����~ח�Dm���:k�}E��r�=i�w��ꗦ�F��:�ʞd�T	�.Z���{�u/�2���s�Xs�X�ԕ�9�����D�K5C�8����u�u�V$��ko���7�r��yv>��':̼P6M��x�x.�K�0�Ƀ�W.'�Ϋ������&��ۖc�S�6��T�ODY�ž�Cݶ�M�h��;�J*1z��P׊W�?�k[��	��}��[����|q�9��R|Э�4�r��)f<�eH��ӥ�Vƥv+��>�H��c�i/���F���ng6���`x�t0}�a��H)���ڣ�b�R���9h�B���U��}���ߛ�����+��:��m^��e��[n�(���u����ߜ���')ٺW�ڦ�E���@|l�^�J��<ڏa��O=a?K��ti���g:1ׁ��`�8�'��{�b�qy��T�^��:��ؕ7���<�3���a�&�w6�Uk�oO��n�M��������V�q�_9�$��@bd�l���~�{o4�G�]S͑՜9����C��γnQ;?�3Ψ�b0:���j=>go���J�ԩ�y ������Ȼ`�L_X�$��=/8�ỵ�'�7p]��OK����U2͑����q�`zL�ã{�[�U����� "ǉ��w����%��ը�ٰ0��H(���}�g��R�_�o�:�K�p��X�j���
�-� ?��"4�skS$P�����������?�Tθ�"��|��t(�h����首��J L�K|�}��1I9��T���!-��B�&ibb׻2t��ֺ��Ɛ�a��Ҵ�d�2&m�&J#kC>H+��]����>�N���a�B�%X]l#F/��j.}�17�C$e'��E}c Xo]�������QK]!�E�0���Q�unk*!Z��#2yK�� �ź��;ɋ�f�c��-�j%-��iZ��
�Ȣ�ǽS]-@���^�b=�@�j�?,�����`��Y#�h@��G�ygښZ���?
��In�a��+r��Eb��w�x�I9��s��8r�w!�ȰX}"�{��B��gْK�H��|x��m�F�X̊��3��:[-�d#ơ��:;m�H����3j9h؆6B�����E��צi*. ̟ս��E�8_nִ߳X[Xgbx����-I����c��czlupSi�L�����ZjsM�UR:�4��Q�_�}<��z|�M�9Xd"����U��);�=�y���uK� �;��`0�7�V��]I��� H�,g$AFL�r�ޏT�"�+΀{i�����
���.��6\'숥����sw�2r���4K�ۦ��\J �V7?��<��[��w'�
��3����H�$����g�\�?�  x����t�J-~�f���M~���b��\���Ŗ<VN䤩:�jy��&7�f���P��g6b7�m�r�b��^=�Eh�_P*Ԛ����������ح���{A�W�;k�9 ؽ�1��	�ټ��"��?+�~NG�y�.p-&`��8�� $�7��7�*�ZU�����[,)��w�F�&����D��	i�Lt���(�%����� ��ɋω\�_w+���xg�aĮ����l�1Ƙ��\+a,%tR����;B�;[zEǇ0/N�����P\N��i�P�G�y���Mm��Z��[L��i�ÙP���wZj����Ȑ@R����y%���sA(��'�\���̥�4E����U�ZW�'k���[|ν	���T��y�����Jg�����n��-�[E!n�z�zKGu�r�wLy���b4��(<����K^g�]G��)Lq������W�Kso�E�.g&rK�5T��������:�SRRAk�hG�?eT�w%�h�+L�_�����ۙ!>�嵚�z]��&Xo���讐Jc��\��`��ڵ)`�X[Th[ѹ��B�J�Z�*���T��tl��>{�Ჟ����-�H�KF)[h�;ܦ��1_X6�W/R�\��\�
%��ώK�r��L��"������vr�K��d�&�`o�������=�4g� �f�s��&<�Z��Ǎ���U8�6A5�r_�������_���.�3���cDʵ�Ō� "^N eK��f��ܔ��~���tk��������W����0�4wu=HI�л3���x������#��`C��i6��}UP׸�hV��)]_�������[��Wt�#����x���f��	}�'��b���N��/�b\�a8�G��~�w���p�U�\2f�׾�g��<����7k���c���^�2h�>�B�Q�*��ƭ��/�[�L5���?u�fi>����B�\��Ҋl���e$:87�!l�T���߰.���<�p~
�t�I��������sہ[Jr�V� x�f-6x%�p=��uxή9;���3�k��o�C��nሜ�5�2����%l�Ur����9*Fi� e gW���#��j�H3������q�w�i�O����_�w�u%BE�9���DiW ��D�)�ǧhj��a�#Y
;��%s���^�O	���V%Z�Oe�gU�=�<tn�?�������˯z4�Tn�C��ɡ��Z���1y4�o�[L�H�p��}]��4K3�p� ���r�g3�6
V��ч=2�h� �?�.Ֆ����"´�gV��"SL狼�+kk����4w&������%jo� ��pӸ���^�C`%g^"[?qT�A(HD{�|o4��e`�u˺u�{kS&le�l@� M�M��G�<$&'_͊F�	��U��~Z�
-����e-��j��tx��hi_f��H���AGN�e��Rϸ������Ts�~w$\�� ����Z`����s�tn(�#��� (F�OdQiή�3�\kt��<��̱T��M����&�ô���C�j?Q�?Z��;t_뒕�G��ࠇ`��~ �AOs�Gj4��9����	L���N����X��G�T��D��D+�u�_Hd��������.clI�3�(Z���%��.x�	��j,@&�M��,�:�Yo�;%��?hO�=Υܜ��@�)ˇ�!���.�ɵJM���b�.>�sX�L���	�����]��^ɑ�?\}���5s����s����<���m[�z�I��cW��NKxAS��N�y�f�}��⸨��Km-��5�
�{�bJ�3{��
&�'���?E"��)X�s@�D�cD�U�P������lvV���a��]���g�\S��E�`�~����P_e�x���δ��y��<+5�A��g�K�,5��^VͲ�l���]2�L@�:K~!`�����I+�~�� GI�%'H$lyk��u�E&���D�^?k��'��a�����y���ʿ�6B�#wf��G����,�zi=�AM�8,K=3}�L���=)��`?����m�'!Ht��9���m�&ȍ�ht.���g(�ʞ�(��^ټ���S5p�]��ZG�\�N�!7� >�Cf�g��<��+�ʷ�)�?8��i���p�kC�Q�)MSZ=����`��	6z�{�0�Q�y�K<@20~�������������V����t�����3gZnq��I��Al=�7#�|L;YZ:��}��n����"{�c�u,�8]!
݄�QŘ�Y=܏f�D<��!'�*o��y�]/���*���,lKd	�C sV2õʮ������L4ە+.r�����)L|=��-��M���Xh
��պ G�k:�}e��<�|Ұկ�1bA[(�9��4K��i���Ol�g�_��I	����&f`>��96�^�����9�cF������c��w�֕5!m?-Q���m�"�ZՋǿ�Dw�u�IH����^�}�՘��K?�@��e�0Xg�s��H�&���O]~�����C�t���o�&�o��!�i�|:}�"[�d�F\���Q���"}��o_i��e�Zv���x'74�W�]�~g��&$^9�ڇ�[6a�_���J���H���}c���j+ל�ZYo�V8I�e��g�}��SůFn��ߖ�"�e� ��Ng�'��T��úW� ��|�/�.&�?���5�h�g*�?E�x���P��������W��-�>��(:�����"�Zz�h���.�S���[8`�yz�L�+�4��>\��U���h}$�5��a�����+����� oNz�in�����l�4����%D/b!FWVЌ���je{M�����O�<R!_[P�^�ہ�9}�Д �E� ۿ��$��y|��9'L$���_Y�3V�����t\��޿C������z0T�Kڪ�M�����0х~k�H��#�C+��RW�FSo�w�(�WM�54q��P �'�lGD�Z -��e��FP\9�]{�������Ϡ����Vƫ����UT�6�L��q�	��&d�X��	���";��>�iw���y����p�q��Ahx� n��wɚP���Yt�m�|
�G#=�y�W!`j�;�u����C5���iD�����6g�tu�&��"d�7�\3���"��z�	� " Nɇ�P��4��R� �&E�{K�H��4(���u�t>1��*w����<E{r̻�j�Y���iq��w��E��yɮ�7{�p ���I��*5��MOG��7�a0G��?:�ݥ��F�A�
 I ?勷�V ��~m�6ȥbh����V�Д=���c@�y�i�X��������Rӥ��}��-�F!��c��ыR 4���e��u�믋0ɿ��zP6�d����}�&�ul���!��ٖU��������5�L�a:�e���+��C�psGV��j����� �*%׊'��2����t�f�[å�M��_ 
[k7�*��0�ȹb���[�](UZ�c��Z1���C��Sp��`��;�޷�0c��o�"��ϺU���ח"���:�+~�����H��`��m�9������u���⪷֤WʹŊٮ�&�0�J0����|�ù���[Y2��;���Os��#����쪴�M������I�ѽ�-�� �0�L���g�n��������b��{	�t�ţ���C�F����I�q�x6���R�j�f�	��x���>X��u{�Cթ��qj�7�VD$���2ʎ^@	���Oj�A镾Ktq���Y^"�w {4��Z�{�)�c�k3�~�����ֵ-�䩔@��+�"���_�~���a��#ڋ�T���g�xRV��.+��׹hc40_�b��G5����`9B�.�I�kׅ
Y����;����灝���U��c�|W5����v����1�D\��4m�.�R��������z�L�t�@�re$gWC���5>�����Aj����p@�P�� 5��3�m���� �Z;hob�����T�?_ �3�0��e����Y�nɳ�i�FO��L���^F`:[�Г���'�
0(��!�``fי)��=�2*!��9��v�K��/v��<1��78\�w�8�?a��:�|�?�ѱNo�>CjDA%��b�+�1������
O�ݪ1��v[`s�����f�c!%�̾��P'���}K�+��-a�bX�I�䆳����cM�|��(6�l���BP&��󕉹s�%�i��k[��J?]�v�+c�R� n�~� ��[�F֚Uo�B����>@��Kej�� ^:c�gi��	r'>�����L��A@t]�3,ƈ��eAJ>�Ek�CZl�!x������\=����W���~����q�ǹD*�YZ˄@�I#@��^w�7cߐU|�V��,jI���]O��2�^y��9�v��z�y�;�Tw}���co(��5n�OwW���lF��'P����lEV��Z����iI�>�C��ճB�{{4�Q�7��2��԰L5w�4f-q µK�,<E#��xB���wb��Ʉ��}�Oz~������f�šN"���3���0^�R�6J�a�w�тu�t�.��;��.����aR����y:�p�*�n��B��vۅ�����#uga0������ήÍz��N �ډE,|�Zp_��1�ɐh)�(�[BYW*��p�"PK&��(`I��څ�}�x�lzɨ�e����+������Y	J�ox��ЬP���<S�e�ф,��4{��t��m���Z���r��9�\P��S`��F��ߓ$��pso�;h��(���M����<\eXT]D@���C��C�N鮡CQAR:�����:���|���<23��Zk��F��.���m��öNꮨ��j��XT�j��5,���x��.���L�,Z<�eG��oQM�,�������B�_��On�1���$"ҤX�� ]���x�6����@��g�� �s����
���(u�a$���O�&�9��݁���ql6�C�����P)���n}8����qU?ȕ��`��f�㨷r���5��p�<:�ڍ�9�@�Ӧ^KY�4c�;!&�Gv�@�[�p.B�aN�Cy��-�ʥ}�Y2����c�W�(ZS&���������=�@�#�3��R~������WA@�,�,�h$F��P���J �_���8�ʡ4)ܑ�������UE��ʡt����������P�Ii��5_�;x���hc��)?��|8��F��]�~��5�K<f�� �J���F�]݄ÿºiD��V ��ih���DĜ�� +N�H��,��i,p�}N!¬������P�
-�D®���%�жj�.�54X�h9�@ ��k�փ��Xy�P�2@ުr˘=�� ^��"�T��[�tfh��ه�G��Z������]a����ԟ� e��qڕ�{�������5w�Pn%B`Y0p�;�T־6\��
��U�L�&�� �t� ЄWi�QaΓ@X]n�S�]��'o%����oM��3��s�ZI���`h3g��Y�;=����K�?t��n��U&�Ո(��xx�Uc��" ��E�\.�vZq�ȗ��#�n�%:��
l�@���`��Py��鳅�X~��ž��3r ��b«x6!&Q���
� ��g{�΄7�wt���b�H~����i+�3%�Q;��X���sz�S<E �w+�_f�py���@aK=$� ��5j��J��	���a�V�2����|�a�X��Jzu��X9�}i�V�M��v�g2�K��p�S�^�ҜN�i7��d����;y_n^�����!������!3�� ��x, -�(�G>�	?���~ǚ�78:! �\���0�8c����w��]�P���^E;�E�$�+&G`XT�^L��![1
�!���C�M h�t�;v#�~S��@ .��I`��#%�=`��i����Dɝ4�>�rΕ�.>�Gb�]��óNw�r<�4Ϝ�2�������������6-�T�����S=����	��C%��OkD�}-j�`�5г�a�̌�<-:��g��B��8ؐ���r0*�^�Ċ~�QȀ��_��v��:i��\������������99Z���t���s�4���iK����hxI�S[-K��$�
��R�����/�V#}�d��Ԟ�v�wsv�3[���Co��˺m:�S����~Q�+���[����unU.�@NP����JM��ͮ@;�J��}�����=a��&��f�3��9bv���m� ��L>/��swS�'�c7���G�f����&F�%Lu����v8�A��CYK{�I��g��F3�� 	"�u������x�� $�G�z>Z��ɰ��jA�6J �ӱ�d|�<�Z��c	�������'����2��:(}3ш4���CP��62A3���E�-��q�3��d>QXVh@�@��F�K�o��?N�M�YPpe0	`����h0�߰0:�Q�^�O>�h�&a��Q,e�.�4���O�Y�*�f�J����PRp���N����P�L�Y�$B��y5�%ܓf�i���=��?^�ץ%ǎfR�6���j�
X׈�U}��u�+>M������l�L-|o�	l�����g�I~��6	�ƺ�5˪3�������ԀH0������w�*�,�a�C/�+�w�� Q�U-��w����p��Ӡ���t�%r�n�=��uI��r��ڇ���D �h����+����A{-�~��U %��T��hB�S��!�|��"�gm�azy)4ɞ��*�f�ƽ ��r�.�0�pe+8����b��zu�z:x�b��{u��r[��jk�oe� ���_U�b^�d%����61��7b05�1N�g�������S�J�v� ����g�=*6h-!���������'�.�l?�����?���N!
iue��po�w2Y�>���a[^�hT�d&sR��lB�ȧ� ��'��Q�c�S �����#
Ni��#:�l����\�}'y�d� )\�����ݤ,t���2��1�^���)A.l��
���UR���(8������b��zqV��I)�8И�'����u�f#���p(��S]���hI��kE ��u� �=-^Xb�EQ&\ɂ�9
�� ��q���PQ����eHJ��q�>dJQ�Ӂ�+,�z�8Dt�/�d cX�Ͳ�x�5���q����?跴��zJ��m ��]�*8t�`}�JsS�W�ju�q�<��$.{~��o����w�?�G@`q~�;�{�:,�h���^�-C��b�B�< M���h��Ø��O�O'�>�zQO
�|�"#K5��1E�C��*��ů�f��q�Ѿ3a;zG���yDwБi]/�V�ڭ�\�����~?��K}���� ���E�|7�hH/�8���.����]��;뫦�`s�V4�]EA��hHzx#��&��`�����D�ܜ
,U��W:8�{�]���38�TU�d>>�y��b�$(</a��-'��(YOXl<�_}}�q���5�T|����ER�l��r㩹7��3�D���i����d"͈ՙ&�^v����g�Dw})��g e.���d��x�\0{��v�xZ� �OL�uF�H��0y�\��l�Ȃv�����V�p7T�� [���5{�t���"Y�M3�>
~����|x�^P����3�'{(����^��8�<�2EU͡�)����� �|(|���n��0М��U�{��.��+��A"
i�G�B-ஒ��8��p��7�jm���?�Ϲ�����[�ħsa��+}���
�-/�V��c�L����`qu�C~7�*0�$��.@��7f�?�O�n�����Y���:�[���X���������s�[@؇����	��C���o$���N�-V [pd<���}�[�x3��>M߻��dQ�K���0�.�b_�~�2�"����F���}gތʽ/�H��v=���l���� {� P/Uiף �����	P��ۏ��.�8��E����]Y��h+q���w��/#�����?@������������mMBy��Z�����F��K=�q4��^=� ,)� _V���?��;z�Ԥ�?QsZ�00~��
�咼��?k 2�A���$�{���~���l���[�
)�c�?��{��6��kh��K\�0� �4�����&Μ|��+�����J��J����P�#��u����L<��<P��x��(l��wi1嬜-�)i�A����v��V����h��˭�*xl=S�;Ҏ��cUmt�W��JU���[� ������!Q���v��e�iS�e��zpLl�j��¬4.>���=���hO�-t1�j���;^H-}(����k2&{���������P++r'e�F=��8*���w�6�F�N5�m�V�_�ُS�\�ϛ��r�z������$x��ċwmK��[�p��L����ݻ�]�s��C�a��iSZ}�E�O+:oz6��9�&H5{oX
p�����/��5v"x��>�e`��7SSt��(�o1�ї3�n[]�D����*���H~��ϲ��ϧ�� |U�!�%�ǡYۍ.���yn�Lw����xe~Uw�G�e'��˩�H����f��Q8^��"c&c�gyΛ���c�hgY�i���!�3Y �n��~E��$�06��0[�"����E �1���ڪ+�xO�p�%����M^qކ%�)\��w<J\�n�w���	�W��)5ԗ����K�2�B̎ ��P+ߦdV�'��}/⋻�P�)���ZJ��C����aSՖ}c�l�O�ǨZKɷ��jrfS���<~���}/���ϑ�uQ�>*��ΟH��5d����bRR�,RR8kUۘS?za��L�8�h�
N��w}z55�Ng��d/��\�@f�ШITe�P������n��Ȼ)� 9�of��X>��E�؞:Z����<*]�~s}�|7W�j��	��zV�6�> $Z��[薋~(�p�i�U���l����=}��D��;�<t�A�\�VY�Ӳ�7f���!��>�Eh��NKW{J�������gf??����FŞ\��W��ۓt��<б�
�8��>Q�V��	VE�fzE��!������$8׭o,�jX>p�X/ѲC%�J�����U�*�2I���	�]7��?�|twG �ج�z_9�ǎg2fY]��t�r��1����L��k�=�d&�u�P��\�J���y]����q����(���tw���V~�W���f�#i��Tpdd.�����om��M�����4��
��6z�J�0u\<t��O��lmK<c�߭�����(��q�P\	�g+W��"�P���X����#1��)��x2>Ńm�9�ĭH?s"��a(�LF��~���y?vf@4��un����1Y�x}*S��L�''�����!����A�
�F�V;߯��G@����b���� v��^�C�Z��nB�-&��>�H3��P)u	�����a��s�RK��t�	Rms=ˮZ"
��?���jjs���5�I�a���F���q���d�A~��� �N���giQ[������;v�S'��or���U�A8Ɍ�-�=�X���?Z(�x�%i-*���y!� y,[q6)��X"=����X���q8v�<Z݊���/��y������	%�>3���Q��+�n���%�C����w�]b�����+$j�����r�uu�
EQ+��5��F�qَԽ��1�>����E�_ib�k:魏���_�@�t�/~e(k!�{G��ä���iP�WVWI���y���G/��ٝ�v7F�T�=��UM�%AhJ͂���s�W���>!�T�L������HN
���w{��9ك��NHM��>R�9*�o>�i!m6�k��>����>���j�(��v���W�s�L�A��AM~�/����W�r3�يi���r��#�̢xS�WF ����8b-����u<͕��<P���Q�Sٺx[k���8MI���i�j��?�Uq��Gl�s0,�ʺw�GF^��J���A�hs�FSP�8@��\ǭؚ��k��&	D	��W�f�g��9*x�����f<���8��fc�N���ji1������O|�s�滹���q2���N�"����\�zJd���dD�* .5���,V@�.���?����2�\H�\����SRT'=�啕�^6�ϗ7l��!���9TV?r��&[��Gw���u�g���V�}�,L�^/=�jفv^�Щ%x��d�m���D��̭��ܾYVV�����Z M�5M?��^u�6�����~�Y�*��5d�HF#�\�>>���V��L#��4w�lIP�{��v�	���� 	��W":?�D$l���w�a2��sTO��X�f\Чz�tA���^#���-͂�Fr��s�[��%o�`4`e3����Y��J��,��z���t��02*�}���qt�{�Hg����q�o�]y�É��P����]W��ĴZ�c����nGf�<���}���H�_#bw�(M]/�yr�d��I�U��l�sx����tnH�۴m���ї�!9=y�;��s�������a��R�Ob�Aq��Y5>�y;��VnX�����6�$al����&�x�r)&�0蠥�V���SԞ]�B��ʼ���ԶU��|,��E�$��c��KV,b}1�c�$i�[�zQa�<���Ȯ���~��GI=�n�HӲ3O�K�����p����dio
��4�Lu�F����������]���9ţ.�� �P�I =�"�,��l�z�,�v���a%��43oe@$<C��-�V�3%�����%�Ʋ���֤��Ws5����;�W�y����|�u�8әܻ�ժ�E ��Nkd�j�nƖC{5���wM��`V�H+aF�п�y�vva�GKC%��ﯼ�a����T�KA�)�pF�� snC�*�6�hr��K�����9Q���(�1��,2+iH���
��͒��9u�FѠCr[����it���B
<,۪�RpJZ�W�)�n����c���K64��f!%��o�2>�`���h&f�7cG���N�w)T�{�M0,� "DENw�s��l���߮@�Ϻ�+5S��d%�I��>5L�w\3��F��]�RX�$ƭ�l���P�tLgM}$�Jz����M��"��TGB�6cpP�d�ShEq��.�����
�B��Z��gtnkc���Y-U�����n�*���o��_��U�I�x�H  ^�J7T�Si�k�۪����ZΗ��ŧ�!��9����k-�v�t*��=�!!Q����9|%���C� "����B�K���6��-��5���������bn��7�9�'?t�<Jt����\SD}�iV�48�vZ�F_��WM'ڮ���8�3��p-c�)�-��D�X���L+/t�}��['s5�qy7ݷ_�ĝ��ʌ/�JV��U܉�ۋ�E�{�|�9�`�pbb')�3sL��Ƭ����@,{������_j����(��:F���g���7
�@+���y
�`4�e
}�r���k�)�e����f($��oBf<h���ڪ�곅�\YZ+�}f-ڔ��w�C��i��N�W��W�v��Xw�q�à�XOz������1##�����,}���@����~��6��ʙ�;���.��?�MZ�7A�	�T��H������X�5�U������?������44ߨ����\UD]�г�UIB��֟[��!��y��*���]�q��nG�s�32�C��C�����ed$���K�8W�W��㎵k�^��j�ɭ��	��ThD�e��[�ݎ��^�)�����~�{;bl&7k�߉RT>��pR��(֎�z�m �;�[�+�\�4D���Q�0m4ꃏs��,�Q�R�-���}��n���g�����؄w�=���d���E�7[���?�k�_���A�4~��Ay��">��Jܰ�v��]�[i�j͚�`�C��[��|墘�bMO�ϥ"5�_,�ln��������u��RI�0��^Z��;C�y{����7��ƌ�<���!���W���VG��[I��C���/M@�AKG�_%Ռ����w�F�͔���/�tPFg��|�͓/f�>�̷Y�i�i�e
��K�-��L�(E�����y7E�s�~@���������p�P-�pyW����]�+
5i���e�Fo{7����0�LO���C���=���/N�4�j���o����@z���˳��̲���jKB��3-*e���T Ŏ��Y�:g��;�VG9DS(����$c^g��Lߦ�#�3d��%{�F����*��#"l����D�����s�g�J�Y꾧��l�ˀ�{R��Ҏ<��sC�K��(����[Y���2���O+��V(����ɻ��Z��� Y���g%6�\�y��hZ.6�y~����xGU�W˪���js�3�׼���A]�>���p�p�N���Ե^��"�;Ȁ�/��.` ./@K���,�}��=��k뢝w�����!���\ܞz�&Ü�.��ee�O(Vsg���e�7�_8��T�����Y����bl��b,70Gs��(�~�ǜ���j�+��e]��H3"��=՝av�܅iT2�ǈ���f���b�djR�/v��ǭ����v1B��U��jm���\mW����Օ� 4tv@�`��Z�i��c�j{G�΁S���pFƸ�op�z��1I/QYmҮD���Y�T�Q��c�����v��������B��;�0��jsc���(h[䜙�r��
���$����Ò����5��)�'����]s3�����
5[4�����A���Կ���:�O�H�F-�a�DV'Y��
,M��2���4��*7�Ѿ�村�{P���S?n�Mq"n;YFB$e[ꡂ��!�͑M���E�{h�̬k}�c��n?���e
�9��h�_�p5JY�
������j�U��<8�-p^�no�̹5E�T�r�<�3�>]cg�2k�*�JuY&������O{nD��Kq?b���3-	=l�7,����(e?:��;x��nL�pQ��W���o�p����,�R����5�F�8M�4܂��	��A��U��ՄJ�ѽ�n!,�I��Lm�i]	�\����������&t�e?�r���KMP�ʳ�J�ѲW�o�d�L0��yD������0z��m�����*�)�&=��,#�*�T��~uŪ;8ay/�MF�Ⳡ��#p�;��ʥ-��V~u�\�ի4ř�|c�/2�1��̫�|�UL��n����P����i-��s��Q�}����݈[#xaf�j��6��aI�'Ǭ���Z���hwp�Lnoo��W��h�֏��Ip�OP�U�m�h��i�8��īs���R��������s���d�m�c����t{�;�z�A�:�~(�/���P���|I�*�c�'}ZS��N��F�N�z#�v��ɺ�[�D���[j?���~uM�地o�w]��HIuE�幫6Pןˍ����Xz
syg��x��F�D-r�r�r[䙙�-�G�
H�z=X����;[o�ڬ���֨��6C��[��BŌ��対�_�lK���F/0��VD�R�lq�~�a���X������G�栧FL��yx��HFG�
ň[�ʇ�q��TQCx��W��┨���12��tW|.�PT��?���p|����G��8j�;	�������TiۙG_�s_�u�&Dcmw�fp�|f�c��6�'���Xo�)FEE�IEPpی����0a�u�AM���:3*�
y0�Ø�ᩣ�0>D�9�|�U�������⭟':`?��P3"�u�8E���[�����ߎ���˕_
+8i_�EUX�c�}uNk�:3D�<{6���jB�ִ�TcU���>7���4���/�
�b�Ep��qثdw��!���~DG��M�&�SnT�T���9�������I�Wr���K՗��x)�}XG�Z)�WjJ��;�n�{�z�p�`n���Fj�{�ݳ/�+����5ii$��8n��x3�}D�sDV�.��;�r�l��M��QN~kC=D-���ه�cx}���l���q\#i4s������&�1�B׋KUȂo���A�_*�����1�2��˯�߮��Ti����yR�����e�ffy泵�崴&���婗�"����v�}j��믬d{a�[.��צ`7�Eb5��d+ڷNMv�PQ{(T{��o��ռ�G$�ITR��=�b��.*���Y)�7���S�q�Gf�"#J�����ѐĲP���#<��~�/�K:��/��=��]���%s,�)�e��\�D�����m�
w!9�@��Ӿt_K���s8�q�*��#wN�)~⑗w����4l$�/7�b�S]\m��nY������y�B&��Po���,�����jP��`�����K��c�-�G	w�&�;�g�)�TCf4��=��^O�45L\�V�����Zn�#w����!	ĬFu:�"-�HSh�`��3 ����;����ZW^Ub��y�=�u��a�k���7p�����?��W�E���h��{A�����M(�r��6�^j��sOn$��n
;wJ��g�$$��|�gN��w3|� 1ЙH=0�ᩜm����'1�wNo"�V��5����ō��e���B���Wz�"�'�ѹė�Q��ѝ�ոR�s�l��ֹ��kWD�NQ߽n��-�s*p������z�y7�hw*�Atb	G�����X��Լ��R��Oj�'�v*npO�V|t5)�����Tu-}hߋ�%t:��h{��qM��G���������K,����B��\���ќ��
��Zd<�36ϗם��.�=f��+�~W2g� 鼓�9��a�t�m�J�t��Ŷ'xD<+)�n6�SBc��!BEW�)I��n���=�Q-	O��}b�(IG�m*(�VT�y�����A�vM<�:�]r��ǈT9����?Od��"��8��
k7���ɓ�Dy���5.cn�)����G;'�/�t����\62/>~��J�'��%�Ԓ����RP����)_�4��6	������ �:>��b��:Zuu�����Z~h/��mg+g��[����\%m)�+"l��8Li�*�MS�{ʞ���D�v��}�O�����	�!\^ݝ������ ����3�����}����?�+9���{d<��O��c��q��D� ��Bhs7|=.)����f�e��r96�A#���O�N��_�u�B9|��~�!�ֹ�T�3�b�g9�(��_"΋�e��8�ً}�]��w<��q�s1��-�G�g��[c��;L��XA��6�q���|w������k)��5)��Rk��X�w����`'�Ks�dv�X2����;o� }Ҧy�v�\��Z����xN��uJ���.���2e)��e;���7��T�0<��s�u�!ꈃ�HƢ�+�[w/�E���ܕ�4H�sn�)��f�qi��B��Գ��d��!�@�n�tWe"��+Gl���e�A��1�8�実O��#��`���2��U]vK���G�� �G�h`@;&{`3����Q���Lf>2~ei-Go�G�o5�fت
Xx�Y*�V�k��!���a/q����Gs�r��3,�nT���uxߛ�w�f8��!;I~�{?r�ǆ�2�����.���)�T5"�Nh[M�%�1!��`��*;6��e��_朴��S����ܟ�8xی)I	���]��G����i��-{�bMJM��/�ǔL��uT��k�;&�����V�͹��m�Y���@��HvsFÁ�iΥ>���$��8����Z/t�)a��B�������YX���ERk��40�}�-�[!�!8l'��shJtz&��m`�MiA�PmE�juJz�c#a��Xr{�D����4f�nI�˫�C�p�����N.'��5Q��>{����p����$�H��Uc���� ل�m�=�\�j���������h�iW�}dDP�^���@(��[y\>]?�>+����l �=�A416�����K 'J��A,�S}̑���ӆa��+���<W%��.y�b��CZqGٕ܏��7뺐i���K���OU�����)o�\� �����GI�r�(�ö��y����d��'�п���+�4=����O�	s4X���W.7���?�z��O���KQ�ud�����2;-�%>6oג���=E[s� p�#��
/�d��6R�'�j@��%M`�&��C�,V���g��j�K�u���n�����s��
�c���v���J�d�O�h�NT���n{�Sf�;��xd47��E�dm��[tK��}����p,�k�$���8�:vDc�z��s|xI��/�3랬2���O���o#�s�uW�L��0yp:>��'lJk&X�2�`�z�5n�Ѐ^��+�G�(J�^v��-v��@���z��]�V奷���e�4���.����nbqƯ��J%�;~��܎*6������k[V�����Ŧ_ ��y�B
�v���K���)���Y�Pyp��U(�{N��X���Z��8{�h�!j^.�9gB����x>���,!.=K0ٻe�BD��bߓr_����
Gf�x������2�(D-�Vu�PF�qi��{�#����E�x�#���,�)o�+G�������=�n?;�!�/�(U�t����a��y�Lpj���Mr����9v�НLD�ˀ<s-�� h�y}ڽ5ö���&<�/u�9}�h�rw:����7,\�h��]/|�lQ�p���c���E,��_TO�����9�G}�z@J̚5�僡C�%A�WC��Kn�����&�e�oMJş��J*r˓.ɱ3ub�d����LT��=��1>��?� 8��~�FS� ��8+P��M��G�� ���� ��|���e�q�� Ũ�[Y�}�W��k�r��C�(-LpԾM��fӨ��.0Zb�W�?�#�-�~��!@��~P*�jT����[�P��Y��X��2�:A2�Kj?�%����`�G7�՚�gߚiA�s��ZZA�w��ȿrW{�{b��.5R���x�%@��=�޽��
T�(Ʉ1B��h���#�^��o��TX!�L�j�W�1	��
��:��e���"�0�H'(����Y\KP��+�(��w�)(=-ٟ�P¥U�m���b����]�ټp������|�j����Ҍ̵�ag�z�%6��G�&-o5��Ԓu[ܾǎf�����W7,�ӕ��f�R�_����
y�'U�/��ˍ��j����oJf}A����$��&@R'���T�n���+34[EIK���J��-E��\*��o+�������배'#�������9��K_�W,ki���3�۸r�ƾo��{Nܕ�-��0آ�(K}�
R�5L���eKe�W�L=��4L_��O����fCe�������3M�6��Ws+)�_�Xyϴ�%nh�-u������D��?2�	����Q&��y�{�rs��t����&{�|�o�(�ݱ�8�m�?<9��xq�sV(h}҆?�;�2ͽ$L�33�9@��:�|�`����rĝ�S�	�ǜ�hAV���">y�@\���!�%��W?�+���	�I��N�K��r4�����#ӌkA�6p
$��R��=�`��a�$Q�����"�"���u��`���z8M	��u��W(�����{E�n�Z���N�J�ˎj�����`	9a�(ժN)�����*<4!�S���D��&���ٽ�̭�`�b)�{S{Y��N�X"!}$�-��wV}YǰD�{S�ͅQ4q�W�8*�&O$Qێ��½U7�+�dp�Y�-( ���������,��\��m)���j����w~]z;��e���w/� �,�(��md}��N�&��o��sg�� ח�2�~Y�y
s��gX��je�ϴ/��k��v.�TT�j�@�>r�B�?7�t��������:��V�I��]�1ޫE�b �͍����cMw1��m�Q��-�h�〉�,~ADɂ�ߺ��+11��Z �y*�� Of�e1����Է���N��������:� ��� ��p�����#�Co�.ԫ�=�T�6�i��	(��[k�Z&�����
�|s�, W�iU��r�Y��}�&㌹�[n��`%MI�`=�����m3�U\�lJ���|~��b��A�)�#� �n�P)���;t�F�I@7j���%�x�AZq�k�p4�%��ƿA~�֟��T7��ꏅf�w� ����/DcTlj@��f�-����
~���+۠
�{gxF8����gb�h���g�C5N��R!�
����C�C��� ��݀������?�=�2ni(8IѦ�\�[��� F�
I*����������C�?|���@Y�U�8��uHk3�_��N�Y���e�e��E�0J���{�[3�U1 ��2���Z�
��xw��_d�t�b�@7�j���7�`ʣ
ʗ`���6�XGIF�����@ɎU0aoϞ^��u�h�S�x�� �a�b`H=3�k�sG��	L���;���l�5u���غv)���� ���Ji�����W�p�&D�>l<H�V`t���d�d{�ǅ�I/�)�(t����Q�¤���ΰ�u_8��NbU��ȣ�k:[�y�Wm`@�X �����d ����쏍{43L�E�u�<����Nr"�t=���"Ey�Z3P-��=q��_�*����������M��"�U�P��O�w�f������/u�RFт-x�ڤny)�Ufb�?�c��<��f�N��w����E�ƺ�������g�v5���Q�5�Ƙ�� ��@m^,#W�8�c��&B��|��%�n8���t����O�
�]g*�Z֬��Z	��C ��*��yξ�s�`���+��C,��0'����.g� �_�f7\�'�S���t��f>7W�2���2 aS1}}+H�^x�'�]z�_t�t��Yjͩ�ۿ�v��_?#-(���3gz���E&�k������QU0n��~nK4����^����uK7Y�T���ղ�/9v3j� ɹN ��S
n��g	F]��Oc�B �Dke���X�,�W���d9�36w��e%i�M�5�C��4�Q���ųJD�()j�Quٸrsj��̛}��������Ćо�g<�e��1�)V��C��ke�R���a*�a�}o"�^F}����4Y�Je8���@?-��7|�^������F��oH������ӿvEN��'t?���jrJ ���LT���jeF�Y��Y0��?cPr�W��\v������l	�}x����J�\�������^�~o9�|��}* ��������y�^;yah����Z�_h:S�R13����ݣ{��S���>��-�	3��G��j�L����̫�s1=���}�K Ϙ=T���t䯒�"n��B�
-��e��~��s��6}*�
���d�)˽�a'm�$>�+^GD��C�N�Ձ�/�c��2�	8�B8����-霉XPA�y�-�P�=i2��]�Աǭ~���K\kt�G3^�O�
��e�|�R9�q�T���ݽɒ��r���J�Q�V�Κ&u�jrH�]��jt��O��֮���L�T>�M��4�Fv��$K%M}����!>��ƛ*�0w슬��a�)J=و����@�q�ɥ�@<�^Wz�Ϧ4�5NW�<71Ơ�RmI<��[�k���b(���@q�}|��8�&C�c^�>3R�빞jd��mN�}����# ��۾_ѭ�؜��Ƚp�$�Q�?>od��ʚMz�C����$2�`�rA_���Z����p������~my��m�쟿��'XT��^c�3%�?z�,�:�CY9@?M�CS�[7T#�@iZ��c��C��vS���v nr*m:�J
 ��=�s J�����*?��ϜME��~+4^'h��/��8��>�|@/���qS��:2��E<bg����"���Z�5���b\i���37}aw@`��R��"�,�R��y)�	��4�#���1�[jE�J1ڛ�{�-�𴯯�O�Akm����ڄ�w�/�K�g!��2ߜJ5�}����-�Z��C�ѿ�[>Pa��y��K��.��ps�«}���5����u?1�1��S��l��&w���~����{��4j:�f�I�x��ev<���;�.T*	���_
���Lߊ )�tʲ���yM(D�t�$M�<e�H��ؤ�ͷ�_�y����;D��_ �����t�_��\��}�w5(T�SO��bH�Mk�� '��8'�M�J ���U�����J5�yw7�H�!�a�Q��,�̤O�p�]�E�^��\ޯ���d�a()�^"!�^v��� ϻEn�^Ϯ�����y�4LT��9՘�;�6��/2o���һF�f`E]���K6���A2��@&r3����JaF-@�%���������H� ��z{�s�v+��%	R 1��{����g\�CSSo�C�h%!Bz�f ����E����(\߄I�<��3��P+n+����T!g��WB��2- �ͯ�>��]G�ƭ�ը�P?�`)�ǣ؋tE�["ń
`x)�_��$��ME��>S>�:�ð��Nwۂ;����{淗�#6������G��L@i����7�{�T�m��d�}�C��8YMw.���d�T���� U��
��������:�7�-l�_�ս�&S�j|��B�w�
.�*�ꨴ_��m0FE`��W��o��W3�RWj��ރ�T����'L%��ΰ"��ali�I�o��8%�h4 �L��sI��(��d�'�K�]�x��`Cm��!���V�N��4moY��d4Y��^��-�A?Há���9����>+|6m�.����H�Q+�Jm���,X����X��w�/�eZz�����)������R�ث��dS*��^�	���8F��q�R!�O����\7�}쑟�}Y6 �6�}u768'�K�bނ'Q�j4�ڙ*��Jt����g�e&�>A(��aW�޻8��"?�h��9�B́�{IZ����K(��O�o�苑��u������ͷՑ�G&BM��=�lզ�1���0_񱣸��W��W�a �Y�gh�d��i��1Qo#
�۠��������HÚ���Cx�����n�HQ^���hM5@����X��FN�W5d��tnG ς���#��$�O��7%���'����)s�b���!��f\��0]�A�-˛?ZI��bݮ�K���C���7�(a��?�|#��jO�ǫ}�p����� QD�?��o}��S�ܾʥ��UVG�y�*OL�o�X����]�IQ����H!1�T֛�iL*S6@�xbQ
TZm����V�61鿹�b\y"��&��0T⋽� G�U��^����呂�E��� SA4��ĉxxڬ�7=	�I�����j?T�藬!�`���:g�S��-��)�9L~��� H ��$t�H� ��@�H�������z�t�qF����/�my/-���*�:���S�}�=N��'*x�����ь�K6^:�}��o)<a�_8�'�z���hX'�O�q?�r���#�&=�����o�;�/�W�RU�䡛���롍
A;�L{?�\�2K���PRR�w����s�� {��!���R���7��A�S�է����hUsi��w�&__U;��C�6��%-��O}vu�9q��S�f����������� ^�5⏬���&�z��%�8��l�3�K�5~��`�	�f6�H�fW�ȟ~M�H*��mcMu?Q�V�!Y��d��5�I�tp~%��,����Y�gB�0_>��t�]����ւ:O���J���T�uTT��=>��(��4���H���Cw��)(�)����%�Cא�H������k���5.�̽�<�~���9g<�S�|P	i����!�tHw�$�M�y���1��f���[��$JN�ޙ�)H�~%8c9<�s����0Y�j=���%���ɷ��"��U�(�Y:
z5}���Kj�����jZJ� SXz%�U-VhI����3+�5.D��G�I�D��Y:Rl?)m��k���;��	w�Hk��>�����u�aD�,y��,�� `x^�^&����7C�!]��+G�bH�m�`E_;��j��ύ|}fa���wD��O!'c����Qw<3с����h����R��﫣2xE����AhJ�e���_�в��J~z�"�'o���͗�~�@�>b^jg���84�����s(Ƙ�	��T��M����#���X$.�3[��������ܖ�S�'4�މ�6l)�HQr�
�����1Be��]�ݔ�[>�ۑ�Q��Dh����6��<���RU�oy���a��85��H*}�+�@y�&�*g:#]'�n<��iw��~]<�g<>��"e����Z~���o����x��Q��TFN��-�����.�ȭ����L�ˉ ���tI|���]�!!��C{[|���&F��W�	���.�m����[fo�^���<؈\�g���|�ga@��g*�r�'/����]�sF:1;CN������
���JO*Oܠ5nd��6��劁���ɜ3�4�.���`�3��w�L�����܁�	��3�(�kG˻�ytb��s`i���V1:�v0�[�P�7��U��c�T���d�?�����^@��X���4gs�����3��RR��\�����o�+�ʢBWOy������5%RDF���Q�Y�A�V�<(�N���#����Q�0�չ	� Nr'�Z��3Yb��OM����%L♓�Usk�����f(忛��TS��M��[=�w�?3�������_�x�l}��ݒ�����H�M��_�_n^O�OI��M��D=�k�fR���K�]�h���fݦ�`�s�8�C���~��4jD,� h��7$�\��u�dg���a������t%.J�/w���9�(#W�\�F��bm�MPJ�`ة�c��'�'3�e����Kw_v�M?,��3C-���1y]�xY����~�n�J�|FL��=
vݮ�&e�/��)�C�V�g�
{"H�a��w��2͂>�MV��::�%�����&8����·�Q�z������ܐ������wl�����|��cZ��rvhk���L;�S�q�(�T̐�ꭝ��'i�\m@$s�	�7�tϟ��qd=�3�~Е������6{uٽu%א���ZA$Y�\{u6R��S�^���~�i6M�#f�y�!e���wYaL%{z�c͵`��.rj9��ir�S9J7�<p/��^��0�F��i��H�3��g�tO8����G�	q�eC������S�����r�B�,O���2BOп@E���J�^�0�j�w(�X�R�V7m=D~���S���L�i�����h�شD���j��h��1�u���P� /q-����v{��)��h��rG����Mb�E�i���8W�o�Ј���O?u'���=^���/��!�%�a�������rx$	�=����r\f~O�Q�~ck���:��\
/�}��n�-�ɼG,�R�w�Ǣ�p�\TP���c�3���Tݐ��������=y����|^�`�x�ZkĒ�;��>j�k\�;>2� N=�y���苧�!d(OK�+�����;�M�"ڸ���C����1�_���DМK�<	%����s
��a��2��߳v�{�y���xؾ��d�~0cROZ�ӴN�i
+X����Cx<�D..�J��(��7� �:���J�+��c4�+�����J봓g��v#e��t�U맏<�ᷲ���6����-�5;6W�Q���)4dgp���5�΁�Et�Y�܄�����*�hа#g���tnQj[O���]��fvY����H��#mm3<U�K<�s�ng1���cn�wk,9��C�X?���~��K�a/�W���EO]�EzojɟG��~_��h�"��@WC���,�������%Z,�9)ɂVFy���Y�[!�=�(�}?���z��tjQ��J����~��5�5�~�EN񥮰�A��Ŏb�/l^�MΗ�w�lxOJ~Gm� b�)�q�_�=�4K��1*�!e�B�K�'��i`�.�q`��y[��Q8C��،�'�V�}
*�|Պ�[}�������S��К&#I��%����*�K�6��o�E+fn8���s|�F��r@,�d�}���_p��F�fH�,��q����k9�C�HwX�O��4�tC����7���W.�q~
9�e��gzi������	kT�7!�U�N>�ǟ-��AfzQ/u�^��6_`�_���dZ�� ��_CrCADwy��<��<kcdl��V��U��/~Z���o���$*r֋�������Z�Bd�o�o�-l��	���w/���s{f:Ѿ��´>��B�����2��K~���@ �ȵP"J��Ժ�-ϩR��!kv݆�H�l�T���n$ö��)������&T!���X�V���k�#:![�qO� 1�@.���c��T��KJ.���1�l�`�wW���k_�bاݰ�zW5$ˢj\�qm�m�����<�ܔ�w���WR� 	���iN��7l�2�k3�Y�S"�[���_�@���k�B3�S{K�r�`k�@�0M�/jkS>�Ǖ���azY1l�7Y俩˫]��m���1=}��� ��m�P�+*
옰d���I�޴���m��u�`R�K��.u2p��jW@Q~��wz�]�u3�e��jc@\Y��6��<+]q�<N�U�Y�H�m�~��J�����5�E�����8�-f(�;�%�I��(R=6�4[>��q*�'#�o/�﫡�J��g7��(^�΁�l�+kX�N�^��T�K��ի��u�R�IA�qE.P:i���3QG�q8���)�6�M��<�E+�Z�5$�X]�--7�Zر�������[3tB��ǋ^��#b K�{c�e�{�u0)�'��v������-����5�������6e�����K֎��켹ї{0?)]Hk�����uZ?����Ɯ[?�sh��z7��Y�vYܐ�N�.�ʂ5���}�n���2 -9�t��zր̅J���9!tdE`}�]e	E�˃��"�VL7��Zm�HzZN�f�WWH=�����~������l��Z�`�����#En뮤���/_K��t�0X��ƕ��`�pM�!�J�:ԩOf�F֠�8&�nD�V��#K޹�Ρ7�����m"�Zb5��EhnC�J	[O�e�:E�M{�2�?#����}c��:�	z+� G�����U�?���@I�s6���>;3�W=�u���$d8����L�c\�i��[���M��hw��ܣ�s����'�>Hp�����y�O
��+[���d���q�7�A���:fP�/�{􀮯�|,��%k��f8��d����.��8!���ۘA���,D��q��f(�� z4Gր-T���V�� DY�lB}9�por��Qt!@^�g�b6��f ~��&֜��P�5E�_�Vh(@��/���X��W�iv�n/�a�q���%9H�����,���~������˳�ź�YJ�8M0�g��ǀ��iE�&�f����f�OJ���A�����ĵ�>�z�J�c�Y3��*S@l{�>�g��K�s-�)���T_[WI���k�b��w5��:�vG+P57�:�6�ŔZ����Nkⴼ2"$�ER,7v�+�5�"�I��8����N���!u��yEk��WO������?��}oO�|;�<)�w����9��� �������n%.���)aI��~�D�$�#�Ks�����$��ë~F���5���#>�>n�h�)9@ҙ�ȓ[�feH*�ZN0� >��
A�4œ2^���o��N.��Gj�a�b]�@�5��iύk[�̆��r���ٯI��i�CT�hw<�T{B�P�Qq�����FHԺ�Ȃے3�wR\ .�ص��a�J���Xi��緥`��;���8��j�ђ��I?l	�]��w~�����<�ne�&�� �!�g�!r��
���U[�r�[.�5�X�\� ��:QD�C}-oNd.���A��9��%|8q�h���H���c���8e�B�Gd��<w��4ˀ+���ۊX�>鱥�~�W���QZ��b�
��4�O�ͯ+WI���a�.�ٍW.R�悻l딫#Cy�]�{ö1"d�xD ��c�LMAn��R���#
?��*8L��QC=��峇*&�pq*�y��U���&f�Ja2�{9g�}:w�Ѥ2���}���k�� >�c��2�?/��;�P�[��|^L	�hX�~��n�
�����'���t���i���ؠ��%o�s∽G�m6�*Y >�_ym��a7+�E��!	]��婾m�:�.K����
_S߲��'}}\��NR?�{�.v@M]����U��_n��D?b{�����YZm�U��2|�A�`Y�к&�dӞ��S�%W�oW!��ׁ�Hl�\��Ť e��CuV��R����s��q�]��A�8f��M�$��[��J���ot֌�+-oʹ�X��.}�^�x}ڍ��ߙQ���sM(�9W����y���S��:�w�N�DG��x��]ih@O?h�����#���5��G J�t�i{���~�v$i�\x���}�~C��
`K�16��g/�#�;!����ߓ����~������K�f��{B|�qh�k�/��
�3οκ ��2r� ]�+�0D�������S83����C�~n�?p�)��M<ǟ��u�A�¦��ـ	9���fm�f��+��`�%��Ȏ�o�}����D�^�#b?|�J~�DK�������ʆ�s��*�8���p�;�Y���zKg� ��w�������!`��!���t����0��b�oi���	Yڜ^��&�*�Π ��]z�؇u*�bf�����-�!��Ƚz�RP_�#�vG��Hw�������ŗKd�֬#j���'l�d�z�hH�g���|%�.&î�������zU�/d�t��F6=�+2�v	�⽪�JQ���[�vP��q�_����_�[~"��>oSRf�T��]��\��p�$'_	�HYJ�W\Qq��^����m�r:횚j�À���&vJ~<\~���pm�J`y�RSvODV�-���:oI���(�a�7�Zk�"7X�}�~��Ś�~�8��m���/��y��E]ӗc��C6�����M0��ع�Q��{��V1E_2�\�x�&�L�޻����grzz�Hâ�^�c��L��MN�%�p�@4^�*������D�{AT]%l�M#I�U�/^/O�óY�� i0�s��9�b�: H����2<�����F�j���H����і�"��͛�y��_��\� ���ϡ��\��e���5qh8�B���Y�	/�RxA�E]�/պ���W�E�L\D�V�T<6��GH�>��öXd����S͍�~��|��W����yK�^(T���L٥}];��g�6x�g��W���p���x�|��#�C@6�J�g�uS8z�=��m��}����,�G���$�<����{��J����$�_��)]/m��p	�.��z^�٦Z�PK������,��h�U�T~ɐg>!3����`��o��U&aK�v�\Z�,l岼5�^���*O�Aqq)i�߆l)�nV�"��x�kK*�YX�tã��F���������l�.����d��������^��~|����4��@��)2Q�����T3K��H�<�z�h����ߒ����KTr[qﾝ�]w���!?�-& /���ۿx^xn��S�a���p "՛��H�p�P�XDvZ[��d��[��*�]*������^�����7��8��#�B6}x��e_u��l�>K��?��-��g3�%P�o�]�7o�n�qgt��Ҡr*�[	UH"#K9�wLWx�ȼS����RΏ}��\w��:QͯE�����K{���$M��ȣ�Ջ������gU�(r�Z��lf���j=ʚ�2�s��#��ق�F�W�~.v�ڑ8�?L?����.8�:0D#�.��Q��$NY��O8���"7�'d�*��HVY?Uʒ�4k)7�9�Q���p�}�2�M/ ٷ��N��R�}l���!X����}�gp���aỸ�_���)WW��z/��ڀ"NH�<�C�7lFn5|�\ɍmmGq��8��N��%��i�U}V�L���|���sW��6�����݃t�~o�P�o����/�`~�-c��:I��$8��y"B��5��M�8����	�y9Ҷ�l[��ÃR|���z��4�񹽐��1oaB_إ�P��\�I�\O!�2"�w���Nr��-��,۟_�6ŻX��C��.��/����B��KK/��}v.�3��8���H��FҠ󍰾?f���}m�ێp�4��/�:P��w�F.�!;����P@��";���r1����˝�blt���f��a�3��3!ELŌ�(� @�~�&��렿q���&�q�9�i�ܴ��V�-���LnO^[�"b#���a�ڣ�	�� ��^{�A�_�PJ����g��R��B��M�֞Y[� �W��q6��+
�+�0�����P����������M ���֯W6��p����<*�^�dT	�A�H�F��PY����G��^�=⣜{�d���AV�Q�c~��u����b`��C��B��J4�"#�C�h��$���_��uV%���^�!v�'�?ЈpD�]Sԓ��jj��Y�!+�[���c�����طSY��0���6��5
��v[)���x���?�;MM��w���V����$I�Wd�O�?��8�!�����uk
N ��H���G�Y��-�xdwP$-��2�|l�����o�¥?�x
��\�HAEֹ&�vw��:_+�Dd����e��v~��P�o"�����é&_�B���~��N'LO*�֠$����8����_�]*�4�������YE�%O�f���7�jB�n2)^�Ԣ�!�?��z��Mt���j�cO#���D�Ǆ��}�}�����3�9��()�|i�}|������݆�N�fL����X/7�������??m9t����Mm��1~���9�򸲜Ԃ/f��-�jTz7J��{,X�[|�xQx�&��߽̓u[�{�_�S��z��}�p�����p6IW\��#6���߻��p�������г�F��wx*�/W������nY�����ag��/��z�WH����Bz���r�t��KY���pM�|���r�!��v�\��;���`�qn�K�yP�>�{:����3=�"L����M*����_c.�u����WK>z���K����zӗ<J�Ǒ.!m�S�����f���]���K��%�4ץ���w�U��ly�)��k��C��n��8��c)s{�=C���!G罭/BQ���w�����d��k�w,+d��N��h{u��v���	�V��Eӎ��f2�?���R&��3�B=���BV��ǧ0������Cu���v�3�ip5z�n�Q�$���C]0��X���̍����nđ��9�'�Ւ�e���7I�H�`,�=`�Z��?}N��V��3�9��um�
�"K�*Me!�q�잆�m'͇"���s�Ƹ�:\2]���x^�0��aw7A���:ڟӟ�rYq��K��CU���L��5\)�s��\h^���I��J����Q\a^����`��y3�+8NL`3k��hX=Y"�T>\|�	]�mG�:�ͩlE��4�1/AF���0v�ѝZ#ڠ�z*k��[�`Ζ���RZ�{�:Z9��;�%��!����L�RU�D���g󝉫g�S����P��զ[��Ǧ��6`�6�;�֔�԰��-V��g�4(
�*�5�c�T:z�y&�����O��ҭY6#k�GzZU�{��� �@g�cs܎�KJs�P�����U0n~�^$��#Y��:E��;�����*g�x�%G�S񐉆��)�5Ƈک��%�[f��o�e��-��VW�[x
�3�'_vY��T<���,�F��2_�R'o��$Sl`����s��r�`/�O��7:8),°���#��׆�{�"^~P����*j�Q�ꩦ�I�+!���P�wW���t%��Ab�j�!����#R7�͆T�z>>P�����I����\^V
�Z���;�R[�!֩W�w񇳝�����+��g2�b�};�7�"�&��
%��u^Ql/�����LՅ��~��1Trs�����E|OK]�	�1z8gZ�ʔj���K�E#���wc�/�k
S�Z*�|_�{�����Z�{Θ7 "�/��e�9吕���ul^\HK�C��&h+�W�+�o�Jr��\O3jĸI��{h�Y���'��l��P4\K���\�>G�a�[5���=��/����-΅�9k�io�E#��j7��w�_O���̽%���u�!��( Ѝ��p�[�׆~�@z��;�6EC�2r�?>UԜ� RV�6�?����Y�tO�E�-X����̱s��ϪX�b�@
�J��f��P�G���99&�l +�IYd�+�zZ�_�y���/�$o�t~kB>�R?��d&SKQQ��X��E�U�� ��ѥ1��5xٹ�p:�s��|���Bx�)y�L�����sQ�sp)ǻwb�R�3da���R�0�i�:O�s��4�Z)�Dr�����D�B[�/l
���杧�����P@>�J_�3�M�JJ� %60�/a���|���s�n) n:�+~�u�G ����O���k�⴯�p�((�l����6��?F�����B��g*�=�Akdr�^ ���^��|Xp�V�K~;.ּ�P"9`�s@==��~�D���u2�Ձ�3��P-����c�+����{yY������f�c9[�C,m['�ˌoۗ5z�/�����p0�<D=�j�*�է�μG�!ok��t��Y�l:jd�M��E��P=��`^r�E��8�C��0��z��Aϓ��5/ޟ���'�������| ��Y���#�Y���W#l'+Q����zy����n��i��.���8��Tr�Q�E�^+�
�@/���nWrug�T�W�Jl��c�Z��a���b8ln%�p��^DO��y�t͓�Om����\��Z'6ئ��o�<����8���\���x+Lݷ"���0����8��7����:�]�"�C��s�t���j'�1��R�5ڌ��EV,�4������0�]���]3q*S³�w���~��n�����Ğq��C�ݻ��>{���}��Bfs��}��Dd8�:�B�r�ڒ	���	F��]y�p	��z�i��8�����;x!�I��0�i�R�iQq����M���1���h���qI�A�4(�)�$���2& A��q;�|��9�a��9N��\�53W�/W��u��O��/~q$E�d�/M4;.����?�ˈ�� �=���ѿ��P��%�&�����f�4�18���)8���𓛸��MhI���q�w�Zlf��:^G�j�k�[�R�������+��ݝޓ%5�A��S	���y;n�;Y�r�E�9�!'�g}Ь,
q#���Z��w�����Ku�(겎$��٘��i{Dj�s&�'�k���?�w��:drA*5,� �nj:6_����@�B��N�y���S\��jT�������b.��2��c�q׶qv]!h����"uѤ]۹���Z5Zy���z%��_�����y�����9�6����#�1d<m��f*��� 'u{ �Xim��:�WC�h���d���P%Z��W��Ω�+}���YdE�E��l����V*�ߵ!�O����ӥ�K>���I���M#��hrs}�{��y.����W�M��O3=U$Dy}r٤�b���K��r�ёf2���c�G�\jэv�b�Β��"Ɉy(���+_R�]��1�H"�J�ڙ"v�|!�Dv�Q)e�?��y���IS'J�ܣc�j	�4N�Ms��;z�-q�8mA�࢖�͊��iÇ�L��7�W�ٞp�r̕�{ԛdP���Sa�̕'�pb��������]��s��=-P7���x	3�RLޓ�~���8���V��7L$�{�5Ar5A2���m�m�Faɀ0�*��ń2��	�K�'��3W���|�iqQ �&AgAA������d��.��X�R��4Z>&�|H�E�]�4ᙫ�tV@��^8.�NWq;�"^�����u�TI�k9`�n��!�g.�w�����I+X:V!0�-,H��Qq���S���+s�V�Ã�P��Z����wS�[�HX^a�
�_��ʝW���UY(��{6Y�����Ib|wf?����t���ތ��&���V��~	�����1�q�C|�0�"jC��UZ� 	K�)��ջ8���_����5�W���\��xi��ӺMB�G���v���	Έ��p��B,ȕ��@���N6f������}�h�k����Ǩ�ȢDΰ�b�`��[g������l��e�R�M��#���x������X���U��v{(�ڤ��=+W�u&\�w���QBh��d���CY�Fo�ͦ]<��=��N���,�q�;STa���y�s������J�I�4Y2OG%����/l,^�Z�^���2¿�1���«��h��6����>��l�l�gk^?�Xi��]�4�Jߛ��5�9?o� ���H���װ|�����jN꛵s�S$'!�[C�0D?��M�&3�J�(��8>��u���z.9���4G�d<�%CN���sXA�QPTV�g!
Gn���1�ż��r�C�����=�\��:瓺:iP���O������g���_��3�ӿ�zv�s}�VR�v�"�Q;Onj�T�Q1X ���� !�sxA�Md:nF����Ռ�R�Z)��}ﶴ���
��\��a�,EO>ਇ�*W&�{sz�B?���R��6c3���I�z�bu7Y�������t���Uq�Q��Ϫ�������YK����"�|2VA��� ڊ�6l���+�-v��o���0���A��}�A���ڕ�o\#=R���7��I�R� o�.h��2�<����$=�u�\���6����?��yoT���h\&_v�E�a3}�X���}55���T��u�Itˬ6I��}�h�~�3�%S����f�;j�����ٕ�qi��;��fm��_e��^��7�&��[�w�Hί5���}�����̕z�,Y��ci����8�Xÿ��莖p4�L{Vn�v������s�%pnB!:T(����f�np�FR��<�G���kX6�((g�'�����:���� ��ԁ WS�[[���h��a�;P�����_�вZ�B"oB��F�5��c���װ�c�݇l͈�X7>����8�ȁ�R�q�C������f�[��k���ˆ�8Q�z��rh;�eB��	�a:ڳ�F;7�.���>g����ןo�^C�l���v�`ZT�,	^��qǌ[bV��C�;١9�qlU����k\�$�ԇe����Ҕ��ԧW�
յ<���ff��<t��7�����C5����PS��wz�!*ULOg��,`p��޻��n����3�t��q~�y����׈����lYR�]\u���k� �VL��j� N��` �a���f.1�[�{C}#�����v���ʧ�a�@���k"Uo��A�8���ݜ��)��a���x%�	�IJ+�Y��Cx��z8�	�Qa�N ��¥�Vj�[O�e�-��8�6I�f	ѥ��g~��W�	X1���|$3�w�U�Ң1�#6�1j�1�q$=WRd$��0!9����V|��6? +�M�3�~z���ܥ6�>�5V����vW՛��C�)"�%bv��LPQ��[��J֤m�m�J���Ŋ��&�B}��UUV,E���]�s���0罾�����6Fb����+|Py}AT4p�9���'�����jP����+R�ˢ�?w������FK��lA&�dB���ɕ� �U���`����A��Ӈ�	�[K�����';f�-���Ũ���zf�h�Z�ߒ=�a4���uu�螯���D�cM�{��X����,��K���	�DƞPY_<q�ZP��]H�hߍ���%r44^�-����r�����Wvl�1Q2�5�O���K�X��}�|��E�
�]9�*~�;�/m$A�ܯ�s��|ٴ��Z�iP�Ϙ:�_�n�^e���j�����ݾ	�n�9]�MZs�y/�P��B[��l�0��`G���ӊS�W�-˒�
ş�Y@.6I'��A�FO�څ��^���T� �`�}I.]z�/(�����^Y���p�y"��u��P��~+�c%è
y�`� }�5tBs�L�#]@IӰ�����Q�&,�#�_2:nL����<ޅ�U�N��Y�~��!ω��@���c��4��.e~����`�]������������*���X4��K��on8�7<���6��'X����ԯ��߱�b?�6H�=�+�e#��btZN2��:�o[�����c�e4���f��9������zK�s�D/N�&dń�Kl=N
D�θ�7y]����.K�1k��r��b��^��i93��Xu��c��%b�0��M���ulr���!��|� QPXV|�j"Ӎ��`��^�4�)Y��L��O������\K��g�a,N �_�=�Ҷ����:�='v��VՃ���`�e|����&$d�质g�F�kf�<���8b^h����I.wJoѸ�D`~��[���������R�=N��uehi���9CR�0��I�2�w�^�X3�Y�m�	�/�\f�(����,�)/u��=���E�!�]�|��ޤ�_�Z�]�V3Z����Ia�a����^��g*�g\m'תP)yqO.���Z[k=�����S��ʅ���J���}��.��]�'�����z�ᬜ����G%���D���o����Sd3����2�"�9J�/e|��s���B2�z9���.p��X�E��ak� ϯ,Ȣ�������,����Bo�R��o8>��6�^��^��\�A�
3�}}�rYru)��<�Ru���s�i#A�~S�W�I��!b��������Z��+���� P����;w9��b�>F�Ŝ&i^�����W��e^���4�?�m-�-��[�r0k�ab�ޢ
�������G�'X��d�� et~��H��+2���i��D�ؐ��>3g�H>�G �۝ȓH����򍚻�D��ovR{���dֲ�bbB+���ԑ��24�À���7�,?W�7�+�,@�O���2v؟���ǎ�i��.������j7:|zH��H?�ܻc�=�2^�7X�K�;�qL��ʭ�z�G�ʧ��[��Wg1J��  ��-0��uI_������h�b�4�m� �ђ�cu�qi��ca��������j�S�O_p71�r/�1�x��m�"��7=G��,؎UK���]>C�y�~Ó���_N�w���2Om1@ A�v��gn�怄�>�h0��4ZB�%eK� i`'|Z�E��qL�[� � ���^9>�m�[�G���y�`��k��Ak��)���*YO_ �fw��)/{�y	�H��Mt<s��&�?�4~��.p��挅nL��̾�����1]R+ ��^ �n@y����Y���'v�=_��@kx�|R�Au���L�nqt����p��E����ppS �?|��,��}���
��XM���QT����_qB��1��:��5u>�ۀ��?�B�t�#;��
tM95@��'U�V�i:=�ٲ����6K�t�E��Fh�N��6K��ȳz�6���x7k'q�������D�K/��h �F�%�#_K�M�3R�0m��$�0�'���ɂ��2�E����@!F�8W���<u�w��lK#��	��[큇@��� vW 벒:��n����c�)A��g�O3��[���́�@68y�=�53�(��( R��B��m��dq]�on����z�p����C)9�Y��l��Z{`�f�{�[X�Fj��@��;D\�*vЁ�RH�����O؎� ��΋������}`V�FR	J�P@ ��Q���Y+z����c�h�# ΍�q	��i�\D�	zz��	�`�bH
�y��~إm��!�FA�#�\X�~�D!��,�T�tf�{C�@���������Q 2�p����q]5"һ1]jl���W%�x#��G�bRvì�U|�q<ewv;3�O�=�� ����.�VL�a��M�b��jl�X��Ѐ�l��9�`>�r�R�Ka�fh���1r*T=s^��"���I� �:퇨���T/Yp�s$3���\H]��N��J��s����v����J��>�>F�c��2�z��?�ktúK>6��tO��Gpw����c�zΐ�>6�|���@�奚�Ά�������+�w�D5?�s�\�� �p,]�IF	�Ë9��UxR-����{ CJ���,�[FO�Ѐ�}���I �4\��l��8�w�"�$nX���;�	4d,�V�z7^��M+M#d�zn��I�Pr��t}����BP� ��(˜�F� �x��d�+����t������כ"��<�f"�5]/'s �5E�D�������ɑ0��=�5?Y^����" (��|��|�LC�0 ���r�G_z�*��"��"���Td���F���].-����~w�W�! ���C�jFZ<�FJ������M�ο�&���P��N@zJ�^�Nz��Ao���6!ۼ^����!)��m�fd{����4��?�j��}�HWEG�?
�I�5��ij �~� >u���Ew��^6��uq�B���`�e��"��7s���>�x� .�ר�� )R����B��$��>"Ý� 0��Cl�E�_�������j��9�C%E��Ay0ɛ>ϫa�f�4R�*m5n�E)�o8�dV�1��i�ŷL~u>�0AQo�Sp�5�����&����?Uz]�������z:�E���os�)�q�/ ����b���s0S���ķ!o�ؒ���`:ɇ�ڲ�@x�E�~vW��Ğ5���u�-Iy����xa��Z	u�Q�����2;U�ƕ�����g���U��YK�k����+��RϬ��'�?[�l��"�>��N<�'��J}3�8��"#��N��!k�+��_���Ɓ�5=;�7q.��Gu�Y�N?�<� >�S����/4�;�cu4�\yY�C�� sK��+i\�BF���W͡���%�=�#��K�4ӡ
����`*���$�3 �_2��Je���C
M�s蛐l�g�ygV
�����O6$�ӑ���&�3DWxN��:a*���!�`>�b�!��A�@���&���饏�?w��0t&o���"� �3�|��%�~G9D�P�d��;�9�� ���k��U���	�`������ޛMG��y��F ��j�t!e�t||ɳ��@a U�Ò��!��/�l} IWے�3*w�Cj��ϫ���'�9Z���� ]}�nMm�/Q��9�5:�n&�LESAr�4�����mFރ&�N�V���P���|��=���}�']��W$
���]��%��"��cb��J�Wc���)�����GVKv�I:��Q�<�C�O�������p�l����0+�3�[��9�35�M�!W��M���-v$�d,���@?�"���$/��A�I�� ���@���0��Ϲ������y�A�N�������J��$`nѪvs��g��=)E����|R�B�񚷄ֵ��:�'�Y�C噸�-d7�|�� ����.��5�(/�+��I��}�?���|'p1�Z�l�n��q�<�����������z����6ʹ)%�.���j�+��5�&6q*�C����=[��))vP۝�Ԕ٢�n�}$<�ʘخ�"���~��ν��۽Iw� 	P�K��{]x�H��*��2$	���#	���l95/�L���Q���݂�`��^��D���@ <��[�v�qWGj��*IK���@����\���� ���h���nYЎxx���(L�xĳX�k"�
�ÏHYb�~�d|��ë�F�5�	�!��Bˠ�S`}+ W�������$��R�b� Ȁ!G�N�k5R�wZWZ�g_X����ٺ��_L��V�;!�/A�f&��_.���xjٛH̀<��ǃІ�b�^���8��S�q�����O�
�!7q^��S��~}|���ϒ����v�_^^��w��@N����'������>��+?�I��j7��/NV@꫻fѕ7ϒ��R/o�z�{ZV� �h} ���\���Yc8�d\{jTN+Kmӻ$���"�=uc|�\ 5�ӻ-�xg����ߞ@�m�*=���$�\vv%5�� I�O��	g ���y�8��"�??m�d��7R�� �wmj�C�ȿ*Ŗ�Q=yc;��@�a�KwqL���
�e=�Ժ��C��j�;z[�X�$�%!B}�S��-  �.0z�a�.f =��^��-�4�B���Y��_�j����v&Xaxg�{�k��mz�.����߼�Sz��4�5^�e�N��|
����[��%/���������*{�w���k�
�J�()��+!5H7(�t��*J0��%H��H݃�������/�%��<����9�:v�
�E>��`��:�|p��񫺋�'��k|jK�=A�tx0�Y���~b��^*jZ�CSS�G�6�/֊ 5A"�CM��Mc&U�<tϗk4�Rs��z|�d�^,�G�?
��zَ��G,�q��8�6칥)�6V.�[%�F�\����[�@X��*�իk(��k��R�}p� 9aTH��о��R�x���b���ܱ
�0�ڗ�Ap�q�7/�fN=ɍ2��3�<�
:Cb_(�]H@�{%�J8k���$� ��B��+�����\��ҵ����|Ќ̚����a	���/g��٬/L����K���M^�Ҵ�E㬢����!hy��V��������rїpr,7O���rj*�� ���7�Mg��8�4fK�4�׌�/����]Ys��$[[ȹ��+w����\.	*g����Y�ad��	k���B������A��~����.�F�K�U"���6J�ɥ�h���,��+[ˏ� w�D���k�y����0���Y��9�� 4o�
�Hb�z�<�PZe[S��F�4�%��k3�i=���l�`#�h 2ܵ&U�3=�����Yz��4�Ȏ���X��E"%TDn�yN�l��-���d�"G{0��W��'������4��@8�ö�"/��i�FJ�h�x���=rTp�h�Z�Z)�)i������}0� RW4�L��?J)���4��U�����(�B�)Z�Z�`$^7�i�	R������4w�~�"s:\���-���[��g��Y���K�{J�����1���7��]�ӊ;ߓ\s�tp$!o�ǵ΍1n�*�mEB��#�^�ڐ2*�q9�[PA��a�U-�-Jq�k}��,�cڻI�p��a��A�ݥ�7�k�2.��܀��z���t�e�x�h�u���J�,(X@�?#:�o=�\{�*�.��ʲ�D����T�`����̷����)���w?��kqK<u�dF�0M�<O��pd��S��چ^���A?����s���է]m��{��&,j���>�Hnj�(J>\-�|g�tt	�w��:���U�0������"���B_���n{��<5����'�ٵ$��yy��F�+��}u�����6��3���@��`rz,_��yf��P=0`X]��kj��Z��V���O�k�#P�j�e+9�.b�Ƞ����L���Z���9��|�tS���(��4cLO��9��?�*�mE-�ѹ���B�j|���`��a�1y��ޱ9���^�sVj;ƺ��|P�Z�,/�т['�?�P�V)�L�U��I�Z7�jsX	k� ^�{]\���	/���p�#X��>[�������6]"��`�������g�T����{���G���kn���3�ס3[�����继>���ꖥ3�1&zYS�J���&�OL�s�-*��0�S��Tp����`��#���o�j�Y:��x-2�����w��#"�����nj��b�uf�������9�J�w�.��x�Wzf����&��Zu���竤w.�a^�i����ବ�N�xs.��9��E��k�Zڙ4�l ���>�"
�xz
>@�Z��Øp�,���l◡����^ʠ�,\�e�uǶ�Mw� im�$��?@�_@,�w7RF|(��	��I�����|O�0:y8ͱ2��ri=2lg�6��s�����!�k;� gQ��T|�v��We��h�[�j�C��k����*�����D�D��ރ�*�q��
�UN�nh����
JP��̾{}�����"�j��s����-�vZ,-���Qj��_g�=ƞ���(�=��{#:��*�O�4��I�:P&v͡���\�	!~�7M�%V�R�V�!����_lL�nӲ[���S�~2ʲ���+�����#l?V��Y��{\4s�Zr���$S2��H����ܹ���r��>�����ˏ5��F��r�����i:*��bCu�-�L$��:��,���{�}Ò�����H�������Xz0�C1*�3��|(~w�����T��d;�'$|��6|�w��6�#Ԋ|hC��AW<k�hxt�exjnlڴ=M�]7j�
K���.?�ئ�:������v����pc.sG,��ˎ���>��Y��)q�`#S{�ڳ"V����/y0�j��f�?aZ�Щ�S�c 9��X����gǦUhGd�yi6�
��]��{_��f�zT�����0��m�{y�o	ݧ�%ʡe�zD�j��r���m�l�����|}�_x�gN&�C������RV��J������I����R�<j�{�J�R�s����U��Z~�QJ�����+槗!�����V-b�JqRt�C���Y��I������8���<q���B�䨶>.�|oR��Y��8��Ak��H�m&�qK=fم�3��B[}��*2n!`n�����ݳ)�H�C���`�57٥][dK��I��p�]�3��}A��_Ѝ����CA���'�o�}8��{���SM��֡�	�3��y��܇�WI�]����
u�'�V
���U��@��9�z>�g�|�#C��b���Cg�2V~�
�W����s>�h��-�Hya�����j,����1�˅#o��6{\j�Oi}k�d���7{��wk���Q���-���W���.~�e���G��<H(����c� Q�����6׳�7�5g�Mrᗐ���)�ΚZa��VVr@�?h���]�V^eG����-s�8�m׀p��ܻwf�K���&��H���Q8h�2=���R��g�˰�n�%�)ei�0�	�Mk�g����^>m{ѧJi}�l~f��9�} t�o�<�7d(�A?�t%>��T'z��kk4�g�P4V.5L��jt��{�Y}Re����%p�D���v��a���S7F71ez�E��?�5��ԩ���,�@�����s��^��+�o�\E�38�H\����*4��T����]\4Z���(�W�݀��e@����zf�s��ɦ��r��s^ �=n��<H��T��>�C�]��ċf�����L����f�Lx�=@��F�䠌�j�ϣ��q}��f�_$�]c�.�]H ���}�G� �\���n����R���Ʒ�	��]}�[��w{��Q9�ܴ��u�ɼ�d�jAq�%I��H�)���L�Ύ�e=��c-����v�ԺTB�s7F���[Gߺ�G"��jUX�??*��f������G�i�8Ӄ�߄j��^��T{�pԝVUN��JP����C�R-�����6�@�h@�Uv���C�@Xٹ�1��4)g�q��q�Ƈ��4D1��)��}S|;L��S�9�%��Fd2P��d�lX�N�2J����W�CUuD�L�B{��0릳��*kN)�J����T�Na=/���q��g9O��D���؞�[^$�^����?طW�m> �O�#ӥ*`�4�8@ٌx��x�Rlz�T���W��w������9�,����M �x���<���I�ra+y]��8�,�hf��<�Io��K�0{#��H"��J��)��8m~qe�l(�gt�C@i e=X$�ּ��~-��%6��'��IQ�l���&�h�&6����@�a�Zɨ��)�h{�Q���k!/5�U�h�*>'i/��i���PΞ6��<��X�o��f	�j��x��`v��Qϝp�I�l�re�aݸ��,l�-��]�����YI�Myǟ��l߷7�!����ߠ�3��R�Te/��D=Fw���G���׊��?�71�U���dܿޞ�Yɇ���߃j�g2P����M���y\1���՜�&K�ϝ/�1�I���A�Y��� �?k���7?������sv�XkFL[j�8���H͗�r�L�{߹�܎Ԫ/��ą����C^-#��g��eC�暄#�xD��ӭ��63��5�Sj�����#/�~�ٯ�����D�yAm�8�WCV0�[P�)��2��= �њ�(��U��(�U�jX�t����"♍_�9q���1��_ź��/�|��җ�A��!�[D��\�W=&`<�Jƹ������U"0�����s�9�^�t��O�j��A�-W�@�WA�C�F9;��h
�9��Aw�5nb��q����-kL|s�F1���N��u��_ډ8=���*���N\nL�pZm�^����b%���wz��������l�,�e��{>2 2�q"|h�O��t.�8��>2����}��g�.��;�-�cX}�3��<�`ڞ����^��V-�M=���������u�lsai@�݆T�p�]�?�L�,f;}��q�G�H@�cx��'��1�M�=�il3�i ���4�>ȬG���37w鐜.̓Q΂��})6w^�B)<|��Ш�k�co�mD�<��:�����ix���-$�u��w-�m�|�6J�*�i+�����`;�G%����BH�â�IӋ�Ui5���[*�%���?pf���w�K�m�o�aijB��9�N!z�V��D���U�<���]����#?���>;2�����'�>̹��j�}bͼÇQ�g�y�I�ӬrIx�򠥛\@s��5��P����~���!w��1<�Q��ۧ�s��E��<�!էz������L�v�/�J�h��bHz��W^�ėO~"��-�x����}�z��)@hҎG�WU�WӬ5���T�
�t��a��LE�9\�z�K @+�!Wi����X&�uB�.�,�����^$-SpW�0���/��rN��G2�ʤX��M=`����I_K���P�,����ї�"��q�x;k%[������	/�{��}Br{d���a(�W{_R�oI�%p��Q�ha}����W<cF-��o�֖O\+���X�� ��L���;QD�?���r�R��~����n4J$>')m��ָ�
��"���R��z���t��|��"vYH�Y�q@��`͕9���a����}����L�B��02�t坧���E���%�;J��(�|n	�j���L��Ŀ�Q]<}�Q�_�g�9��"�L��ۗ�E�v�,�F#�e��a���.����]��̩�03]8|�є%;̈́��,Dl����)&{[=hҖ���|����3��nSƈ��ѐviqm~���6*Dw�#ˑ�uN���݊�Ѧ�>Xً�5�c�`n2N�����~��h�iO@�mo�~w�odӯ���w>IQ�faJL���N�MRw��8+Pwڽ#��������G� )�H�Lpɮ�p�].ݝ,A����]����E�+;ϋ\:k�z����7=��,�X��#���J�^�%Y���R���Ƈ�#�����w�f�I����%
	�+6{û�/h���.��f]w�r����۵��A��O�6y�,�V��}૭Uu��n��˃o���5Ɖre��>���@tJ/z&tkÛ<Q���ׂ6�r�g6L�[�p�t[��Q�![Kns�kSsy����Px�W��p{�E}���_�7�B�͛3�㚑G��zE, E�(�Ŗ할]qX8�&�Ś�C��oc�}������ƁC�̟3;��W��	W�����0XB^�+��Ha-�h�m����9��c��{�uǆm�Q��<P��mV9����a�U�d\Ha��K�'y͎����k���p�#�dѮ'�h�xS�����n�h7}�¾�_�����rX\���8縔\�{����iףyö˂��Wo�������BSE�\����y�d��Z�wt��:��HX�T������U�\k��j?��$J�t��������a��++@攒���CZ1��wd����ut�o��I�<���@f5�#��#{?D��RÞ�#�C��%'�-�l^7��M匡�����s_���y�$s�Ný�ll�!�vrsC�I�������ҦέE�.9ϩ!b��
R�Ҡ��G#��A����Y�|��s����UlT$�R�~�
Gx�
?���]^�}0�;�X�����&Clo��^s�Vd�91'[׽���B�7o����W�{[y(�nT_��Ơ[���p�a|3^AxlXׅٴ�}>�y1����z]N��j�@�4�3��ǂ�<�J�� ���:�5�Ҧ����Ш�[�&"J�z����!�	M?�=xKJo�C>��Q2�u̾�b�6�_�X���3��J^xoȎ�t�pużC�H�&m8�
mM��[;i}m���
k8R��'���zo"��Xv�h���VN����:9�K��%�|���ڛ��(�)��r6�`��W�-�8E+�_!6��gX0=�5EV�1�Ey�v��G:~��Kǵ*�TԞ��哸bDz��tBn��~�vwկ��1�Z�<�ʲB~�n��`|��Y$���%���=����}sF�NgA�?h��V�
�V߇�,L��f�|���t��̕����4!�s!��ȅ�<�d�Eڴ���PFO�׌�'Ǻ�i�YT�s#ji}lȯCV�+�n[|��'���
#+^,U�!8���
7T��3���./�?��\#�t��j�������;��,)���r�M��m̱��q�q��)�6I�#I[6�I:�=נq��۽+*$Յ��N�_�:G"�Zz�/��b��h����D�X�1Wۂ�1�<>�ї��7Y�=O�}���Ǌ��Ő��+�ߓ9�
O a��m�0Ye��Mwu�j\���t�%��,���?_�c�T�۵���m�1��������$��K�%�����g>r��ba�(q��,�U����u��w�?�le��I^�z%��y����q7��h�2��t�}9~S�}�!CT�ɳ-���M�j�^׎6|lg�wpj�4�(�R6�2)�֦q>>w�X}��OҰ��Z�S)��zT$l;�^��j��^*U��Jf3�,P��Ũ����euv�Ѹ�&�
�4�?�Q��Q�ub���G�g��q
�HN�������}���QoNg�����\�h��:.����#�$dbatn��3�j*D�(�O��uW0L�X�if<����8�g�n!��e, Y��o�b�j]����O�􈣮}=B��(8tj��j�b����$�Q�0�Y����\Ͽ<n�ɱW����P�W��O|�P���ycd7�݅sl,gk<E���4<���/IE��\bL��(�
h	$��+�v'�'�Cs�="������R2-5�G�n�M��Թda�͡�6R���ֺj	�6��z���C���%3i�n���&s���gN-�.���|MG�y������,�q[3�5t�q�G���4�LY�`H,�,�GV�u�Ů)�;?8b�^zMG��'�#�l���e1T�v�$�#K���������4�4����ʕ���Ԣ'�b�<=gr���>��l]�ܪW�ͥg�n��,.D��1$ ͪ��_��� 7��;��u��.U}mb!���#���'?�@cJ�u]�������A�<G��5H��N��Pv8�ܶ���c��'��֦D�?{nu�P ���^@��&�>�F���4�B\̊��.��.P��c��� �{����H]޲�E^�r_�(_ɝ7 ��5e�H������<�A���B`"�|���'J��K��yDӶ����Ӿ3�r{�r:��zP���w
Bq�v@L�����\����+b؎��?J���[�1붐�cv���[���[����Pq�Q#����fO`���I��ԡ�y)��Z�+n�C�������v�?�L�ӣ��cs��=���e9�$�o��3u���e�[�k�mb;�D�?��2�o��gcc91nv�Co$��/�L;��l
�z2uW~��߼Ƚ�nj���0�#���kM�@p�����덋�!D 0���@U$5iM���p�9����F&�(��|}���m����k�6-�|g��0nٓ��opl�ҏ y~H���)���X\����%z(݋��)D�z�����և����nw�b���⻿�!k	i�.��:��m��o x�I��-'���.�݅��M���mE19��IkL���=I������}���5?��zl݇������;[���?u CX�����FrN+}�K]�i��27�$X���@ ��u��:/w��C�)�)�M@�R7|o9 f?ݏ��;���p�`S��=�.x,ys�RQ´�c��sF�i�u�d��hm<&Y������Ë���y����޲C�����c�f+P6�*�nP������8���\�[�Ƕ����P��b�"n�T�̐&�h=��L�gk�%�녛�%������}�M(��}�H��A�IҴP�9ⴆ2t:�I\�hgXE�a�1�\��,��.�����@��qW+_)o	O������<"��C�G���=�|�W��� 1�I�A���W���<�Կ��G���3�k�q+�C�"$�\��}���q6��ƫ�2eZ������$U��������N�h��V��b���E��Q������;��œFW�8��7�"VkĂB����"u*��2C$`�f㉜������б�V�����>�gD��M��)�+��_�3}����,�PS�Q�t%W�
�J�����S�4�5�%4!2[4�/�H�7�����ך�bb��q�B,ح����W�41��: �@a�w�RW��M��Y���U`�K������O�sW5@�<g�ܴ߹��[��pm a'�O�ʗ�������[�����{}b��߄B��%�x�# ��[��ܢ�Q��|����A�M��C�KI�I���Eoi��Wc���@�	�	���A�Dw��F���(�)'kw��zD-�2B��r1�f�Ŗ[˔���ku�I�P\{��/�^㩮yׇ����m=�X�7�x|}��^v:��Y�=`�SeHP��~z~���2ғ�d�'6��b43���ڜVZzm�ߎA��lH���S���;�q�$A��LF���J�=���t���O�����! ��Ѱ���h��L ��[�s)�����viM p����ޖe�PKc{��T�p�%y��@hl��(�ʻ�%Ξ�uܩ�Bb��*�daR{ ����Y����ԽS�)'����a7=���qCu{�}�=L���f�g�	�����11��	�e�j�fGc�KöhA�*\~�k�#C��b�K_#�s|Yf��I�E���c.g��3���GօS���{HEi�16�UP�L��XV?Y��X���4����d67���hC�H��%!4����m�!D^�D�h��tA@/>� MW$�7'V���\w�?�N���}�70���բ��+�<��0yl^����W�I�*ګqu�b�^,%4�ᦕ��FKG��V��֭�d�we�>J*���5��Rɥ� �K����V�T�.�9Mf��hv4@m���w�ED���O*�l^7V����{(|�Bj�ܺzms��sT
�)��E�l�L�Q�A�b��F�[�l�,���EPx�>1��,�u	5$9��!�.+Qϲ6�Q���qΘ�L���-���*AU2y*�B흳<���] �C��~��1PANf�����O�ev�ϭe�����u�>�O�H�׿o����Z�� ��.$���s���a�P8����"A~� g��P��<�_�s"9u�Fupp[l�	io�z�d��'^�I�t[?�iw֯�*���AA�4��(G<5%�Uj�*|�P�������M_��wB�����^�?QbPy+I9g0=�\�����,b��E^'JP����ڽ��rĮ�n��]8��j�t�g�U���˂���{_���a T�%��Z��3��������ҕ��� ̻����٫B/���\���0��P�q���3��� ���Խ/6�UÎ�%�2` g盘�����L�D�z��Ǎ�D|k�m�Osc"z~D��,���M��5AU6^X0������@�r��!Ǉ=*d>�$��_}1��z!���b�[�e)2ۃ�h�F$D���th��ك~����������RE��
�,����ER�"�=�=׶��Z�((7�����ܰ^>̓�l��nAn�h�n'NJa�Z�M 9��(5�F}�Ġ�����I�Vbe5�J�v7'{�a|Y}+�S_�)�D��j2�p�F�åK�������������4 �4d�9������h�/!�!m�lp,R��{jR&�H�!3!w�f�:X�9�;R��~���>��:O#�|9�
�����z|�\,��8Q�L���m���3���tIQO�D���p^a��}<R�z�É�C|��
���w��G�t
��|�[���tN�6> �����j��&7��6��!��+����s?E���p��W:97�]��E�z
K���yc�X�C�l�e<j8~����b\�E���<eK�Q,�ȢO	����}��kٛ~+�ز{�O�삲M���� |@=]a[���C�vleޗ%�~�*"ZK�*����R7  8�kR�|�Y��ʯ���Dc��ʰ��|F6�$[>]����l�:D�,�u� �4���ll�	�I!z�M�@�d��`(aY�=1��A�PT8�*(k�^�V�W �
H�T���8뭝�M_��Mz��|C�[�ʶ�֒Ĩ��g!;�7�;�WY>Uc**��+o�
�w�[�n�lΝ�|�]�Ѽ���34A0���5�����}��3�ZQ�OY5��ˮ�����9��f�
�V
V?Y|ZB��LE�pCR�4y\�E�3�/�N~&�%2.���UW͢Nf��"(~ ;�0��-x�q��
Қ1R�z�ix�pܡ������c�%�C��!Pf�Ӣ��v�̭[� ��������zD�;潄C�MP��uleB�7�E��/u�u�I vh�<v�hL�������
������\���և��b1bE�ۭ�F��<E���o�14y������Y4j]���QTN+N�Ya�߰�6A@�odRְ�I�� Pa:��)�x��6����&D�} ��	E����}�:}��gn��M�tQ�J]�T���������qq�i�� �e���Y�4]�U��,T��R�R�F"�Ʉ�ܐ�_�8��y��GyF�	� ���* X�ᴣ.�c[{o�g���E��]��܌տ7/�9��X�V�l�,ѭZ�ף���EKyP�ۺ��2�����-�[T�f�M�O�:�V}�{���i��������7�-���r<��|�&W^@��d��BC��U���!�֚��ؘ��I�n�S���ɺC_��8��QlT�,TT�ڃ��zG���\ֲ)J��1����J�v���'i!�9�l�c>or�X൛�6����MU^��A���dW�QE���3e�3S�n ��	N6�� n�(ġ�G��{��_J��8+�<D
AY��/�
�na\�Z�e{���?N'�#��<~��//p��Vp/�y��:5������ὴ�8��EM%z���j��\� w��t�6��J�PD�Ҽ�B鯱gYφ ��M{���q��Z.���b�V��(��ڷ��Ӭ�6��hh���=U"�f*,���6����O�I~����?��<���_�	�h�[d�wb;�D��J	������u5��P��M��w�~m~A^C�NQe��,s��^T�?�Ǣ����o�x�1c
�����Zw�a�hk�q����Q�=Ӿ�U�v�LB���������i��<N�2�ô�-m��_m=�!�l���x2�Iqbv��20}�b6s�yƺ�y�w�u{�;���<q��eP�a�~I۪?w^=W�������Y�Q�H�In@r��-��|&���~2�l��4'ws�}�t�p;�'V�0)H`�@Fޘ�6�{u��-X,����6��$��
����>��鷋0h�G��T��_��°݆�E�n\a� ����Mt����Gڥ�;@M
{�f�f!�M�q��}w�f<��@0�u��7�����Ow�A�p�l���tDC; �i���Wڃ�%{29 ��{�� p��)9%��N����c,�
��B
L_]�0�6Ӆ����y�,"��OR�)]dn�ǬY�����5�i!?Dʾ��+: ��Y�� ���!�.��珢��6�����"ڗ;שs4��	��}YO_����4��!�"p/]��AW̺!Q8�����DWD�$3�}� ���%���t���E'��#}`��\���;��-��l.ˮU%���R���	B6���c��;�ڊ{H��IXЬ(�Ӽ���.3VM�v�&��I*��4��OO���+�9u��F�2�J/��!/�����n� I(�f@��i�'�j�Hw���y�A���C7V��*���YU�>����=��=>��AM�� p���e�ݮ�͒��ڔ>��;�BFBH,Җ�>E������%�����}+���M%�*X{^��OJ��`(�tu=��e���tW6���}$J�(�܁� dm5����	Z��	�����e[Մ?O�r���
��(�X��\��zH��?D=����O��zg��� <��Fj	�O�|�"G½HK�>�`�9�Ib���^9�]�^�ih�/d�F�q�ۏ�n�JL��uK�1���ʦ��b���Ni������EƫOZ<�����F"ό��p�]b���%����K���K���]�{�ƣ�U\�u=��1���K*��N]J)3	e]���ruƌs���s߸F��[���R2e[��äV�۔���;D۪�6@�)g�X��8�w�R2R�g��4t&N^UyJ�{ZBQW�*���K��5�}s�+�AS+��a	R5J��%e���D�݂ΈR����F���i��&l�d��z+Ñ�&�M89�9�e4�{(#�.	A�w���R�
TM-TU��T�6��_��k�K}9�/:f1�l�J�
�K�a�_�a3P��`g�A����W�s)��4`E�K�ܒ��ӭ����ɝ��97�
?I"�ԙ�(��R�v�����a)<�\��m㭗-ꋘR�έf���Z�wN-jo��PiD����f?�tGd+,�]Fm�"�C�W�ȹq��?�#��r��yu
���M��%���-y���gN����2��;7�u+;ݏ���C�)����W��,��.G���Y��a)��Mg-�ǌ9s�e�ˮ�x��p���3�����4+ݮ�F�>�N���wN�VFrY�Ԗ �MO�G>�lWm���� �� �f��?Y\�$��#�;��^��Jբ��	�O&�V
�7�R�O�	����E|̯i�z#hN莨ߍ�l]��ޜ���'��5�-����C@¶#%� �:�AVF��b�&+���w�y����҉�52�0:R���/�dX$�P4X�P�`x�6�z���ɮ!�U��L��_m=��I��!�Lym?\�ǂt��#]3�J���	��*y�3K�~���r@.>�'�>��k���k[��O�gȗp�O�)r�d������K/�j*�Y��|�����N����|^ʑ�#�.(�.G��Sc�L��r�`��3ZE�{�3T��_~'C�#�'���A��g559���-����Cֶ�7;��h� �v�� c��b���a�:ؒn	{�m��?�=<<��v=�V��d"ԩ�$������p�0��ɣdr1r���?d����		#D�G����wr��a�f�3ϝ�y�I6J���o�����U�'�I&�?4.>�&�4����7r��{nÊ�}��,�a�Z�� R�Kڨ0�����n��{u�#�j�D:8���Q-Y�z/���sz5%��i�+Y�Dh��oKJ����Sz�D�1{��/x��r��b�%�C�V��-�p?�,�F��!�߶II�e�=�߹���
xg��/-��Иl���N�����ɡd���s��kUx��PS2��7��h��?<�t�)}f�!��8�6g�5*���i'�n\}|Nvr2!��?s��h�C��������xv�z�WP�`}⪩���[>��b[�Q��+>WU���2��t��{&/T^�KsR�$P�n���X�>2d�_j��Xʴ�����̡ȳw�ېV��T���	��۞ԉF��ɅO_��X�?�$��mTR��Θ|����Uv"i|�pb:/����t�C�ϕΜ�T���	Ee��	���r��-� �/��E ���M�D�GϱwOՅ�N�l^�#`EZy�I��:)y�R�o'uy�;�N_��b$��r6dS����ۢ<6�O�X��2�7R���ρ��������J�ss����!qH��6>U�ɷ��%F6�-vR��X�*�t�*�0��Q0%�D=������.P�����^�w�*��2�
*�e9�1���2��%2�)sW*}�����Ry�5�T���7����m�%Ӷ9�v�����̉7Be����N3�S��F<M���F�%Y	1�Ł�LYO���;ysȢuק���Y�R�CyN[���oFy(ֻ�Ԕ�<���
,��[���滐3XF3�5nfe��F]qZ>/ {V�?��T��,yy'p�Y�����L��d_�D����K�?��l�3T�xDj�锕�L-��E�?��<�V>ן��m�ԭ�k�qZ�D����
's������;�[m2�;s�a[b/||��
D�4�^�����yˤ���_�yW�"k���PB{����ͺ�hXϴ���*�FU"|��oR~����~68ՂZ����i)t�7��f���~�T��<�����}�	�X�i��ÏvE����7K���idmo���⬪fKd]ѭ����Tmm���|�E��?�����ҏ���'�Y"��Z�w�\�1�����Y�]�d�e�xB�;�^խ9
��D����7!�O�d9���4�j��u��9���oŖgk�fXh�KrV(R�߾�F%"��JԸ���0����N�TF�����,�;.%�=`�����3y��j�X9ʮT.E2�%%�����q)�@�K���|].��^�
z=̋�KA���J�/�S���C
�@��m^�hm �h~+�_�s�!�ؖ��P�MQW�oY�Y�/J|��\�/4�hx&,�E;�����*҃[)��c�\��0�����z��\S�������?KE�ī�	ʮ��ؙ���K�.o:�}2� 
��#�}�2OutN�BW�%�������;[�Z�U�o��k���j�"�� o������<�X�r�����wF�Z4V���[��á�q�ؕ�-4�tJ�;+�؄(���$B�~��Nm�Gct������መ��h�r~pLM�`M%6.K:��X���F#Yn�lXkx�D�����nn�r`�+C��9{�.@C7��*���LKQ-�yԙIc��(�y�w�y�~���1��Ē#��b`�c�tc���>���Ѣ�A5��g���JH������ٟ�>��jM��(N�$���lu����	�K��u:�-{X-OjE��pbၩ�ce_N[������9�"vk�,y�i"AQ6r�����2-W�j��F�J�l��W	��?DN�Z�?5Y
R��/���ʪ����u�"���
RuJ¼�"ʔ�
��H��:�-wZ����1�<�Q���M!�b�"w铸~�Z�.��ߞ��/���ѷ����*���gk?��61���.>�~��K>�^�|���WB"'��RWi5��i	&i��)yDCHEWH�K9��7��ȫ�<��V�h�q��]M�G(�!�����7Ϩ�3��Fz��
�(	.|�~���c��Y�m��{ܷ`F�?��z�B� �z	Mb31x��s5��*Oc�|�sK��@��WR~Ց���|ߙ��I;*�ܮ�$��/�>�s'��*����-�^���G��m�J�-�}�����t�*�n�����v��i����ɥ���V�_o�J���pR�\v0CMQ�x��%&9&n��:���c�X}4�*��!������_Ӿ�Y䜡��jR�62O7õ� `�M���Ε�e+��vj���2�����^�{�b�uR��e�n-$�&��-�
�?t$XVf�C�k�K�+�G;�fpm<�e��Q��{9͈�"k􂬸j���ްu�1�F\]p_N��rF��q*�.�r�Y��.�s��`e\kՋH�{7P[.�V��ԁE������C�k[tYa=b�s���T��ﲵ�:�|���}+���/�e�'숷V-K�5o�`ظ�W��XK��F͙<9��H�{�?Ru�@2�x,��{�T����Y�b�!�J�ǃ���uֻ;���OKWv�ss�sd��-_�����$!��m��S�;��������Dpmg�\ĵu�]�{�ח����Ù�*�V�s߿{ԕ�:J[a�Q����!_��V�+�οE�8����E@q��n�g����\U�����&�Oо.;}��Ʊ�m}���o���gv�O;�y��9fW���W�X/�bu!={�{���H#-�3�e׹��ø�+B���U��~K�\E��u�s:�Y�'e��s�I�a=2d�"����0K�i� ��q�.˪ i��-R�O{�'o�y��^x˜٭y�O�_g]I_��z�b�+:Z�;hy�'m"�g��FD��+ьؽ��I��O��Mw/�J��
|-����5l���yI�����tӖ-����Z��T���aI�f`��g_tt�N2�̾�ZSƎ�?�	Yt��z/�Qe>��b��٦w8���C͙�[�-��n�Oz�	���X�C$SD��A;��_��.�̬lX���L��)<$���f�,���t�/�;j_�}7f��߲}���9����W�`��|ΡEu�S/� �`��c�U��A�bQ>��6�-���-B�z�o�Pʇ����+g�w8�o�7��<G����?�a�E�ĵ����Yҗ�%�+'QM;��ʣ]׸���ԣ�2���(/FX]�R*�zf�,���G�Z��sn���'B����V�>�搴O�/+3����%I'�w/�ED�L}�.�y�Q��=��||�8���jFcqE�܃MS�>IJk�����̫����
��FL�"��vS�V̺�r�-
���3�KD��Y�.m>c�`ZCM���X�� ωΫ�yb!bC}��!�յ��8�켏�H(��4���Y�=���pV_�zee�7�l*x
WB���@(���?����s���o���B��5/e��:rժ�˖�n`��e����&���^C˼��5��rϕĹؤ�Ï��?�j���[v���w�_�6���F&�্�E��rT����h�zZ�0a��=���n�i�ڪ���Kx���O��l��皅�%��3�5����������`��s��A[��X�	c�e1�9.��
�/��E��J�����`�v%!�}�L�Q�]�B��r�6������Uw������Q��hΛ<LB�{��GG+
��(Úә<Cm��j��=�7Fe�������j��Ml����s���H�,�,ɚt^����aQ�]ۃ���-*H+
H+ݠt�]*�94 �5Hw%C*��94�ߞ�}��x�����^׊s��\�x|�b-԰�7P�SK��ju3V�_�D��v�ǭoB�{��ů��c����Y�.Z�7�!���F�j����d��r��~����Hq�򑸸���&�f��u]����m#jN�Is5��S��R�7��L>�O�����w�Y_�2nF�q��/|#��]�K�!�+H����ڎO�-�����H"���ϗ^������Lx_�|ҥ�2��������`�l��
����Ս$>`������|��q�Bcu԰���]/�{�،�BG��$�Ƅ*�8���eH!�ז��q1�+��8F��z������'�w�F*��"I�9D���M'i��)e̤��Hܣ*J �֥�}�o����������l�����N\�1�ARnPM�}p��Ҁ���I��|�B`,#�8��<!j	`�g��
e1df ���J�N\����Ё�o����ZP��=,�Z�B,6� ��,��G��>2��&�F�t�Z�֚5�ҥ��M�ZUl4v�������j��k�$�8�H!�a�iޭGg�R�x������+�}��fedj�mF��u��|�rq�7�J�9܄c8)���u0�.i�"�<}fM#��C|� -��e#r�)��[������Su�g��n�o��N�d��R�R�jX�Xgg�0҅w�g�^{�����wi�5�{Z�־��EѪ}��0g0�l([��|g�EG���u���l\)�ʑ�:��r��'�qQ�	nM����{���IsW���B{+��ܞ�J�K�Ano����2�Fʐ9���f�! .�3w������,)�1v56U^گ	^'���Wx��c�w���=��U�dy�k�]R�y!C(>�C?71���c4vP�t��{�����c��m�������	a��&�O+h��T^.2_{�;��j���&|	���C���m������֬�U������s�=>i}�^��J�������)(X�P��r)�@}]����X�y':7�lP�ܬ4���"3h/ꖂw�Jx_/R�x��2R4�%���
BC��p�D_CP�aG[�!t'ld��,vס�4��z�߄E�'��Tc��1�CW#B��@j���N���zM��M��ff6={3�O���V�ޮ1�;@��]�QU�q_�#i�M,(����?��o>K���B��ۨ�&�"q��e�x��:�H6��z2&��&����(@㦚���i�z��A�Q��b?�8����_Rɡ�"��Ź��wXك���#T�2IEU"��s?���V����@B�9X��Iˬz�%T�� �c��i�Q��Re�x�˃�v];�@t�i*��\�tU6ͮ���5�����Q����������� qe�{�'��vh�?�W*[i�z�v�~$��j�� �_#�#=�33:ȵ�W�'�i��:�j����@]sL��Mm���4�:�ڢ�(J�$n±|>/�,�"��J�!�}(lt�w�1ԛ�F���7��=�n�xY��K�5�c(��YŒ��ٛR�� ��G��P�r!����O�v}���2a���y0����� *����Y�ڐ�i��$����Ħ�p���U�Y <v�x`�D�Y@�nJ�Չ"��8l��G�	�$�]]SVR��DmP#�q� #�˖_��r�@�+uM���2�Q�44��LH���G�6��Q0Ϩ�L�B.ĝ��ߍ�b��X���s!��`���Kp�e)�Cz�l�̸�˫^��dVz�r���!$�#$�����k5���E�`���>��1���|��G���i�П��I��j�%k�ʁh�x *�:�����Bü�U��������l{�h��xf�hޒPtfY�3vEh�="Wo���a�:׆����Zl9����8�>�J�Z��m�[�r�����TY@���Db6ʳ*��(�R��	\�u�4�K�ƳHV2�t� �E8�Z�uT��B˟�~ҟ��7HC��7���~A��.�2�$��F��Ifw`��k���h��+��1���ˮ�cD�ܝ��)�Dt0y~�v/�k=�,.y���}�B�����\�k�I:s���X4S�����z�/��	�-�?�.�?����%�6��
T2�%�'�4���J����o����`3=�y�yC'K�o'�����߮��P��/#�Ɩ�,R�M6W��)���'\��rԠ?=��%r�ɱ~�_?��v���qބ;6�&��w׀�G�t;��~�Ѭ7 u.���EHv��i�S˫����=^!�[�v$6����^�_:N �1�����]O���Ҙ��I�)g���/�HxI���ѩlg&��ǐ������~r�/ɂ���Ҷ��\Dd��c���<~L��
�0G8+N"K��W��$"~f����Ђ�/7"��D��l]�I�a�L��s�f��Ǝ�����xJ��!I�N�=�}aCA��q�ǥi[�R&�U�0!�"���~� p�ب<���
����ir�	�p!G�N1����6��{��!����R�&����ˉ��۰��G��F���15�##��|�з��m�� P\��R-�`ܞ���?�Y�1���eV��T��
׽�ODp7i$��q��AΦL�tM��Cz���H܍�n�"��c�鹦{vcD�̥�0a]+� �M 7�3sXX>����s
�����qoX����,��S�]B@���p8-�9���:���xo�s�F�{bK�g6@�p'��Ў�.>��?��$8�ё��F���B$N�P�·���o�v�f���]����:�U��ݞ���C�K��ε�!V������Q��<�w�G��q���{J� ��i�%�M��Z�j>�4X:ow�b��/X�CP�?ӟ���o����M1�������������{����;�#W�*w�3��x>��3��� x�&����a����/��Z��9׌�%�=�1"��H��|�u�S`�ߠ�!>�X�wQzSw9Dۧ��{��5$q6y:���\wA����we� �.��٥��/�~+�FP����-�j�Nfr����:��Lp�q�1*�ώ	�o��Q��&1m�i��~��eW?�����0#��jA��%�oU�N�� ��}��k�9k��g�ט?����Y@��k(.+v���I�i�Ƕ���DA2@�� ���4��E.
H����G|s@�{��9�eG�\����	�3kT�L}��XW4�na9����;���8��:a����զOVN
0x0S���@�xU�oTFX�6�Ȅs�Uq����'=)�Ɔ����=c8��pH�u�� W.���^�\��Ƨ�ILW����\�H���es��Wpx_�@4�R���
dJb�\�������IVp�p?�ְ&@��Y6Kj(���6g��	�b۟�>���X��L� �nf)���v���6��[����lY�x�k�3G.ɦ\�=�࣭�Ll?�� K�͢
��I�m}���?r�NT
�S0s�̳}�����8*��HRQ�نl�]k�mJ�Q� ���w<��7��������ɋ*�<y���[&k�gE�g�ɇ[{�	u;
�D5�]��:'�� �t�Q5�ʇ�O��P�+��Wr��;�]�T*cD�li��X�)�۟'�����a�.Qnt��Â{ѕc�7q��KO����`�;�]��Ӟ�����28ٟB������w��15�+�)b���@qLZ��ION����)���Y̈��l�~�m�
6��+��s�f(<Ȑ_`F�:PbG�q�;ޭ��Ii�(���x0 F
��� S���]A	��	R/ `��{������]'0���02ՆIzV��vS�\����	{.j�*����dP�P���JK%\h�������r��M�3�oH����J;�$�C5 �o?:��2��<�e֙������sk^gk���w挞?�n����������e�bb��1
��^ m�?�"���ۙE��D- ��l�{Y�2phx���eL!c<P&�>�����G�� #����F0��}&[!���hl5 �v�F�,:z��]��}�kNem���}�MM�9���L�؛�cJE����������v���������gM7��Y�%����W�k�,E�H�e5j�x���
6?��ߥ^Ti�������V�F�հz�|���I=�Z�4b�&� k��&<r]ߥ�����й��	@F��+Ϧ}�Հ$�C#�F���l΍��Cr�pS[78j���5a��οh����� T�.䯶SS�ƨ�/f'1jb+����0���Sz�հ�?�Z@����{��J�Ȓ+�H\��O��엢X�V���KPK�#���rޑ� �qW�����6���F�����\�Y]����,G��C-���#"5@����Z`�*D y�r|v��^�S�o�	�ΫO��N��B% ;<�@�p���j,��Y!���{�����1�1�/����V�*��m�Ll^l����_�n��m&��5'X��>c�ܤ�G�h�W����"�XW�Z#Z� ��?Ru#~?��9���!"�y�ra2���i;|�;ke���S�	$:c���]��̡��|���whAB��{��ƆLH^��K:0k���P�����m����3}8��%y3� �[|��_�3|!��]�hi4V��Lɟ���a�v��$n�]Ǧ�+d�\�Y��W�y\�����|Q-~/F�%��n�������ˀP_�Ϲ-��M���-]^��Y�'v���~>f�r�j�BpG!5��.�-JX�t�����S�>�$U��s]z��{�V��gd�
,EJu���m�	I�w��xD0�MB�������M������&\g�\�]��r�I�O��~=���/����A��.E���L+�Wa��E��(n��m�4���|��gυ�e�)�M������"&����z4 �d���$�?��sn���<��uX�T�q)'�o�<!�Ax|��^T�h��l9�j�������y��M�~����mn=�����ϲRf0s`���NW���ށ���|�`�R ��xz�\�8���	z�c��kI@;r��<��[���ܕ_-�
�M����A���[��**`�=��YA�W�@2�aي��,p���Xp�
§��k�x� ��=�YE���o�Ub���,�}�*W�*�)>#r�rP|.���\����`�V���e���o����ԑ��f���V.:��B��mǡ�q[E� ��E���\�������{\�q�~Rȳxr�f-���|̍v4͑?��	)@.[*�e'�%�8*��Yrs�K��)�͐��3x9���*�HF����:�Jc�"ru��r6�V���{�'s~��+��43�&0���l�㔠{і&����wҢ���˶��l�;p�l�~n(���JZ��%.��-�*b��d�Z�ڣ�!��J@UJV�]7v���+{��xEY�4�*�K�}9u��B�Z�^y�̋ �'��a�$����a��}EN��粦{6C8k�����	�v�m镔����O�,D_T躘ϊ�\�)Ff�k�6�v���H��g��� :�M����D��]s�MN�!>:�*5���`Z�xW��;�У��u���I��Utѣazn/���u(>q�kl��:;M"��q�=	X���{i��qw'կ�����-:�q�痁�E'k�M��QGEq�t�<_�`J3��5	j_�>-�]t%��F`Z�~̱4Kh� ��V�Ǿ��e�ƾ3�ݱ�¸�y=������t��5���:�|��s�5Ҏ��ڢ�5���.)Ώ�nӭS����j��A::܇�|��?~������4�S�K�Te��Ib�������o1[�|:ox���/��Q�]��ʾT,����N��}������~7�U��ؓo���N��
1���~~�uL\J@e�������}/dr�'��b����������]��ޮp�_5����б�{���a|\���n�g��h��G��+��f�;S�3�grL�#��<�&P]?�?���y�����)V�ⷺ�q�|x���������2�С|�Rw�ϤS��Ej�N�?�S}�.7ڲBp��̦�Hr��?�^�	���Rjm�HBUeͶ��O��p7i.��A?���<���x���a߅���9ѓ��}�RS����W�G�:Y����J��&���0��%(�{i���Բ;��בrQ��d~���G�ү�Zat�!�4����dH�+Ԕb�>s�U���o-#Y]��{-�7�8	J]���I��F�[�1��6���l���Z���45�*X�^��9���F�"G��/��o�ѹ��f�3yBY�|���mMJ'x)�H�`f�ڿ��Tdsl0y��͉�߸��w4�F�蚉��͆?��uHb@^��e�Q ��W�5b�l��Pj��0�"���p�˗҃Y|rcϕ�4~Ue�: qDk��_MLT��UlQg�˼%u��~����lh�gs���K���^��/	�@�s�˘C����D���볥k}��	=��GH��ҪOU�$�T?��g3U�F��-[�l�ت5��vc��,�6b?�5��l�F��c�(֥=��ЦZس��;2�ˣK�{�<�S��*���쫍���x�
���-o���ENW�2���J���jI�^��Kϡɫ�����?�y7q8�%���B'1�,��M��%:��CU>C�=U1K^��j�<k(r�(p+����d5?ey�\d��Q��
kO��s3����q�|6��ٺqREk���zĕ��cj)�A�y6��[��n�1��#�o�=e�,���y�kf��`������!0�%l�|�};�p3y'bG��roD>�a )ʦh
�݅]���σQ�!���i:��p3U&z����}��4�+u��XuT4RV#|=����I ��[����l|�I,`z�T$�����*�q���ע{���bL�I��b��p�Hͭ���c+�^�b��X"X}���G�)<�����iI�L�.�3h17��c�ehR��������;6S�_���Y�M7�*{�#��������P����=M�87N͔[1�l���͍��fe�"G����fމ"��tQ�G���f܇ѩbsI�j��LȬ��ٝ��-k$�����d��e1�Vh=R����#M�o\�\�d���7��l{��&t��4���ury�x�r�ޮQ�T���Ǫu��4����Q��p�����X�1[�!�T�E0��_��F$hvk�k-𲀧�*��]MsOi������m��<�VZ�Y*Z�3ü&*�����b�jɦ�0dUQu5�#�)�{Y��/I���T�o2;9ޖio�����)w�W�]4{'����g�To;���|j�#Xe�Z�ؖ���Z#�M����r��֖kw	�U+n'��vw��=�J6O�Ƀ�wqXn��V�M'4e�\�9LO�
��ּZ<�1�[��N��st�⇒gJ��.&P@�j�=>J>�1W�~c�}j1��we
[�m\|f��B�-�߶�r��$��K�����^���x}��E�����2eP��F��z�r�0���^��d��N��{ޡ��5iS���W�jk�J0��6���T�~�r!�67k�Ko�C���~��@�ƴ��>��`Eb7`
9�aH�ܯ��:a�7:RC\��/��u����%멡�Pf��F������j��>U�h7��n�ݿ� h84��
.4F���c� ��cuI����]Z��V�n��靼wő�P����^�����;���T6M�n�E�x1��Y�S����{�!97�}�&d�Ƒ'S�*�#Q��X�:���2ļ)ɞ��O^� Uyf�`:N�Т]c��C�ՙiژ�7�p�UD*��M_����l:杤���#�"�_�#�o��F��7.��zU��
4ׯ�{�/Ja��TfX%��f��wG
��
��խ'N�g��7Om�o3�x�j�F���0�9��H+����9�}Up�{�� `�s��X�BT���5������3�Dq�Q�����v���8���c�p��������}����=������m��󪼸'JUc�qo�Y(���w)�3yœ̜f?����6��`��A�H�!I�4��j1��ؠ=P��g�+[O�$�3>eX6�ux�f��Y0�P� uZ���Z�,@u��['��)ļl���l��k׊o@�1�,�u���Ň(���WN���s<JnZIe(-�/���C�K,����S��Ν�����h��N?\v��s*{���m�uf]7+�{���!^R8]@���O�Bc(���������!�1�S(��^L��/s�?NK<�<�@��޷��q�'��Ƨ&LO��.�B�j�`������v�
^Jֳ�K����8��Ӣ^�|��F�r�	��80�+9�cN��q���.�-}Z����R0Ꝭvo��o��G�()3ʵ:uv	�����#Y��}�U�V��}�Tɲ4c���x2�n�'R}��5?�U<��X� 5��W���*�_-
w�ލ �Ǿ�{w����Z�y)VI�����*|� Yk��G��y����;m��"շ��t��e�^�^w2�Ui=�>ڞG����u+��U���6��2~���*�W�"�ni��ѱ�����	8�	N��������	M��G��W��±H�^��v�hsh��[^�M�ӗ_�8Jє+u��e����3 B���o;,��� ���V�O�����
�
.�ގ���-wL�=�qx�?���J����+��^V��H��/N�x){m���U�S�]�-u�u��=:��@��t���0����A���M#9�C(Z�ka����=��7��ڝ���S��˸��6i�}ƇZ0��%3olH|��58�Wz��䄥#sX��ͺkq0?ւ<.D5k����+�ā�7\�Bx���(fn����WN[W[y����n���%�!9$Yϻӿ�q�7pn3_�x�]��jlȵl��[�$��'��c74(1Gl���|j�U�mt'fzn�mf�?š5�q�������U���gU�ܭ����R�g���k�VQ�{�5[85�mX��}H�9G��TB9\)8�B�r �߹�S��;��o@�i�Ywg^�ƾ !-;!ޣ�Q�d�����
�fm��Y��_�sm	��K^�7��6�*#��U�6M�C��xu����Z�9'?v	"u��R��V�0(��25~�itUm;k?�|���2W"f���oP7���a����z��#�#8!�����L��ϊ�[�"�	7<j'M���"}Y�)0.�_'�O����z�5ea(.���l��R��V����9�J��g\Ay�|vl�u����.�ݯ�U�k"�C�{�,H��ߚrP�C�k��kl��2���ޛ�
>x\~-e\o�'�p�݄�>���*�y���]әh8�w4^U�&�p��S�H��m[I2�t>�lw6�t���uD��[����������:n3*���#X�ب�?W����R�������Y��f�˛�>��cu��cqt͛�����ԳC��s��x1-z�}*�P�K
U���4���i6�Ǻʄ�=���]C�%GAȱ�&)ȕ�<��� �i�T����@H��>5"]�	��[`)-�I�1>�	.$�̱Ǉ��C�ŭ�Mg2(O-'�O߬��6�d�N7Kj��;�YE���C,��_�E}���Hb��=`rF%����+�����nsL�:��N1����E����ً�q��I�[OԽ]tXm�O�RS7[�3���p�L�?+��;�&|�X!��fJf �U��ix��f�M��2���/�i#H�4�qA���"��&���d�{;Һ2d�b,�=WID��Ĉn��K�����)bxJ�+�9�e,�P!Ӵ��o��/����w��l�x�y��ӬXagو&_I��C47L��v|#.�,��ay5�;�hpK~.:�Ԗ�N,��u�-�QV�\+3Lq����a�:�ӆ����5T3\g�k��>��q���7��`�8^9`���*[�f����~Uکg�O�p���_G��sC�_M��<�E��,6�t/��=ߢꝿU�;1���z��)d:ڬO6_���3��G�W���5=�q�f-�Il���!�Yn�6�LХ��j�l�	i�4���i���X/]'|����Й��H�O��J�����+��ݏ�����%����zކ]�t_�&Ԇ���4IYW�B�].� p�t�@�7@��ʴрU/�A�-#�:���VoB�r&ZO���9x�����x��*��F��e��z��)NŠ7�<��r�@��m��.�g8n����z+5�^���̾�k�A}p�p� Iw��1����~��v<���*�7��<{��Eŋ��@�^n"�/-5r�Y�}Y���W�h3�3 L�"*�Fn����'�:��9H�u����Rbx�_�|�g�цm������/e�d7�:�F���^�6C�Y|P����M��䆁��>�����y�Bud��{�M��05TJ�4�dp�!po�����-�Pe`v��z���ۄ����0[��(�����R�(#A���r����cH���j���K<��l��GėR��:��Tᓣ)eoҡ6�9���I����[k&��^��x��U3����%��gQ����ns� �s��(�S�s/�����K��a���.���|�����G�z��RDN��:s/�!y8r�WW�0��б���n�1',�輺������/�+���Q���Ț�Ιqe��_]�;"�;�V�<@�� =.�QQ,��g�!�2�1�yu�[�+�|l���;?6�E��.��s|�.�
����!�A����'�d[�����|$��=��CH��\�	�����[���Jg��!y[O���٢�H��_7_�VC��i\�d�ԔWz�
�����d�|�r�3�y�FJwl�.��D�E�����h��l��h�S�B7�>L~h�[?ᷟ8̙��-�.���ۏ�D��e�uҧ����=���q��P �B��X�v����hn�5P
W����Z&Y��n|���n���^��R�e;�P5�c^��եB�g.!�=�
5�y��^���(�B�8��k�(^��_���D�g���Ck�͵le�W����ս��T͔ �iȉr���T	�Y|�=
4^��F��y�O�0m��b�oq �$�f��w�!��x�4��͵��mZzO;��gF��5�
V{�.�6��+�V�a����|���{ϑb����x鷱}\�w�y��ק<UY~�J�I{; �-&>:��cLv.~�+�����+E
�0ś��p����|"�k��%cjX��a�n����U�ӋQ�[��{˪%�z�}G6��A6�����;�]a�ٌ��)8���Щ���R+��3��~�i����������r���כ�����;4� �"s{F��<;T"ŋk������=�sU�g�Ha��	�a�=�i0��@?������V\�m3�mV@b�b��Z��أ�|�����g�����E��<�O+y���j.�vi�B_��r8ד�#��s�ԇ�
��6H�䏞����p�t>���` �(Z)����2�@!��yle�C����VϷu���ک;����1&_W�.E�p�/ae���3�Uu���bX�Yt�'���+�p�-˪�����1�L�Sp��zq�ucm~��9�0���uɄ���fH����/����`���7�s������.=�;'mi��Ƀ��5�H}��Dh֨�uY]������MMP�zޑj����طN]�Ң�D�K������i��t�����ks����|�]�N>�v�+��y�î�r�1.�!��P���� q����V��B-�
vvG�#��
�:p�f�M
쫄�����Z�?�LLS&�;�00`�w��8V(m��*"� �ʪ3
����q_-%�x$��G|~5��>&�o��d�Ad8Ya� 7:�)�����/u��N�{)�]��W7���Hf�`Jk�L��#����G��̜#��D���r������:��<���wy�L3�Ïv�g���ԝ�s���5��`�7VZ�
gu<ť��y��(��1�7��-�D��Ԥn}�<5����ob�7�$�k*b�����AYo�8bi�T$��v�m@����l~F�w:5A�.R���:JqP��$�v7F#\�9�l��H"zN[����$��}�DN��5a���^�p��{���+��}��?�آ`�A��*��{e:ϯ��f�ݥB}O�|+�1]�C��A�k�(�������ŗuf�t����q��%�ɢ�9,H��0�';�+���F碹@u?Hi�+���M"c�*{w��_�s�Iq�,uLWL�o.�H������}���D��W #���!��I�U����Q�1ý��9;�E�%�_�/�d�����
u))��;+ص>(ay��z`�WVV3F}�k����5A#?���j�"���?|x�C_RXh��P۰��ț�๛���ǚ_��cA1�����K��lWJB���u�˾�)�K����qN� xOÀ"�k�?��C`��7LK�&6�:oK�W���m�����6Ԁ�]՜�T�V�4e��k�)Q8���w|#F���o���f��n��>��O'bdԬ
�YƩ�������6�m���y��Nan�@Rm�*[��2c9��d�gUw�1�N:a�Ȃ<xn�č�9G���)�������˪���$Fw��ߘL�h�-�d����?�y�4>�Xz�f�>S`���z	z�C����Xv�3�M,?Ğf��k��~��g4ط)��ˌo�����-|1Q+��<�������Z#2�P���d?�})vY�fa7]o���n����1��E�y>|I(HCl�����k�0!��G%�h���^Q)�v��ۦ:�
�!���5��k�f{J�,�tr8���(W��H���f��>^u�y�����F��0 �9�2o �8��_V�]��g�*���M
8�.���\�ۯ88C��?�Qf����#�3K\�/B��44bc���7��-K��%G��Sg�ݲ�-�8mp;h��TӞ^�}���h��i�عu�(7��cn;m��Ѝ�y]��()k'��Ω�%$�,]�C�Ƶ��_��X]�?�3�)�+����mg1���a��KY?�����ɮNŮw���^-��<8�0�?�zu9�X����yo=_i6:Qw<��d�����4Y֣���������*��ܬ(�Xj
P�t#KG��A�	�-�`,
^IR��J���'�~u��4�R0���&��u`À���'2L�8k_���lʻU�Y����n:�v*Y�W�S�K�K<��7$o�(4���<z�XA�x������[�W�e���s+˚�P��Ǹ��kQ~QE���;e�=!�'��a��͓�ҡ��#��y��ja�ȑ׸�p����~��x��i~��{��ce��说��I�U6[E,c�󾶺� л�:y�洛cߋ&���d�.T4@B�Ȁ�Ы�{�kg�I	6�@/�n����$��1)ְ�P�����A-��%k�V#��LSg�139�ku��SR�*��w�.s��p������\�$2�ZU���~B��ɌQ�N>�	r�x�_��υ���=�*\�oO�S|~�@	_��^�P�߈̮��q�u�~A=�o�\�@'������wY�cOk�#����ꎐ9Qb�QZ>#V7�>��^�i?���HrT,_?ț�W��z`������\o��l�j�7ab��w�If����w��&����d��7Nji)�$%�u4�߷���N57�{�-���׋�z�2�x�D����45�J&�f>m5�Q,�K�;�b��_h��Ƹv����vU6��Ć�>���Ԫĥ�^�aS��G^�B����`����ʺKq�C+�e���o=4��6�/�2�_�U�=jӯ^�-�r޵�����0��ۖ �p����w'8�IqZ>�����o��)�Q����xcQT_��#��k���뎓{ݷ�6�tB���{���Vs\V�{�NV(cO&����5�	F0��	�i�7�I���~N:�J`��<�2�?���?��������^�n��te�F�[��:��<����e7�gS�S0�¤]#��t%wu*�}��M��,�Y8�ߜ�We���a[�a�ȃp̃Q���ͨ�1��w���됀�^�+L��Hl��5,Fb8�2Q��A[��_x|Պ�.ʔ�i�
0�UKH:����^�l:�=6���W4����t.텕ӮO|K�UF���3u��rp�ح2Pzͷ�5x��A����ubI��RR��!�TV��CCS�9}$}���	��*���>
��c�R5(8��% �h��Y�K�SNov�����҉y�n�X$erK���-"��.�1�n�8���=8�ߎR�m�(t���
���=�Dk�w���#F9\7�D�!Q�=?� �;�4� �b1�TfƱaQ�|J��~�ZN~Q���18�^C��a+
�E,��0�cI6��<b5a��z���t_>�^V�CwYݻ:~? �2�z�R̼L}��VL��liD���=��J�q7)�k���(�eЇ(���|�E�BȧC�.2��s�ï���.zqB���D��E�����U�mԠI�=}�,��Yfү��A׏D1��/^3����0���G�8��nr�~
N�H������LGǠU�N׮�'S�`Р���8k��Fk�X��f�Dú֣���ũ8�T���e�������nY���B���Tw63P��S�X:��X5(���Z*���-���(l�v��b���e�t��L2�6�?��{��7�9�9.q���׻���3��#98��7깅��|�S>�9*޳�&e��z�6jA�K&@O�^w0AT��IPA��S��^�����\c��w����
%�EE<E��b����ɫ*���gC3����uRuQ�e蘯ʬB�����r���Q�F<�G�\�B�,���w,R���gS�k�{�1��'c¡ڔIɡe�NB}� ��kS����F�"�vh����h%F�����Ļ�-��<E��*?���ґF�/�� �p`�8�<D1$Uq�@@��qz�LF/��J��� ��B�D��ܬ�R��{��@ςv�KƲ�J��03Sõ����4g��2���;���=���=�r�\-��;ւ������_�HE���7p#F9�mݩA�����{[h������6#_�;gP�.�G�o=�Z ~�a�{~Pc��I�r��<��"���jk�~u��Q#!�9l16ȣ��I���;�*���WqX|��v�n�j��Z�p�D>�Q6N�o�
XK/�`���Z	f||$g�tx�$�9��� z&d4 :�H}#����ǭ²���T���Y�~����ɠp�gE
�����ޛ��Sݳ�l�%wF��.������b�貚��u�oK�ϖ�D'�=z�������J��m#y�B/�6��Q�"�\���r\��70�OP��Ҭ6�X_��^�g���:�_q��s�_R�2�p'/�F�I�=���Ai�{�0�"0c�����bH��Y(�l�7�K9�t1��=h��	t;�;�«)��Fa��=���iF�cmT�QN����%~��m��/#��x�Y��眝�s �/��x������č�e���e7~�x�ܶ�~����-h�uqp��<;�R��|��6豓;�P/I*��n�[����{�g��_����r[Ͷ��~�Ty̯ሪ��9��r��깾
��0.N�9��7����q1#K�.�ت��ݓL4lR��} q�����[.�i|$��<������'X,�mu��'���c�4ru�2mTƄF���S��(�E��^���J��J��B!��`������Gπ��3�M-��)� ��m)���j"�g�^X�s��w����(Hb74����i��w�a���U��ԉf�<�
�E$��1�i�����]�t��6�ݛ�_�.�s�9�d&�w�=���а�\��2!�A0��o?c|g�ډhMɷ�~��7bD�}2H�v�tv�l��<1�d�f;�<a�	�R@��8o��|�|�S� ��˝�}�tQ}��/aZI���{�&�x��eUT��?�O"M���*ل@� �����;�|UڰbL�����|I��;Z���+ ��E���_�P�d���Ė�Ie}u�}ʩ�c<Ps1#�����PO����o���cp��i3������&�ā�C�vm������W���I�%$<�YQ)ö�y)�Z��8l�}�2�R�T�h�*cXQ�M�@cq�����x�*��
����$����e�frO�KP�p�{����r���P�B3E`e�~	���pP���<���/�I�U"�ܷf;��@ͅ�!�dƐE�Ҹַ]�6�u�޳��PfS�[�H�T��T§gʭ��E	2`�&kX����sAIo��!1 P��F!�+�d��J��xc��氯m��7 �d��M�}{:{@���oB�[XZ�Uƽ0̅�6<e�\9?� ��H=_�{ �_/E6���a�����i�ͷb5(S�����qQt�ۃ� �%
�� �JJ7�"�,)a"!)ݵ����HIw� K7,������~>���s��}]���!-�9Źq!֚��F���Q�y���i�Y�e�j��-����HhI�IPS�`�����6Ԕ�Xy�	ւYR�z���ɼ�<^����s�i�4�˦�#�fV�TS�@�<�W�&c�`M�@"%�t&&���`Zsǯ� F�NN��������+֫r�VO��(|P�&SJb�|j����B����w `�K�e]&{L��%��dD�������/bU ��8(W��vN� �\��W��r��U��M��?�64�3"j�^,x�m���II�T��@5_	�����Ë���9Q����h�\�z��l@�B��#�L1��\һ��/�X1�Ӕ������g�%�����"Rw�V]����	���� fI[���ج�È�w��Óא�ߪ�
�����i���sɧx7� c�-��6F3]YK�/�G�1n�K@M22HOX�)�%��N���Q�8���seD'Q��ڇ��U�`�ϰ�t�u��CO��ʫ���@��ʟ٣�C��UV��Ǹ�h&��"sF�S���o�)��K	8r!x6��8$�ڂd	�ͥ��k7�����Ɛ��g�4	�_��?��q�Y�ɳ�1:����kyB!R��P�=|���-~��ܻC̥��!0^M�H��v+�xաX��l�ZI�v$S7�;P(	�WA�'^���g�>��	�"K<ݤ$��Eo�Y`��uͲ��;q��'��8�ix�dW���O��=�$�u�����ń�Γz<� _�\\�sU�O�m� ~��X/����e��9{�]ѯ�CU�п�S�Yzt���o��7U�W��b{�,�%1_������dI��zP��_���·6�Pg
h,{w��·W�(�:�5LP����W�2��ۤz}K��B��'�xi�< �46�K�9�}����7�U��Fzŗ�<�7ƫ�	,S��u�g���9���{0��XA��u�ax����
��K	q`쓊�sgDWn�D3J�|4�����J�?��{����)oM��չ��Ե�$$μ��7��R������k���o"��a0�F!v'hK�n�� z­.=I��@��7d� ��&7���6��f0�8j19���v{cV�����J���o�9ʍ�m��Qa��g�h�s�X�S�.H&>!ǷnN�C!���̈́� �G���Ҩ]�q�8�˗���T��x���Qcum��]%��F�ü��ݢl؀DF�X��{�Q�\��m�6�!��Ө�aD�zLf��I�|�:-TbLf�K�Eh�pD ��(��h�l��� ���?w�b�1_�M���s�l0�lb����ߣ�{F7ΙQ�ǣ�=o����(+	�X!��n��G�z`m�r�i
0��aH�v%1�H��JȊ�˟I��- �����7��k^+�}�~��Z�����-s����%{�t�MlLI�ƹ��C�<.�d��P�?��=4�!Ubm!�X4H���Eא��Wn婉�/�
��B M�5������@���Q��:�,��$�s���xHH�V��w��k��ZI�f�@Cqݤ�`HDEY��h�U�~���Y�3rfEw��x�G�)�.]
����F�7D��|1��q@�&�(��jAI+��R��V�č�%C�3���ş�� PKU��	��3�*H���^[Х4�`�R����ȧ�:���~S�������|��2�������6�MQ�t̱v�r<�j�����N�04G��\�gf�&�����:���7 �y�eR/Z$/���L���j%M�1��4�cl���v�{���
��"uxs�����
��g� d��`Y��m[��7 �|�/�J�@]M��R��[k] K8/����OH4OiiY��aϿioO�9%,�M���y��Pkz���tY8�S%,3�}yF\���E�]r����|)'&�h�g��]V����v�Gq$�B� �h՘zp�:�&T��'�庯��4ӝ��l�܎����>����r�냥�r9OG&���[;���b�@h��r���6��7l�N|���z|�h�#$�.ԓ�F?쳸vvU�_K&�������_
�ye�$��X
�r�w!�p��3=-��
Y<�u��/> ����><g�F��A���>�O�sNCB��h5�7�A�ԲC0��"��3�+�q���|H
���ѽ��=I�ck�+��``F���+ r|Dv��\?��fd�����Z� (��fp��?F��k���>�'W�ƭ6�-�,���n	H����çUU^6���6ȝ`ǫ����8����֋�fR��!���R6MY���(�:ӝ�ֵI�-~�^�Ec(fN��c�W��{��)�<&��Y{���F7�s�-��0�4���m[���a��ĝ���9��)��2�Tn���>�Zs
(�T�������� [�A�j�%B� Y.�Ӓ��qa ��H��P��v�%_)�K:d#�A����}��j��)�-��3���_��Fʻl����8���`������w�I�U��Ψ�)~9� ��i�.����?T���P��ԃ�����`@�����N��T�s�"ϡ�ְv�yc�0�!Z�hX4qՀD���,&����i~d��5�̯w$���:��:�� nϵ������l��Z����%X��X��w�B���F�4+���s˒�ͅ5|����⯬|�����?�\���ֿP�{&����b��@n0O���g7� ��<�'6ɞ�� �Rg��P~o��Ng$H����Pk�K�h�0~�0�T��gҲ����弒����W<m�x�?�4➿��\ʑ�ؤ�ƫ���h�ǈ	d�$M3�=g8i8Dww+�-
�`�D1i�ʋ��c�)C�HO*��]�C�~��>��$�u�~[
��/䄐I/*:�6J�:��(k�d3��P�� ALxD7"68�s�x$-S
�U��ȃh��eU���Ld:���.�5S�J5�L�hQmyzL�5��~D~.���,�/�k���6%U�.���橨!�,�o[��8�8aec��i �3N#�7]O� ��F�9q�D�>��έ��	h�_j�z�H�:�^�E�$�G�\���)��߄[� ��-y^��O�R5��^�7Ib	���u���bZ��n�7�����)|��d$��](���Y�0x(���4Xc����Yp�
���cNd?���{���?E�?� o�j��~�9/����s��kU����B��q2�,�PzÃ�A����H(��P� o$���8��z�9��{W�Cx>n��d�P�$G���+���/n����Ȃjz��1\�%�ɛ�1l���q��7
Y�u��K��O �'��kK\�h�*���Au[^e�����򡋏�qTI60#���Q��&4�@��h�A���|�?F� h��%v�������q`ԋLd��\a&�e8EV��W���X��&�7�5��)*���a�bpo��b��S�>�a@�_1��&ʛ����Ow��`�ÿ�ͬ䉒��E+�����d�Vt��k�L�)KY�����K�7�
��h3��` �����fv���QkmXǙ$B�����0F���C�|}�^��~�oߚ#ܯv+����Җ�AnB|���L�L�*G����h�G�ַ�YZd_.W�dlԓ�?�'` A~�ʒ}��E
�H�B	N.�[ pN��U��,*3�������:;<�(�>��P��F��5�:@e(��Dv��N����m���6v�c�BI	��T���h��H��Fens��s����S<ؐ
��o�~���N��4���t�1VO
H˗o?|�D�vU|��q�:���c�%��5�1�l�7��~d��@��־�����k^�6���!>ѽ��e�z8�%w�!9b���R�� �����kÎ>�0A�>_��?�`G���7p�(��52u�$n�~�-n�]2
�ND�����̸�p���,Vq�>��bae���b)X25	!<p�
S3J�e	^%�������x�ziD�o��*�����x��y�OP	�=���6���>��C�4>��	~��j�I��/q��Ӟ5�g���ro��yVu�Vt\z�& ��c����u�r�����
�A�:ncg`)�Zr_m/����Ƚ�G�t���~H��X*m��o'�@㿉����~��m�z����A��<NQ�Z=}P�U�s���;S�k�шLq���P0|�z��s��Uh��P�ac~�_~Γл�ZY��P*�e� �\�>n� -�FP
{���Z5?X�7J*�Өf<EPB�_�(��@��`����TS�P��%�	H\$����h@����6�q�ă �ϡ���4��������O,4#߂�������A�b�z�A ��g�x �^8�8�돜y����ޝ/�B�r�'�oui&�P�觥�)�K����3�����kk���4nL�-��H#�L��&PǕ�F�P"\�ǅ,ZA�t�Ø���0Cm���c�N��ѫjSPہ�����;��U�ux�΃Y���-�.y�K|Gw �Bɨҙ�|E��v	L�R?�;h9Y-�b��v~:��#���^��u{�w��	Ȝ}�`�[�rp_��Ǟ��B;�'p/Y[ФG8��HT�I���_�v{��qeB�A��"t������D�.`!��l!jg�������j腎C�'����n�4�c��I���x�j�D ���lp/x[}R7���.z�֝������ʐUD���<k��>Ðp*%�����p��Bkr�ZO����7�^�ϳUO
��}[��i#;h�{�F��͇Z��0��}@�1��	�Z����H!������ ��"훓@V{���f�*�w���C�E��$&p/0�X@JY���9���Y�Sk^�_�,]ĮL4���jbՐ�5���Ӳ������í���Z�g��|� G}>ힼ9� ,�S��E���r �K�6�r윑�hD�`uˏڠ �`��R���oM�mC��m��fR��{h��1�A���p2��x���M�w>}@;u�{!6�8z&�{�gn�j�G�u_��^�����1ho ��k7H)��)�Q���<Y�m��QI �Y%��~ő1\�E#vڷM#n��
�'�mS�Z�v�j8а F�jh��f=�=�ƍvEV��ނȥP���K��ܵ^�+Q^mmn'g�N!�;��>��9��C�DQ�P0HPF�ê3��KM�m0�Zn�Dռ�hr|��)�8 �
6�b=�2b)y���R&�ò��ے���'>5���4�7R�o�JEq��2x8�b�-��r)F��n&��@��x`IdjF�v�9�$���d��Df47�q`�n�اhgvw�1�*d?�x��Zൠ�!'3{Ug�ě��ຕ[�3y��l����:fY��ц��Q^��_�'�:E&=�sF=$ގ�˅��0�gn;��0b�1$��<]ᒻ�&6h`�у��c���ב�C��k��U��?o�8bޢ��T�!��"=~�;����0� `�3P2��}G�
�)�gߢx �
�
�5t�t�����[�����_M����>��x��á��ò,�OG�3-�������5�𒾗}<�����ʹ�-q��ԃ�{�\��F�#I��]���0p�W:tn׃0����N��X c�W���z�g*pt! vg�y>�Q�v{1K?�hH���L0u������W�W.����r�Pm���vKtH�F�:L0L�"�ky�6���(�g*߁jٯ!�@Vz��P�֚�e�]�����V6��-�ЌȪỻ�%�r���:fAtޞ���%�*��B�cS��1p� +O��xq]��S���EUF1�h�^d�� ?��bm:�燹#}t~��Lr��[�}���򔰞'_�Y�y�	��*��f�B<&%X�t��*��'�#��Z,�� ��e/���}�����w��g(6��1��\˼P�(�Ĥ�٬ M�_Îf�2�Ə�oJ�|0�^�g�}�d�%k8��ih��p)��t?*T���C�U�{+��Z2s�	{�F2�ȶA��@e�7X[_��mB���m���M6�@B����:/$\�C�������]����la6e��X{��I	CM�����_����������ti�[�=�Cek���T��wx��w��l]�kS�{��#�\ ���h��^�Yt�`��%8�!���M��Rێ��R�ZS�����b�y�n���r�e���{���������iǶ�)��Ǻ@�m�[Ww��li�����mt�v����B�X���������aWQ�M�!qo�$w>�Z֯{ծ��Gz`0��` R^ğ��D�������6��c��Pl��;�l��j����TE�mJPS��W�-��Vy�Hm;�ؾ	�,��Wc��Ni[�aP������&%�\��^�꺻����vLץ�|R� ��$|�]���������$s�-&��#��Տ%��J���]��E�6@2]*oaS�l����Z7ASV՝e��m��~ɯ�r�j"ɨ������r��i��p<p��J�k9�k�F�_U��xņm)	
��pcC���}׷}�I����@���ı@0�c���;�]�$ʮ�"�S��Ed�Osɘ5�	�tf�櫛�ۃA��	m�����u�&,�6�ի����<Z�~/��~�D@�ژ!�k�)i;�7^�rWp%�S�މb-"�+������JN�?yΦ�Qc5�����j�y)����폓8����Ӆ�|D�Ӻ��Z� D��y,/l�86A�|o'^�.|�=��D]�JVW4�Y��إ՞}�N;��}!dY�0*>�8��ۺpwl�����du�Q�G�J �.��q�Q�ʙ�_��ٍ����a�Q �6�S�=�v���M(�k%z���:���:�|P}`�!ɩ���Y:
`�0�!��/��<.�ٿ[q*�����
�.��R���O�5^�ҿq�h�<}�y�-c�3A7s�Щ](
�X
,���`¼,v����RϴK�/�]}
�^�7�Ć�N�]/7:�f����s����=��]ʂ�@"�o�<>�_g�8������[�A�v��w ����J����&	+|�cR��F������Y�{/�A�z)��~6�'y�b���4�?Dq����}�r��5���c�+���u���_C�D�3x��0�6�����V������a���vM�4���q����g�_*l�ksJ$;%����
@ZY�o�jxR
�[�2F9V����k~ :0���(�E�������,"͕W$��^D��;��2S�7징�ƴ��T0j3��GV{Í����o�-�����(*�%�\i�%;e:>c���H����>�4���Y�J(y:��T%�k���l��I�8"H=�p_��3���WӾWx�fQͥ4�n^*vqY�`�]u�+7}���t�]+��9��b�Ҝl��0�Z��{E��~��'�J�{�:�{�P�8�i4��o'�t�˓�w���Ffw��Y
���������#�Q>�C�4�Kcb%`<�ґ t!�?�������6��P�'�s�' �f͕���
/Ӹ������2����.�u#^���ɴ����p�O�s�[vj4�o^pH�p��Ps>\���~!���:�=�7���o����,����3\wĊl]��+�&uzh��Z��� �P����k�عoG�օ u��^Ԙu���ZF��PR´�O{Z�b!2D�"�HD����ꉮ���~�벉)�ub��XN��׻N^�����3����翯bcb��ÄU�(E�ػA�W]����?�m�ΎW��sMM~�5l<����.��w���T-}^�N��I;%�x�FN"&���w�{q;i�Ck+�\9P���o��LƑl��a<O$=�A�G�Kf?Y7�N[s�VvYg���{}I�ȡ8������i��%;x��ktq����U$�@��qR5N4�_��0���Td+�=��ʪ���D#rH6�U���q�'ve)�Sl�tI���}�}]{��6aK�����2���Ogoqş�Or'[�T��
��b���G�}�o�!A��{��'=2��s��������kL�/hw'��N�3]G�s�̞�7<\�$eP�hr��;&��>r��^�.l��V��O{�+
Qtk"�� !��i�K�����=�w�$��5Z'rF���w���!�8Wĳ��u{�rq������oq���1��B���ڂFM�/*�(��)��㬢9�hr�)VgX��{�Z���ǰ�Z�����8��Q�9�1u����Mǃ.9�+���Z�YiZ�-HUA+�k��f^u�$��V��D�������﷋Mݦ��7)�3c?F'�/&����'+E*S!|�#S��ĽmL�����'�����]ы[��z�����!��\��ϥ���E&������1��e�~E�����ʨ�JYE��+����`�s��]�����ܼ�5?�M��"U��	"E����B57 �]2S$�������R�OKW)�|L����*O�O���{���z�}�Dfo�P��Z��ؠ��h�S���N�q�ˋ��ϒ���J�.�*�q�'2����9�U'�)R���Wgm]���PE�
��Y��k=�Ǻ'� �B��{1u�z�&:�ؖ*
�8���)\�z���[}����W>��h��M�ʦ��i9Y�ͅrm���OM|
�lk�W��ck#e,"|]��f>z�R�no�z{\��:�P�63�w��$�a�rN�c�{}f �GW��8- ��v&����
�_b���T��k�5�\�7GG��h*�'��X��Y��*`f�Y��搉��HW<�Wzz8px�^�Ơ#���:�k�6⁲!۸r��g�0��� ���cփC۷=��)���L�� ��Ϣ�-X՚�2燄%���A#���<�����6)CRk[�)���?Z�nN˚�E���憓p����d_��$ke�WK�������L��w}�Y�S���ʗ.�o'��I4=T*�)H3�#.R�(����9S5ߤfH0�7]�箧X��˧��Yp.B"�ܭ4��7�F0�O)Yz9��_ zr�{���������B������!"�x�K�k^��F��D����2>�~��ge�"�ە��浢��ւ^[�c=�X�U;3S����K;I�����V�
�K1LH/�})7�ہ:6�J��h� DH(�6s�i��;�>++k������1VUQyp�|�f�%{-s�X!�,�82g��:)�^����@�y�HHC�ߑ�zu��u�Ae{�胼`#�^t��YŨ$Ի
Ԩr��	U�����gc�?�\�F-AV�C��]�b�_��SfYJT-��d,���BA{�e�Rr��:8��X�4^Pޥ:&�[f��gy�6��YP�Ց9�w �ʱ�b�Z�/�@CϨ��l�բ�4^W���Zh�U^Tn���kՑK�%K��9�?K�j �v��o����kU?�Z����G�c�G]��UvEr�����ϟ 6z��&<�9��^�Xh���4��Ͻ���EA�f�ٔ���Y"7�DezV
��R�k�T�*y�U)��n��\�����-t��=���l�}�)Sja)�z���烆����G��)�3Qz�*�3l<����L�[As%`��8��R���?0$2��$!��:�N��j?�H�j�6D��l\������./��4������:��8��K���T�\��Z#�DpN=gÃ�G��S
��f�+��x�+���?�Z|�	H�5˦���q�wϛPR��)�M2�{	?|����{!�百e�Q5|;e�H
7����d��8'I���|��k�Q.$��g����S�?�0��5b3����P�>bjI���p�~��8�����9� ��n�[�zYsQ��S�	3��5�z�
��M�{��&�0�"�S�9Ę��D��PJ�.��"�# ���Q+t�y�/p#,R�26Ϊ�pe-s��_�>���zFD�0�9	ѝ���".nzCO8D �4j�aJ��ߞ۔�.�-M���N%3	R���я��+�Y�}c�sK:�)��Wŉ��I�z@��� ����a^Ǉ?�06�f���0��6nQ-<���g>���R^j�q��`p$��r�d��W񁍰W?�(�X�7^� ��kq�1�EGH�B��.z3�.�ŷ��ĳ���U��L�B]�;J3;4��@��pWXn\���O��wM@mV��B��4\h�ta�5�#�]���x/VkJwێ���rⰵF}!`JŨj|K$x5!j�m�kC־��x����"�X���h�焝]|��?�c�ٶknz� �~^�������k�c���U�y��ٷ�E↢&�+n+/���@H�8�E�f���,7m^��������Pڱ�1=�#{� �l��kk������U��Pl���N�YجU��d_z�U�n��C~���8�M�&ƺD�u�[E;x�o���\�EÎ���&o[��(���� Z�����H(�'4����:;��Cz�wl�F)�
�mڼ�xl=*[��d)e/Ta�7/V��+IՁYY�\�`5"0�ɟ�� ��+v��[)�k'':���oKg��#��6���k��M�)MuB�/�e�o}�bϥk>�c��Kc@m6x���<昜r�wݤ�U�g��݂q�@I-��6�����\�չ��Y�U�B��'�I��肑GU��oG]��c��K����M���y�6��{6������5��K xc�6ǋI�{����}b�C_m�][4lA�4nt2�y"�ٛ��Ȁ�cӕ�SV��Q���M��Gz�й��f�v�"tw��纱"0�@W؅S·��i��f��4��^���	ѵ�;D~a=��y�����Ŧ�d-��h�K�C�>[������U����zh�D8�"�1�i\��XM:�
a"rւ�AI\��c���-���1ƫC��k�s�=?��Q�S4k�Z�����k�'	���|iԨW�N{z~
�-q�9e����~9�$`�1|%� 4t��fڷ�N�ϟ�[eg����g��f�����e�Z��7�$���f�r[ts�m�����!D��	Ԥ�:��ڷȗ�B�	�H�ӥ����+���rK�L�i��tz�\�m��GQx���_�_�R����2�&�]~\L��]����_��6�`�VHE9|xK��5h�~pB�r0_� ޶].����p���Y~09��X-w|.�����>l�M��
NktR�b������uά�����WA�������Uћ�g����#�֗�mM��ra"�!Z?���)��Tʡj���<w�s4.7�i�dI�2��,�^3%p)�Y��E�G��Z��G�ᵤ����`O�BfJ�z��`���+ů�\�--R�R7?��p�����r�~@N��3S�W|vڎP4�/�]�.?.�Ӈ�R;�a�H��?�%9�������U`_���uʴ���6��BPF �x���c^�l����?�\�)ձn�0��gX���8��y�}�Zi@��>r��ō4��)�y���
e Gm,P.�b��¶���&Fxh"�,曽���35����P��7���J����W�~��R�E���Tu�n�y_���̟�xѱ�W-��v[��ܘ��s�GZH�p��C���ٚ�qW��I0��H���A��W#?��%l�
'��&딍X��ISZ�7�?�:#J���|�Fr���J����r/<�pѵ@��l�s��UͯM�Mt��Ԕ�O
��1n�-��ؔD���b��=^`%j�2��^�M[���.{��vmk'c!u�ꔤ��O�N7t^�
:(��b6#�1���**ۙx;���!p���V��.�|������B�e��j�u�M��2Vf��E�)u�d,v���w⺙-�V��;�p�^�rxDn8>>��
����akjG�m�?Q��}���o�����v��D����M�q]�%O.{y���u5_�3b�K�8D%�}%LT+�D��${K띃K}�&�%�W�L��BQ�N���XN�ח�̕�7p�뀠�j��Shm��%�����؍GεAӗQ���΍oM%����5��iJ�"P�I9+�\_p#�D''
M*��atj>�e�s�;[��!E�'�\8�L�[��+��R��_��
�F=�SU���:��t�W�7h�	�����bA�έվʯ6nt�k����>��5�TNC6d��O��Lm��|*�j�
�����/�iČd�'~��M�O�%l��Ew���wvnR	�F/N�<�%S�viKbc�}.�Dֹ�!y����8q��ݲ����`���jͻ�S拕*���#��}O� zC��>É!l"	X=�^C3��9���3�!K� �V)��}���=���8�Cf�K�غWm���Hɛ��� ���J@1g*����LU�МzjT��$�=Ev֞�U��H-�b=�,Ǜ�!�������go%a�:�ʧ�ş<͠WlR|�FO�����|$���*'n��#%�"����D��}L.*�L�v�݊��.v�c��O�����X��ݚ�y.CY��D!|���2/Q�˽|�[o�H�j��/M�[��&�Iu7�̯,N��+�;���3�̕L��U-�D	;��H��%������Ζ�E_=O಄ ��Pq>��e�<6A7���p�pas�y�-ݺRb�Ӂ����l#�m4�O���2ꈸ2�G��;^��o�q�aS�E�:XI�I�&��:�WEg���1o45�(QY����zLa���,5Ә�E0s�����A�7Xho�ܚ]�<��̇��Gv0;��.�]�8�':�8��=�a�_M&�-���_y����P�ss"�+��>�BI��0��V#\|˩GW����ja�q�EZ�U�㘔)��"���;zgq����:Z��X�X1GE'���N� �FEk�/SM#�$�G�߉:REy�'������a��Nb]�M���*]�:�jҡ�/�%����;F�61�x�VZI������,��L�,�iX�<N���V�s��f#�6�; P���T[����	�)H���x�"P�gS?a�y�ǭ���nr���u%8�W5K_�)��h�D�f�W��7��'%a����uG��1�W�T���8(���~�餋����
,^�濒c)��1�MAF��̓lxV�ă����.��J w�l�����Z{&�8?�ؓ��}�n-))�\��^��4~��
<�I:ߙ�'�n �bno9�6Y���˖��tcپ�-!ΌNvҿ5vSSP
�~檿�8�P�C*�tй�_���Ͷ�����/��X��EWQϣ��D�9���ŵV��=��Ro�߫�ZT��j'���ά��;������|j-���g5V�*�S���VR>�����4�J�<�m�g��%�[5ι���!�����_*�2�c���l^u��t�j:%����Z[�.<cƮV���Xݫ)�V���>t�fK���L9���S�J�#�EmL������T�o5�������<\;�����9.轁pUZ\/�������~i�\O[��T���2���	�����
�a�)�ƆZ{C(%L(\�~�G���Ĉ���ߧk�b5�Ν6Y�~��rG=������P��Pbt���G��[�v/�\}�q���{�mb����"��V	v�I�S��i"��x��I�-��	�`�G�v㦾���#���k���`�=�ٔ���#���[�f���������~lɶ~c,\��1�[�u�H�"���v�RH ��@�K��rܿ�� Xo�	̷F��v�>ipn.���y��u:�����?G���覵�3���2��I�� 
釂xCS#�]���l�io�	\x98�Sm��h"���S��^.�ۆ���dc�>�|b4� g#'�2���M�q:k_�о�XLeA�����uyW����+>5Ϻ�343m�����ov�nsv6���Q�1Y\�!l�>�X<O� �� �@��X[�-�&��Y�$�} b����`A�'�=P����������݈󆧍�9�E��iM��.Y�I|��}N"r
Awbp�=����;�������O�Os�T�֫_�f�&c��f��%=����	W�NC��k|&pb�Gb5m��%΂��N}����L}��-P�����O�_�1T���k�`8�l�egz�vz��Ru����뎎mf�k����3&螓q ������Y���&�Q%�J��i�cq6,�7A4�_��l�����O��V(�_� ty��71�`��ó/?���@Ʋ�����������sT���`B��H��{}���ʴ�sA���$�"	`m	F��?�Gz��ېj,^�!����Zn��l]�T����nV��G���|6���.�1�#=ui�=���S[-ec����h�2�G!}3�G϶kS�5s��Mw�	�r�=�(��ܖ��0�����╌��}=�WI(�_~��|�b�u�δC�5h��{^�R$5�K/��oՄ��������&č�8.�:4-1.4\�}���3��g����]L8f�L`=��P˄�3a�L��7>��+��ڝ.��M�߅������k�Bd�;���ż5�}�>�`���� ���M�!zq��ztX�!]wǩ*�x7�J��U%������~��sWO�M�f"#U��C��U�:��h�=\bذ[/�����|����{ff�>iZ>�s�UyW���?7/�3�/�7 *����n8�U[q�9��oZ}6�%ηQY�G����!������J��j� c�qPv���T	_�zF�
2X�^�c�Y�7ٰ�!R�(�N��΀��ٲo5���q��vCߎx=�YŶ��i�MB��ym����~�Q��n�ӕ�,�Q� _��eBWl����L[ݔ�]������6���b���wW�Z�
�J�K��:|��t:��J��+`\EN��[L]*���vA�]�Q���e�1X����y�1��l=���)�p!�7��SE��I;H���Ƣ�;�T�T�8a{�Б!�7�f�R�ʷ�a��%uСńm�����j��u�XO5ԩ1����68 g���Mg
~PB"��Z�̟��H�A�A�����T�̐+�r)(p����dϜb�j�l�����ݶ/�t�p�峬V��O� ���V�����B5<��X�5��Z�:�e(h�i�rI%� PǄ@z�od�����N/~��{���~Y�����ʲ#�%����zD�ӟ.v�=��U%�x��wߔ<����z�i��v�+�5�'�ۯ���l�Q���sI�����M��"�b� ��M���.Q޵�˳��w�u�W��=�0�:�_GjtSL���I�Y��SF|<�2�H��h`s'�Z|?]f��o�����X�̘ޗ�)���!�����"���b���]��X#�Kf~��Z/3�S~�G����b3�Si���~�p��$��i���O�j�}/s��Xt�C���ؕ]��|��ǗV/��ocP�7���Ik�*�xG��S;���9�,�H:6�t�O�*Vܿ��iWJ��)d������n�i+7(x����>����Ӳ�x�Ԡ��֨�)l����;".�7[�/��7%7�ۺ�y����<Yߪޅo���y�7Z&�c�}�CW>���h'c]��rź�RbdT��J���C��z��鶝�`���,�U�e�Tb7�Z���c� ��i@#(��f�ӏ�/f��S}u+F�$�����3���ː�w��~�Ǳ�ZN�[��o�7�EY���۾$-�PJ1X����q8��n����ka��C�4�H�d�o.2�Z�`R�_ˠ 1X�1��A��W��D�>�ue�`a��`m���e�xR���#�_�/l��xC�c��m�6��I��/������,D�	d����]���5�}�����i*�H��S>����4��B�z��^��q����~�ؔ�8<~����[φ<��iB���m�+�),sc�dLե����uQ�9�8�;�P�l���Ŝ!��~�t%�8�����%��^�<�Ϙ�z���!4Ҽk��-���D�x+�}����Д���9�"qY���9�@
��<U���>n��`�A��֨�~Fqn[[p�@��-����Q��nn�me>������g���_G��6#n�������r� )��Md����9827w7�@�}]�1S���	'G��e��BwX���Œq�]��e����%���0�V+�ǥ�4B��o��K��P�c�7�`ش�����3r��{�ߟ��������Yf��J���ħtl���0�P�v��7⾡��"���w�m`-���YYuD�7{�x͌0���g<�g?�"O�M�|��O��K�'@���S��yp��K6Q�^;r:��l��.���h�W�$朠�F.�b/����t�1}\Z5�
��Ð_&��fsRGzD���>�Ҽ��#�@.��u���v%�gI�ƛ�_ e�����R��ɢ]������r�I�y���B�e̟WU�i�Hl���\�����^noWU�,i�v��Iąi�1�WW�����T}��Qr!���׏�4B�N�Ib�֥��]fwB�NĽ/�������^R�	f���Yy�X��?|�O+S��1b��?��y���3}�~�]�6^<(Er+D���{h�J�KFJ�v~�v��W��� ��`�'��)4+��F>������"	�r�VV�j�S� ���u<��c�N��R~bb(4��.�X�gHj]�f�~��en��[۴��'sx�ç��-�h"�B�C��:��������4�A����]���kC��ǐ,F��u�aU�_� "H7@��n)�i�n%��;9t���[��A�����������3����k���Qn�n��������W� �<�K;��,��$h��еh�T,��Oሟ�2-�큯��-ꟹ}���nѨ�0����E��Tx��`D��-����r�C�6t�-�r�����-��m� �&u���u,�W��_0�bc�g�۫��9�=	f�6[�$-ILM����b�x#q���"悘f�rh��- �@לfúF���TL� ����%��ȃ����$���P7���ƖQ� �w%g_��y�݊~�*1�Pͻ���cf?I�~�U�z�"��|����Ƽ�G��~�����TOݬ�v�n�x�:"`���U�wR ��	�?��	�	���T0�� ��u�z���� �۞@ˏ��f�c�n��F���B�L�Fd�x��Wab��WO����L���G�u�g��>�Ir�[�,Q-!��I�6��BC�ݨJ������)���=Ꝣ:���X9��*Y���>��*�ʬ����X����e`��Ʒ���D_�ԟ�����,��� �~�����q�m)$<�&��~0�S�L�x�P��GKv�N�s���%F�}¼o ����pdy>W��!�k�?�ɰ�������~�-D��ӈ���t(]�+0pw`�zy;�d�{��������7��=�z�7��#��ʾ�O������ҕg(k�P��j�$`n��I�>�����{�;)W� �(�c5da;1���a��e-�,Lf�OC+	��no|J܁D�
1�+dF[�;]+���\G�HFsu���^G��&���-�&�z�rdh�=p�]���j�0�U��[�����k ��8�b�;�<��n�s��gٿ����������<M"��%��N6��?��v?v<�Xu�#ܡ��]���{��L>� �5}�T�pʵ�<����7��0z�)��l6�e��'���M,,>��i�$@Y.O ?~D��^� c{�K�ݛ����S7�7�/����K3�;�M�����Ht���'t�����aK/]�c�)r�����"�IfڱIC~s��ݠ�K�r����?�$�xR�5kOY�h�^�A�*����G������;ʭN�7*un9y��� ���$m���iQX� �������G��цS��Z
WA��������3�&~S%���6��O��� T�i{��>��I`Kk*��^�3C�B�lc�O�TE�=�ۤN�hGP��φ-꽓z�]�P�b���O#�3a~�Ԭ��8f�5K�j��2�\60��M�)(�;�D�5r �7� t�p'�0R�O��l=��x�n�;E'�'���'���������9` �Ϻ�1��L��j��֡P���'l��%h��$���I��Nk��~�Ӭ�͹� _&�=%g��!Z��n����4z�>C,.M��X#׳����D}Y1���<X|�"��6J-K�vA6Sy�Y(�����v��eo���HA躚��e)G(�L�.����LY�|zQ�;�v~=�=_��؜�ۡ@^;N�n���?�Q�����c}�X��J����r����_�O��g��3~&��HA��,b(˸�R��В�e<_��fzhz�GA�t˥�cCZ�G� U��iM���a`g�<sGr��0!~<��߀��M<C�=�����S��������0y��>�8��M���P����X�c\ ��y��D��,Ja�_vھ�n�j��1�fQ�_�o�$L��Xj�b�3Ѷz��^W_����Ir�&�t����O@�.	���x�c��̮�h�U�zr�<є�����}W��J�{��" W��$2�,�ҿ��)�H�����Ν��i��q��PP��pHmc~�CV�Cwn@K�#����ћҩ��B��N��t${��������ˮ���c|D�E�� ����4�x]�	������UӪ�d�~M����Yea���Y���"����ߪ����1��60�����(=5�=mN`6��$m!���ϭ��1N�9B�V2V죗��z�9��g
��ǧ�3�hl��ƴ☕�}�;L��#��xXiq�W�0��R�F?c)V�A=<R�C�2�v
;)����5MA`h�>�O��5��[������^�=>�X20jN�o[�R:��.����%l'zy��&���6|Ì�o}����@�} $���Qko��e����j�Nʯ�5M�*�
#���~"�<zk��݌	,����L���5K��<U0�2`t;M���Ҳ~�D 9��nD�o�g���t]���j1XKu
���N�/ݛ.����`;��ǖ�0o�c�_��o���L5Nl�d�L�\ !���!0�$i�NćY��?���Ȼ`-�a��%��t|�.����Q�x�O��m��>�a&���U��Y�40@���7�(��?��^G��m71[!乩�k'h���׮0H������%�`��rm3s��Sכ�W�p([t�	�ƵU�<�����TMm�=>�⹻�N�� ��|��6�.~И��Q�G����u�R:�~���=^�hX�U���R0U�p=�EK�_aX��|�A �yt��:p�|�Q�T�����@Gf{����<�:�q�և�b����[�2�CﳻR��FK�H_D��� �6�k�����k��Km$ v��R�I(ąϋNh6�ʱ3���_�9+��zxG%��/8�~|eS�<���*�  H�u(��!ˁF��b ]z2`�H�ȱ��81����3�-��=�;��9:�ߗ�$rt����۵�Q��q�˫&U �hU���)��+�PY�92�Ѫ\�{I�߅wH
��Ī=���% }�[w��}�*S����$V�8��
N�vu�m�C��9<�մ�TY97@�4�P���ּ�K/6�ּ��۴��(�Ċ��a��P�qV��E.'
�4�ږ�?�@%�{
l���	��k�rZ��D��9=��"@��+���W@��p ���)��߹�z@~/�tD��)�03��N��t��?���_���E���U�~��K�v��6���m�>p���;�Ѷ��[��H�'�2C��+n�⟔~5͢��p�/�u�������!�
��k������\I��8��y�I�!���Y�����/�W���`��%NW�`v����{��*�C~� U�ǚU�����wA��/��� i�j������5�����֯%9�*�&�|�S�a����΀�=M���w�A�~M��7i&�$�b3"�`{�����c`~�=���/D�~����
�X�R$��ơH���8�c=�Q�?��H���U53fOf"7o �4������f�U�4��YJ)��E�Ԏ�ݯ@�o>>5+����U<�:��������W���I·�������ം�w���8N;{6w@6(x�x���c=� e~DɈ#��X�73�k׏� �0�Hj�<�u��U�JG�9?�����{�;0�(5W�х�Ч%)��-�ߵ |5ͫ���'��O��q�Ӌ��>�?�1��l@�Ƽ �.� ���&�Љ���e%_μ���BfH������.��4��%�V	��J�)�w5g�,�4�T;d������O4 gMQ�.���Ȍ�N��5�<f�����{ó��>s�>�:n�Á�/Ȁ
c�T[�{Z�-�	 ��21R7�R�c�,+{�7z�3`h�.���h@�g&��o�7�4Ne:���RzMm*�E@d�C
�����i{~\�U����aa�2@�J�l�� �/Y?Ji���b�2X
6� я��/�(�M43:I���4m@�
��~8G��w��K�=;���Ӻ5�q��)����` P���7ˆ���[��F<��0u�w�P	���
�;'�V�L⦡��s��5V�&ǆ&�9��(@3�<궉qD���|A9�+�V�ɕ�w��Z��I=�����B9���ə_6R��\r�[gzU)3\�hz�����jg�Y���R޶ʁ��AE�A��;\]���x�n ��G|l�(V_fQt@V�z�ޢ	T�ez���_��l_�O�p�!�7���MB�6|=�S?&��R�q9�{�r��u�p�8����EL��h�+U�V�l��|� zRly��c�7\2��`��8U�/�����cϟ �/�=_��&!t����>Ia���V]rf�=X����b�s�l[�|�x��a!��^���p���N5P�?;O��ָ�����*?�iy-C3<CG"}g')m�����wQ����]\<��u��� �0�J�ϋ��I�lWR��º!mb踩sT�|>�LvW#�jB|��w߀9'��'�;�$_t����#j������DT��':���P����M��j�N�J�̂/�b��O���R��kP���?"$����ׄt�|w��{�쪵��I�h���v���_��v�#�5����o�-�oH��{NH�B�Z �()Z�d�(q��V��Fy2XU1_�3HOwO�
�҆q|��#Lމ�ta!q_��$3�T�N��}=���t��	psǄ��= P�Z1�7D ����n8�����G�;��K<`��}.����ӓ)�(���թ�~�I+�L��	�݌���/vE�~�AOF;�pEGBX�:����F�� �dO�=�>@����ٮq��.8�@Kj�3�B� s�mN�����I��RD)1�����0�FB�>�4	1���!�P�I���?�8�A*;��i��|ı٤�b��R_������L��e�iHc���rѸM?�g��H��*��r$���_a�l0�W�B�����8�丫$�����oY��Ot��`<�G��H&���p]�
��o���w�X?�g��R1D�D�Tdg�@=�,�9�p���k䬯~��������}�Х�B��죥�(��t�:ŭ�C��E��VM˻�:x:?j�X�&�;v�`��B_x�sa\���?����s)����G�(*��������s�.+������#4�œo��3��O�����CX<x�d��M�&�M��DmWHu,�a���M OG�앒$�d�u�\�,b6c�&�H;��#S?�Ep�v�c>{e�G��?�s�E8'�F�Oh���X�d�ѬbC2����#����>�j)��}e'�����"��n#IX���9"5�&��l��i���Op�R�0&6 {=8���؈�¨gDd�g�H���O�w��z�uhK4���?�u�T.g+�3ƃ�ƻY�g�eb��~{�N���"&s���p2B�	(��
~� ��~�����-���1��˒��������V*m�]2��C�7�Ρ4���ٵEZ�a���U���O�S�o��n�^_���96c�>��� 0'}�,�slW�U�4|�<K���޽��M?>��`�����©)R�EL %�L}�1�<@�j�0A<Q�Uڇd
����3�� ����LfJJ�X�;T�ނaw��w	w9�k_�w���q"�10څ;�ΔGx߷����]�����<=��)�M�������8x�j�I�Q���;_��~�CY]4HYP#8�k�EV�꺡�߼M��~c��k��{�<y Q����\���"z�t1�:�u�)�y��w����JA:�=	���f��>��f�?�8�5�o&��ږOR���tS}25����o!�M{�/F���R��޻6D����	�f�u_a3��˩H���� LʊR��w����R*~�ԝ\��yFi����A�Vp$���x�uD�"ߤ� �:�pPTuc���P���A#?ׅvQ\^�0�)%�-���(% �.Y'��\����`B|�l��㐱sz 1��_�OD�ǹ`X�/IG4Ғ�j �R�ɫ���j����&Omj��q-�<�XY�:!th5�T��O9FZ;���h_9�s��<������'���/��E�R�O7�.,u痘J��a��m 6u_"�pVuZOήѸ�E��sK����ބ�R<�5�7ࡃv��')xG|�,%��?F�h7����|�0!hQ��b��R��j�8�U���ߧ��m��{��1��g�+�$��{\3k�c 畫P\���""~g=�W���R{��Ud�����k������M��T����lB:��;?#�,��z�O&����Yfa}�\,k�D���*�m���FL[�(����5�l*��SLF:^���D��%����40�t�G����$�Wy��V���G�)9f�-!EGd��Y/'B��/WC���I��N!Q�|�}��������0��e�0�5ea���%*���Mi���J�tY����`��['��lF�|� `���(Ǆ�}�4 �:��ж�i7��=Q�������R��wv1ט���H�|�ҁ?͈�e/��mX�9�ڦ�x9�{��K@&�,�,��'��m�KO��4��5{ �(�',��˩�|j6\lVk�a�?,�;;G�P�S��/_ ��0qE*�b��Akx��g}���*���
Ӛ=p1~�g�@Y�z�]8\�6�i�/��Ã!fp��X��nώ� �i��!(��������Ys�4�iĿ%�/�z��g�t�[wb�I��?1R�k�d��Ab
�E�I'�D��ͅA��.d� ۲�C���O`�߶L���������r���F)	)=dh�F����d7o�r�Yʹw��aA���i�\H�QU�����%�������;��+5���^��g�
��7��K��ހ����()_X�K�#Xdoj��}]1
��YXy��2ā���(8��+�f#�NF�9K3!kg�
���oA-��`�����}�A��	��F�st��*��p�����:/x5ł�M�)%t�PJGO{?��9W�*p]L�юԘ[�����O��o��YV�젃@1�\J�U��,�dԒgTf��tJ?�悼����U!u��m�٧��������.��Y��T�C�B���G�f��v33���F�?5tHԓ��7�S��P�"��Np�rG35�`�&i-N�w~���y��J�BK��m�u��N/l�"6cE>^�1Ȃ�����X>�)HVA�G��e��:���,�75�&`����!��S��sr� l��x:|ʫJ����WD�V��$@�O��d��W�v?;o��Eڶ����2Ƽ
7h�#� #�c��"��� ��AJ���mX���K����ѥ�Q!팋pA�۵�%%Ԕ��RVH���=ղ�-�|�N�S-�-�+xx�H9���3{����س
;v�H��<tl��!��'�,.էFS v/�'�#��p;�n4�j������X�����%���|U-�� �����).+>���8�����t�>"��x���@�,���`�F 쌲�Ne�%���;�d�ibA_�/�0���O����oQO\((���v	��#���X�`��L��������e����;� LQe$6�Y>XO�ݯiD�As��xQ�aő�e���ؓ���M�A�wQmvz����*�#�iRԕ�Y'�G��M��F���o��Xmz:g�*�T���H��ֺ��wdE�.�X�v(����Y�ȼQS�]u�0qA�MCz���V�o	2��:k�p����M��F<E��@<�<O���,l���?�ԕ�иY� �V�#�ŭ[�Pl����`ZZ�,O\r��˕8MV��ޮ��6ёB�oRi98���9�}�{yO?�Sm^����@��W�����y���M��9�̖�V�0>iIN��Bv��'��Q���z�P�����
5z�"�?�}@9�u�s��d+�X�s�7Y�O,ĊϻłU��Z��SV)��#�vc�`!��.�*�`z#~�,k�~N	'%1�y�y�tJ\tV_��qZ����q:��ld`<����ǱJ�kSE���ɵa�a��wˏ/p��q�� G�=�?��p��!��-I����>��h��Of�Z��l��ܜxr��>�y�^��g\��1[�W��c��i�m�wP8L���׆ƹt��)�H�>  �������SL�Wk��E�=��H��L �%���Ը]��»�d��|-~���C0M�B������\>�S:�(������v��y�Q3A;��)�����$���ƀe>u5�<@�֔F�
`���|Cs�Ҕ��j�%�Q��c��e�'='�2k��+��1���e���:���1�"�� ���k�������dS��Z�f�n�y5�� fo�چ�ln�_���]��>�z^۫H1G�z�z��9L D1��2W�U���Q�|��]��(;�x����Cx|���1����SG(`�}�za���f�"V���E)��W�p[O����hr��jR&���H��)�Wjj�]�����G!äo{�;~+���
�B�N�@	f@�_uv}=�L*AJf��_aw��]E�0��������ļ�C:��+�P�SS2��>a�T0|�;Й)�s���de𛬔�>r���H�Ɨ��+C�d���`	@�ڝ�s�Ưt9'\6�ę�a>+��C$���wHo�����'�s@�M,���vV�����
f�����O����@|�U@QN�މZljh�n�+l�*�S��Nrjl�0���F� �ȝ
��No&��� Ǥ*����lV�m��a ��K��́Oy����޹[~���-��x����<lFD4��q��B���틣�G9
�Y�q)6V����}AB�Ч�28�l ��͹8
�74I����
V_}������P𪞫�2�7/�g@��ԏ�^��4*6���V��L��qp�R�'�J���TI�=��5wf~oon�i��������ne������7�T�g�-�(E�)��Ww�-�M,1�q�߷ӽD�U��m-�ҏ�ҏ�����|`:�HW�qrdU�P� �ff������H�]����F��n��x���a��]�"��5�-H�|����܃�J��27�)��9��We�EH��S�d 
���S�)hp�������O����s���S��h��p��f.Jcl���7�|0�"n��&��dM�O�=^��#Pp���66�lL��_�\�f8�$l&-o6+
%9E�x�!q�Y��,�ۓ�{�lD���r��ltw��Hw��.�	����?j�Ǚе�+�}\XH���i�C�t�!�B+tZ��?�0���T(����J�#;?�&����\e�����AFj�D���=��)H,�-
j���UR~e��t�6�J����8|<�tFo�]3Ézt9�;P���{`��XQ�WvR����!�
0���>w
<RR�P�ֵ
Dod¿�#>T6���q��c]���(������ͦ�g�ݎ��e]�ŚfO��XLz�ErES	��f"�#�~�����'@��3���:��%�/$�@yaU��[���;��w�����]bz��<�X�<����n'�k��%�Gv��G�T��ЛE��{w~>��$�@Z�.�0rE]��U�<����ݡ;�YD�|K�Y�ݦ�:ֽ2o� �"-��]�E�@k����Dn��"_}�^"ʶ2����J0Yg:���Յ�m��r�{|7qP�#v����ʗ�?�{����~Tp��b�b��RW�����.F�m},"��:����b���
N~�P��
m5 da��M/x�[wn1˦���G&�*hT a���5 ���4��'|��.ܬ~<���Us�eR!�Gc�Dur��%N[1ɀ�����W�e��u�b���{�#&���rƏ��#D ��� ��EQA���Ua�z�������1�4�l�۩��v��&��#Ne檭Pej�]��@��`��"�*��9*�0��w:K+����@TD�U�����y�p#�G�#���ĉ������$(bÍ����ThSMmB_�UO�9Wu��f�:�MN_My���G揑S��F3�Ǐ�����Ϲ;��i�ɠAf�Rk�9�kP��N&�L�����x�R�åF��vd��}ڹ+����?��x^��؏�ӡ��ް:"�:+1e=,�;��^����@�V��� 4��;����?�E(n��7�����k7	��:�ؠ+)w�^�b+��cT��
>T��9�Q���Ѧ�._A�'?�iQf�ی���p���>����2��G B�0�Q����#��#j�o�����4ړ
P��R�����B�4k=��]Zq�2��h�OP��(x �'~�%ޅ58�:��Mػ�����P�i1
'
i��*?�m�yc�V��p�e�f@~�\��e�/-��@l,����&4z%go�A�:���>\&<!"���P�� jmj�����Q�ȫ�~(�`װ�k�{@�Na`��Qߑ�:��J�%�z��  �G�Dk
"�m���ԇ{���v_p��5��1��d��4�d�@Y���M���m�ǩ	zc���$9P#�Cƴ$����Y�T�t����7�/@��'W�Λ�S`G�tK��.')ˋ<��'So�X�%.�NȀx��jǂ���H��F%���w.J|;�C�
��)n���s ���%K�aXA{6�aLB����i����b(3E�yz�)i�%�Pd��"��0����o5��)�]��P���hLɤ�]�@m�wye�b�hM
��F���V���9] E؄ ����u[J@7�lĴ'�a��z�s��;�7�%d�>��ϛ��$I��D�X\�8*)H	�1|i>J$_T�ٶ���fM�)��L�g�(BW����IB� �*�
��y\��  �7"7�lH���
��@�l(%�ڭW���`��	�ڟ��Ek��d�>ɯ4l[\���������j��f���^����ŁT�[MB5n���H&���:%��Л��G�L4��p�IU�����id��U�b�u� ����$e/�����7o���r���*+@�|��B.~.�c�8�9�F�$�Tf`8��MB��w�P�br]GY�H�g�Uk�_^�����^�(�C�ĥi��kFnYy�����_y8&��w���W��ع��<��F������xM��Oz���?�86�R�_'>���������2�/)!O
�	�'j<#��ۮ������<b1xY�S��*�fǝ0�+�R%���_U}�:A/�K|JC�ˉ8�mm̀��m&k�`����wadÖ��#N]c�~��y7�4�u��턃�EZ��J�̀qQ�.�@<�SF�˦;�h��S	(��dyo,�ྗZ	��9��4�A%g���i߸��j=�uD��`3��@"?c��}��vu�<J��Ԭ;ѷ]Z�>��i�s�C�^U��|�/�k���'�aߖ���R�t���R��ovo�/^m+��f�u��ja�Ɉ�wA���"(���\���'�~dŷ.��<�6䳿C�����$U�p�e>�w?'�=�V�����Ɇ��Z(}͋[�M���B^��R�x���ë���,������k)5��n�L���.>4q�.�G���b�����¤W��4ͯTҪ����5�I/K�����5e�w;��v��>+vI���E���UpPu�K0H�e~+��T�jGBG�����X{���	z��3	�؛B�0��AI� ZR�Sr���+B5���<)�ϸ�0�dTRN��5��捎�x9�n���W����f�4���k�f��=3EPFkU_�g��m�]�u�*7�I��S�t����GE�/�z�d�ob���3����%S��LS(D<7�"<VK1H|�׎�6�_�9`��uNk)g��><�@�X��ߔ�sE�_���Ӱp&�u�لZAd\�${�M�����i�#7����J�Z�g�= ��u�"<�[��������F�:������iȼ�͉Q�V������w�}t�4���z?�N��t����.}=}��f����>�F�7q���U���-��Y�멲��Ǖ���*�ǎ�Mk�+-ʡ��=��d������}�~j ZRj�;����;u����X(|�K��!Q�1��0-�L�{gBTH�b}８�\�����'�k��7�;�G�hT5w�Q������H��t����P]�h��P�n�/0o�뇭c�(l��;����o+��lV�V� ���>���n�qBxL_�Ff�ɉ4 �KFr�Lj'8O�W��]�՞���hK�y\E�.n"��2���m��^�����������D3<����rd1�|��_�c�<˫-v�UP�*�B��o��=�{%�����~�P��V�/�}�$F���;�<E�_�=Y#��������nm"�S������_�\����b����E�{��l���s�I��\Kr�`�2�uq*����ڂ Hk����u�	6�ڂ�ػ9��*���S�*x���9��R֮��xM��{I\��M�w���)��斪�磶l+Knq���"��XK���#�Sb>���6=�ɱ��B���u]�P��7m�Az2cb<���߷�H�Zy��SJRR�"��/���N/��4�>9C��5�˺@5��[�w_��l���仅������|o7�3(Ȣ�c['D��jb�e\0��ɯ<,�-2Ɗ��w������g�j�i�M����3{=���>ҡ�&z��Kv�h�F�҂<]kY$�UF�:|p�B<m��106�:e�z�����(�0�6�L7�F��n���S�{NL����X͑:�s���F�9�
u�|Пۙc��G�S�M=�>%8��Ļ��i�#��v�A��pV���r٢��ӄCڬ�٭l��b=��R��_Fճ�zvϢ�g��z��.�i�g�������Bh�m��{�G�D���%P$��8L���
w�S��g�˒F��{/�̙�]<h��ر��f�&�]5�oC�|�	ȥs9��VT�������q���������G|�z�m��8�������/r�ȝ]lZ��
�珉�'�~n�?�U��`ɕP�6��G3"A�T�/�~�1�V�`&�[�~�r>�
@����xD�v&�`��0�ąO��E\N�'�`gc�[�:$���F[Gwx�C3ԕkl�R��C���>z��������>�Վ�M�K���h#����2� �u���`�o���7�t�ʳ.��{�h�;��S��+I��Ѓ��e�����ܐ�g-Ȯ���B�},E��9.˸Re\�и��R��˼��T�}|�t���ӱ����㗙x(���
�U�p�(h��c\s���c�04K�:����<����Ւ�(~�7�=�>�r�B��[?ەB^\���?f-Էu�o��IP3�s�yU�.������[?gLt6�3$�������G�@7���<�f3��5���[~����z��	��J:�tU㇂�����Źz��Z���0�Cm�h�O	:RM/��2���_�A\>7լ��1I����g�u�>{˓��Ia�Ǥ��'eo>m�o]�)��y��br[k0J�?�g�\�A�8��][i�AJ�J��=ڟ�䆔�[3��8�C Ay��"��bF�(=G9����(>��;n݉��#��H3v��K���B9�P�N�;����d/o:j�Rw�xSYhĢ2���tl�nHcUX���݉���K�t'�Z����P:�2�w׈~�:^��8�/��&XE��Yc�-{���i��\ѣ���xS�g�$��͹��Y�4b#«�D�ݒ���J��5��٦���6I�����ȉ �N�������t�C��z4��w*ċq�#y=�ǜ�z/n{N� *��]��F�-YT�^�ˌ�qS���{�/�9ʋ�=�D�O^��V{��b(�PP[)^[����)����	(PE��H�`�v%T3��/N���o���	,�*����Ȓ���>zъ=1�J�\Y��e'30S��?��dƎ,~�" Z<t)�k^y�i�
0Wإ7�k��)����r����Sc�pl�WLs�.��j3��.?];ѽ<�Xle L_ݪ��4ȻSf#5B>/�&���X�I�]�R�a�ʜ�C����P��w�f@�^�?��BlY~�'���\�h��]��"��6���ʤ9|ns�Q��D��De�;�a����ؕe?����(�?��"rĆȜ�T�֭��m�sCIo�Ȫx;:�'��R�X���3"Wƚ�N�\I��UV)��kR��<� ����j���:���v:���S�L�������W��w��^�Ո��O{�/mM8-o����O\�	Q1$�Ë��шTqb�:�ٍ�N�8�Qac/{4���w��d-�A�2�h۝��UxT���2��N��}�+��Z���ZPM���%��j��$ҋ!�n���~;��%�Lak<K�򪓨%�ޝ�*n�b
�L�����NT��ȍ9�a���\��:&�l],a}qW����?�;ڷ	�����H'4�u�y�wt��/��Il�W&7�#�s�x��U��	���	�un �a/[��#]tJ�/��G#����!0�}k2�S��ͯzY	�&U�.X�Iuh!�i�+U��Z~��#��,�p�T5;y\i��|�<�}@N{|�
]�r?g��B=�r潌��!��P���鎭2��s;$'&�t[<Sa�U]�+R��cZ�-���6�h�8X	Ce���	����d���Sǉ/j�u�i-��s��tO�kH�i�Be�ߑ������,���;���ߧ`��5�iӖ좹�����pn����PHV�ҟ���!��S�RŔ)6pۅ��h���b�	�p��#"W��#!�d��\[��k�������	zz89����_/��,g�N�=.��R��R�¢�֏6�1���K�����С$k[j��N1���F�C����O�)�tJ&@�!�¡_+Q�&���j���f��f�<������:R�>�~a�P��o���T�Z�,��pwe=RoHW�U�Ђ�T����C�g���%&޻�o�$u�ds��Ea�)��4�0�.u��9ؗϖU�����1���W���gs$��X{�Wڇ'�+�>��y��W��-S�:�׵j�7���!�:_N�*�Z������YH�2���|4��r}O�i!���1�q�>E�^��c�hq�wڌ@������R�'���3ə	��p� ����ԉXa����7��b�vɓ�e�X����O�L坬�������f�!��H#8\�ULMTG�+�C!o�1-3�F-��H`�M�h��#y����4G����^E��2����e���G�50Nع��7�c�΢ӕ�\����M_�=�����N���7�c�D�m�+$��,(6�6�[z��w$���l���$J�7�{�+��q91��^�iV��k���ap?J{^���4�%g���Da"�;jͨ`dH���؁�G���G\��4٣Ȓ��Q�G�-/j�tf�%}��Ǧ>���x��O1{;ߙi�
��_/�C����ug�T���a�{�/�P�����������)]�2W��������C��%20L��bb/�/�2�p w�娿�3�e�*�R ,p8]HCۚa�l�xw�$b��!��=`�������1�o$A�D���*���IȚ����Z=t+˦�"���䗆�!�%-&��XѦ�agQ��}��Q���> <��� ��G-`se��l�B��օp�e@6T����h�Å ����2�[��2r#�#
�,mp�Z�t�O Aqe�"��c�s2&��>�[�������\�z���	��R��}�6��3��XN~�>޶��]oz.��p"�J�����V�n<�L��v�����Pk�V/�����Ҏ�z�E:�4�erC�8-�OJ�b��2x�/z�
Ͱ�Ŷ���g~�0�4�<I�;q�{2V�Dj�a�i_7	Q߾���b���ʲFޜ��\�F��R+j�@ A��W�)KM�<i���޵�d���duJ��V�̋�������<��m���s��\e�\R�tl�����QRR��k ?�r$Vyl�@e�:dd!���Oh?ͩI�g�8�s#�Er�A�&��S���+{S���8>�
9Q��1��+Z���x��������t��Q0�i!�����V��d�z�涴Ė��:��V�s/<��N����A?k}���:Y�y�zפyӯJ�9���'���Ӿ�K�nǑJQ��T����x�iQ�������*�	���Y�'����kC���Ƿo�T'ၶ���p�����!9��K�l�_�٫!�"����Ԥ`����&@/T��exq��oȭ�N=Hl� -S6���0�J٥�)[���%=�������8����S��+SLV�!��)��%!�VQ�!��6��5��sE#ǵ}��:ޙ���k������KJ8�v�3�v�
��׌��٫��lj�g�������-?+�[����J���˻�$~-�%��-���_����N�4��j�^�7����㾩�PEv/��+���O#�B?��v�4�17I��8G���D�mex�n"�4����[��������%�(��Z\�,����^�r}�&Mn��6>澯�8CO��:�
�n`��!�V�-*��|�0=�����y�s�?q�{���R���_��k�0T#ޅq�ƥ�|�$7�r,��`���_�sF�`T!��Ý��]ա�`Eٴn��a�u�1ػ;]����(����､-���z����|����R�X���7΄�lbyŏ��7��~e�s�D����H�p`�l_2�y��O�sݹs(l(@�h�v��a�%as>��3	v�f<�\oqA�ށW)oR|y�x���w�1�ьpcs!=5��G��4��
}����t�RN���Ҟ��s�����AZ�šV�%����I-Ӯ|�D�tl���ȭ�W�V�����"�G���T��w�����z�A���5�ʁ�h��TΟ
u<@ma<l\t���wO1����]X�󩋝꟩��i�8�!R�������?�2,��{{ i�n)A�n	E��:FDR���p���!d��;�3���_�_$�^{�uǚ�9���������.�鲹~:���ʪ�����/��ɠS�y8��R�g�%4�VN��5}��\`�S{3�(�8W����E���v�*9���E.V��;dv���)^g0j��R��:aG%����A�P���P�^��� �+?�+�e� ~�:g�� ���N�Q�;,d^���PvE�bW �]Q]����>P�n�E�I4�}����h�<���%�w���N���K�%|�"����pbW*�zB��@�u��ɐ}[j$���o�U彅����uSCtV���37�f���z�
rn<���g1�ȴj�=����D?C88�{\�G��ۀ:}'��>�s,�䁎Y��] )e�Y�V~7"���e���Ϫ	��L����^��p��-�HCh���u(s�	q��s������c���Z[v��.�]���w��P[��k��I[b]X���L�+A`�,s�{E�`˙�쩰`�9�w2�q��[2:�B�#�r�q?�6}^�^v�.E������oK���g����a�{�fJS��
�������=��|<?�-x�VAs����ճ�vGu�8&�2� 2vF2��U�@��;���X����|�J�ħK�z�����y5��3^���l��H�!),�h�E����1S�dH��.t]F�+ey�(ſ
r �6�9Lr�����Lt����s�I��;ě�h=o2ء�}�vW�_�3��~�������:*�x�J�.��?�O$�L�YM��.�;��\	���1�;/�9���i¢�k����	#ƊV47��D��/_���[l�n�AFs�x};ᬇ>����S��4�]X��i�u�|ѽC^^�kG��3r�/8T����=�Jγ��@2���3�D�A]�c�!˺�+zkB�ì�*|w����)R�M�*,��fO�+��V���&�+@+ˍ�
[xH� ��^��<�֞B
-��dU�[��w����ſrpV�����w�q�i�W�SF��~3^�H�l��QR�G�+d,����߿�8��/,�_B(ܮt�����7j��Z��a������{�M��.V�ُ�OS��%�V�*��+�g'!X��jk�>4�绂o)�،~q���H�AZ�aL�5�Jxf\�ט�t�	�J݀^|ы9�GP����ge�ɬ�<�8�yQN}1.)���OD�hd�Z�p�Ob�W�22̕(��,��P�ײ1-����|��:�A��t���1�paC�7�e�@�2�k�(	�W!�2f��ڰSY=�$��~f���-7��ظ�h�p���yq���%���H�E��j
ǒ$נ�Ǭ��$*z�y6H���_���M�їlu�Dm���p�IvZ�M���0�"D4	�K�xɈ������i�X����L]8�}��Ҋ��WOp蒅��0�R���ߔe�vp Z���^X͉�y{ǊDa\Pҷ�5�<��G�9��~O�A�
� �蔐fh�u�-`�Ȏ�ʹ�c�n-�۩&(��,����Q��C�ć�:G7=�k%#��<�W���Y[a��ơ
۶�vc Y}��[��[~�\W�m��Y���4W�}=�s��A�ar�'�G�|��DA��tө��2W葤�}Or��s�r�j�r��k�����0����>��r�v��:KYg�����L��uA"��=�3��F|���.Mi7,�t�tɫjm�N�f�b���qM]����#�Gr2z3�_�,Q�a�f��s��@Gn>���$7��:F@�܍�����l�o���N��|��a���'��ә���Yl���2sZoF�[t��P��Ք�<�c��
e��G|�x�/9`�n��P�a�70��5Z�Q'<wΏ�ns0����ĝ��>ƺy��M��涪~EH���+Ţ��Δ(��ֺ؂I�brLc�oq �\�Q|%��Ʈ�u������j���t�����MWֺ�p�����pCv�r�W�_�6�
�f�-�_`�����"^�z�������R�
o77-�B����[$*Z��';�0�'�%�9����ہS�l��jn���-]x_d���1w�V�]���������(�O���'�v����TH�{\T�9&�J��Ɲ񴼦�¿�/�0��_�ا�;^��C��.V���$w�_����t���`�~?�c�S9P�Ypì����cD���i\rEjZ�x+%�0g^�n۝]�Rfj`��FA�HW{2`c��i���A�A�vU�V�v?J�AZ�g���!(ԯ�y�p�D���MIi�p���}zu�W�ޒ	Ɩm��^��b6؈�GF������X�#����<��蛍݌�C_���u��G�,��~����ma�LjOr���t �=Ix�Z�� yM�p�KN��1 e^ګ�|�,1�g�dK�����z��6��_��Ҟ<��_H�G�V�����C\�������f*�?܍��b�0����/�(�\s�5�O��8pu�ՄF-���M_�J�h*�跟:�Lz��#�C��T��2���,�ء�UB|��5�_-���%���T�L��ڴ�|O��k�]c��ɑ��'&ny�EW�?m�H!O����:7��x�=0�:�������UI sN�3�M��,��oq%ԙ�W��h�T����G�E�-�Z�j�X��G���P"��~0+
��hP_����x��@=�+���������z�噆���<���؆p�����$+�����["�|�
1\�l��1*%dl4J4,�6#62��O�7f8]z�8 �#�	� �����G4ԏA�5������+D�Č^光�'���z�h������'z]hU��b���i��9c(ܭ�Ok�p�7�1�/B�8+�S�=�dK��X��+�J�⛘]�i|��IZuX>���2~��zi�^直S����ʽ����B60�#'ϣ5$�Ҡ��1���_N��E>��hY3��R�g��^��G�`K��ތ��
Q6	�!��?�ң��ٶpQ�vp�����B���Nګ���})͈�l�{��N�atp�۲"�K��}̶HY\){��C�MT��ηK�
�W�����*�
"A?�[��l{��F���Y����ؚ�%uf��݇xn���S"Y'z?l����jy Zm5����2#��P�ˊ������{HS 2�O�L�j2�"?�Y���œ�цd�@A[#*�स�6pb�����\�ֺ�,��)����j[���o��`tO�y=�q�{7�t�Y���=U=mq�����GTJ@�S�jڸ�����#��%��2 �N��������P�F%�}}�	���FQ&�����lC_Edc1)��B���^To;��K{ `6�b;6e�������Z�(w���x\���w;�`t��I�f�ala��`/p�l&>>-�����orD�����?��2r����<�Л�?:���uC1B�_Q�B�2��Ľ'�������RP��T��6
�Lb�Y"��%��m�sAX>Y4'� �>��H 	/�>	P����j���VWM���4������Ι�x�<�%�]��L=�
PB����pw��I�;:����'Э�v§G�&��W��$���"~�SVt�`�+{�%O���G����'&�eT��b��JoI(W\�ۇ�i�!�k��'lG?���W_[�Y8�}sR����X�o.�������b��*���/a_p&y�7i���~S�$�5��W���>{��S�`BI�'.D~~El�͂�j4Q�ǐy N{��T�Z��@�&����ݘ�M9����,ӡ!�)h���8L�&!Wǐ��eC߾�L����q�燖A��[�,�{2S���!_+�L��`��b�x�\�|Sv9s��N����l��2As
WW�	?J:b2]��<%{�ǰ&�����\ٿ��}�;3�l~���!r��GC�Ȼ[�W;8�����LaUb�Pi;a~�L���|l�r��Y`���lٍ3�w` �ŋ�\��r��N2���@ά
v\,F�OL+��li�R���*ʸ~a��
$�`f�Rq'����6=��g�Zy�qOwj�D�ſ���r��E�,�{;j��g7����k1o�6�T��P��y��O$&�����Ipo��2��ox�ZҀ*�Vӟ ����M���J�A����&3,u'	�� =���4��]�Dx g�}�.�[���͋�Z;���"":S�J��0{N,~��Һ�B�g�sd��'��UL%8���~��E���r���81��� Ij�<�����.�1�!���B���U0�r����r6k�3��֢*��O�d������l�Q2�v�ˉ�P�D���B4��n#ꑜ�QK#�Y�RH�/���x�b1u´�w���^�:jB(o�W3g�#20ɕ6�R�Ÿȩ��^�cЗ�o�c�,�|������5�l��{'�@�#�cd�Q����f�oVS:o��"�}/��PE6G��X��m��{k�FXEP��e�qSR�/�+��v0א��M��x��ߦ"��S�k��AԄ�$a��u/f�b;�2�vw�v��X����G+ݍ���Ɓ:-5HN��]�x� �TU6�Q#�H����e9�5ӷ:g�HB�e��f���F��Ԙ<��.bvE��z0�	U��>ge�����*����{@�ף��~��ss�c���EP���,�X�\ɳ__���+���@%��_��]���p�?���U@F�K��k�G"���kN�f�K�I����l���m�&#���q`,�_.����>Q�	/����A�*��/�m���Q�o��/,�W#=���0�Ob8�eX�k��iW�R�"n����$�i��Np��F�?>�`��6���(0�b��c����#k�0i�E�X���j�^�;D��6�Kc����]IC9����w��r� ���~"�k�V���K-�N
U�	¨�?	Ș,T@`GFiV=	Hc@�c_vM�:�a9!:4>�<-���� gE]�Л.���^ԓ`kf
iS�]j���d��00��&�N�	:L�?*h��(j�5_��	�5 9���n>1�=}�M�B�8�s�!ѫ$�k�[�*%���*���&�� ��c�~ŧ�i1z��]4����N$#+b�`e~�Ú�v]�WK'��ɲ�N�.�͂���G��$<Y�1g
c���V
�ԭ;�H뙙�F�I>˒i��5{���߅	p�L����|S(�����`�.=��
�܈A���Y�\���$Z�۴������ތO��s���A�9=8�~��D)Nbhby����B�w:fA�O=ċ>c��B��������W4ͯ����1�������hg�;8���M�1=�n���.���~�����4;�m���Zm�(����;a��Y��O�X���[Ѱ<�V#J�a�P�J�㮋��JfA��c�}S��g߮u�g����Wi��'�+9�=R���i�x�T��F�ӹ�e��8~fW�ҳT��� -��J����2��O`�M�h�[��α���KO$�hԁ�Jc��0��5�w�������ރ�Ɉ�t���v��	�mU�'����c���{�@����%ѫ�jm���"a�%׍�LDA�,��v�K
 M�U4�Q!�\��¦��e@c�ʸ�o���w��͡������/�y^I��b�s3����`5*|�.𙛴����=7���&���l*�����4���� �$����Ƞ�8p��yU-NF �_�,�@P��١Aƶ���(@"��'v5�C��B�����R+�^��eF�M�o:���Œ
�F�g�=�d"#��1�)^L�@��3���������t�,��l��HŒ��5�B�na�?ї$��ser�G���_�~�k-Y��`�0�QQ?{N���n("���$;|��C���u�B9�;� �
�PW�����S�Oaw18�-͏��]|�����k9*J_�J`�T�b�yo �|�F��{55ܼj��K\�|�{�I��6l���
��bX��P��o"�}OY��Z���q�T
<kR|��Bɩ���!�Y
	��z��9��RW���(��X'uVKys���z?�fH��zy�����,�����e�ël�l6�B�����$�g�C+m�[�k=����(�s�����G������wo�*n���g�;878k��
�g��w���o7L,��	�[fF��N<A!n+�OS֪a��rd8���}�8���~-vzwD!����Wc�6N�'�T�;�W�-����9,Mw�Ӵ��Qb;�N;*l@.+Ș|<��oS����Ŵ��h����=X��,HC��SG"c>����K=*rЩH=������[�Έ��;�4�V<� !�!����:6p4�ԨGx�*ж�]����dH,������s[X%��E�q�D4�i�{s�W5����$B�;Gۘ	&��@�LqB��i�DI�;����ۜW��P�4�8�]�[�b��}x��W�k�Ku���S��:x��/q/e>�1��1utC��E��O+l���~�1BM.7Ud�$� ��4j�w�&���p�lÊ3�R����r9EL�P4hiD1U�X3;垺M.�;:
��`?��c���K�4ش�IQ�, 	�|\K��>A�+@5���3���m�SQ$�"ϯ�fC�
��(/(5�睺r�lT���_!��́�=�_�!+i���W�<��9�6%p��-*��ʍ��F4���W^EU����HU���j��'�B4�lpM�����-�����F��[�(e�[VE��:X��9����h�%T[s!�]���9bB#@�Z[G�9\��cEȷ �\RGKԚ����޺�}*��G/���D���أ��1�w9�����_k����
�7�Y��7kP�B���ȽJ�|�$���]ߋ4uuK8z�~D���92)C�u�޺[p�"���1�+����Ά�$�>8TO.�{e3q*.|�����"{�w�����=	CK�"�)�G-�g�j�9 �R�&nF�T�
ʾʡb�Y��܁�A*��`*ǀi���.�t�u|����q��7��/����&6�� S/��N8��}�f���;�I��=a��"�F0��,اX/��HY���쫆1Gq�OCi�� A0���_�������n��	S�����D\<��t,}m�����𺭾�d:X�=
0	��Ś�6�h�Y@`�tYMC���$�"��i�M���/"}�(C���R���bȺ/�;y_��F�k.��7�v�2�oK�4?��zL�6gS,�4�=w�}$�@R�0]�2����OwGF RN��M2t�v$m*�E��y�k����
O��e�?����q&Be�3nf@�GK0�̈́�iG��`cz��؟ ��/rɭ�a��\���������r��"��A���/y1�>�崅&˂7`U4��M�s�s��u���Zڢ���4������q��޿�Q�:R�����`x�A�����c���䯛w/^yh0�z� ��ehd̋��74��$[�IjX�a���S.�t5�>�~
��	ܵN���1����^����̑�ۨ�&����Hc$�NJ�V`G�51���(*˛WA|7J�����=�G�B� ��Y�ѵ�Q�z��h�+f�r&���}��{v��5�>i�:���&���]���%F��Br�ɺ��Òa��'�'t����fs[F;d�HC��U����Xb茥�)z�!}H����;~E�Nz,Ж ���Z�#�_���pA��/�aO$�"UPm;����S�is�t���Mf����̄�3O~��votĢ�G�M�Z3�𻟾 D� �Ԍ�~�h���7EVw+�P�L��X^�Ѳ�����H��0R����{xP����X	9����pMPrC3��[U��׺9��F'!/{T7"�iam����Ź9>^�ϛ�0T�+oC��?t��s��Ō>�14M~+��'Ҝ*���ƀ1���+DU�․�_7Ph2��$@b���������)PGvJzd���ű"���zG�0N'�;�<ک�-��.t�&q�	I];N�J�{����yi%��tT�z���6�w"�O�N��.�����ֲ.W��� s�?)1N�^� v&��Z�Q�ŔwC�f�g07#ּ�)���ڝ����^��~���o���ħ��u�W��kz���g�����:�zt	s9{�t�-F��&m��N	��[�|9����4|M�EA�h�*�;��
�l�m�-+@6sgR�0��W�\p'9i-����s;z[)�����G���_�/�lun���㲽�bq�N�0��q�XQU��i�n�jgݾ��j����[ �j3�F=���O'���Pb=2��>�[�/�w��%�z�LAH|�9B}&�$�,y��p;,I�u��@1��Y�-�q�O_z�V:*��^c=]U�fLc+�\z��/J ��VϢ/��j��Rnۿʑ���_�7��>Cr����φ���GS��4ɖ�`!Ń�3��6���1X�Ӌ�D��A������W{�to���Yz)ʞ{"8����"ZxLO@�U��LS��Q}�8g���>��`�/�m�Yꪾ�*���k��)����7'6�A����tT��;sHc�J՝��%0�Ⱥ��x��^�S���R\<�̻0���>�G������Nv�ʦ,�;�b�b�}(������P�:�b-s�0�l��豁K��f�n!JCn����_��@�mN;�Yj�}���y^�TLf,CZ����+x�큨��*i�P�~�/�F�)���?�������J~�r�Yd�����>�
RfД��a���mq�s����YlDg�?���%�XI�l $�hcK�����������J"oV�oZ�̊���1��pX	 �C%�;?]��g�l�!4�j2%�^�\=F��U�ثq�QF��(Z�rKS��(�Բs����H����ו���:�/_�o�Q� �6�[����f��y��w�z0*���M# �AI�5"W6n������&GW��rp�f��w�c��~�00*�R�b�xI�>Y�����K�YN�7��zސ��>�2/]�3c��_���w��)��	��>Xg�t8��	1U��}��眨��-7�9$F*A"Y���Uߦ65 c5nB|M�稞hh0�w~۳���#:�H�����Z?�U�uLD.H�"�!y�ۘ�K�r�qy�>�c�?��o�а���_��\�1��& ]j��ڜ��=$4�E�?_��)�J��j|��Oc��k��ꇿ�w/��Y����V�iZSyL����V������A6�OL�ꭓ1�=o�\�uQ/��Vﮊc7Tz��ڒ�
�5��Hi��6�A���Q��X|"g6�sׅ�0�=�P$'��+��|�8�W���~.�I��O���Z���۳��(�g�K"��qL��v�ۻ��dV��4���G������1��Y�2*E����I��3Z�J�������#!���R�l(��6D�k�<��d��\�z� ��'[�Bw�����H�����dCP[3�<�,M�D�ǧ1թ��ʅ�Vy�q[�il5:)&�aL$�J�*PM~�j�l��Է�� 7%�����?Պ	��r�ucܣ���a���U�L/�yF�X���.�y��MA1��K^���$���s��=y�<�!�SNyG��5+`:fr�����	�oU+�-\.�\��z��A�|_B�����r�w��<#ƫǌ��Z��lY��?|�b��.,5�!�7�kU��`ɑbk���0k?cD�m�,3����b���E�^�H�`/^����%Nz?�ߜ��T�m�Q�ܫ"q8�o�b.-�D��n)������0�f�!���}2%�zN���G����h�z,rU�N�b�T�� ��<��8�7y-����Bd�+�9�����˾n��X��i�*��̄�
������3?�!�Kv������J�H���>E�,Ϯ�􅽈�=�I�u�'��:�q6�xl-�):�̷ͪ�Tq�?��6C<u5��1*5ԝ�6�@9�8p�6�hy�����'Q�7¢�l��-6q�N]�Oڅ"B-��z	�Z�s���Ƶ+N�ĩ�ĸK�0��M�j�f@"�*� �޲��2�F��rE�%�U����Py�I���s`�߹��[�� t�����΃�ɧA~䍹�S����2��F ��g��ЖJ�M�s#u��(���������r�`<Tɥ��'k��u{!��e�� �Z�g�{,��m�\G�s��,K�D���Ɛ�߀��{�����G�i$@`^��1�ѷ͚�Y���i� �9}P�@�Q�1��	�a��D�1����e�/��1mRޟ%��Tܕ/ ce/k��4HļsՀv��_�lE�eM�M��u~W,��t/��?���9o0���tf��;g/
�,���g3���:,�
{k�3�3�J��;����(3X'$y+��i"�����$+ܻ'�+���dW�A�M�� p��뿻kY/��g$C����尣�� �<gj���U��4���f�Dr�������� >��������đ������.���u��/4
�eh��/��~~{~H��C�q|�W	ϰ�����!D�,�������s�_�X1����!LZM+�]	`P(2ܟzMV�R)q�ZU+�������ɦc����P��,��L�5�f�m�.&K۱[����;}������׳h��X�)��>E}[f$�"Le��T����ɾaR�zQ�Z�!�8�� ��Ğ��V|5��=9}���ztn�;v=�������B!��zP��v+f��I�$���K���{�fx��yD�>;\�n�!�F��������0��p$�*�CV��bVN�/3~L��r�S��5� Io�e�g�Nꣷ�q`������\��nWj��e������H�m.����=R��k�y"��SE֩YD���anhF�㳄Ԟ~�C�q�0�R���*���w�:�3�NƋ�����*A��
�*sN�\�N�-��^�'��GIK-s�S��~kN�V�R����'&����lF�Xirˉ;�54�٤>�mv</�h�䕠s�����΁K�,�8#���-b�"`3��e����-9�<��[��w^Ç��3��|���Vx��`�+	m���BN��/UGzz���U =����D����J�|���x����m�ݏB��a���/}�)����u�7�j�@}�����hv^?�+�'*��Z�ڊ�m���'-�Z0�r��c׆u�;��,7"a4<e� /M�������g�K��Bi@��[��o�
4��l#�+��%k��Zr>�O�T��"ţ��_5do�q'�6a_�"�+�A��>G�R��5��֋3r��*	�Q���b9|eŖ7{�)��pt���Bi� �>�P0 ��������=�ҡ[�<n1�"D�E2?�񖰦�L�Q���XG����B�1xȕ21���'�c��\���-�?S�x��#j�f����ѿQ�`�]��EC�?��OA+Q�٘���.}�4;�����	�<$|���秃��T]f1�%�ǧ��?�7�`��D�\���	x��ؐ�J�,��}ɷ�u_B�N�@���ϧDG�Q�&�P�L��r���f�6�sɈ�ߢPI���b_oz�"J��5�l&������**t��g��a��M�Z�[B�b󒒜�:���m�0�J�1|c4JZ�j>��Z<oIzA��u��o3O6�q�?�����즭L��L\��ٌk��Ps5��}��ߡ�c�|KN�\¯+w���C�z��B�� z�_���񚀧����%?�g�k̓�>7��S�兏V�56�qS���L۴����K9J�;�:�Z�����++�uZ�Jث Y�Yw��X�L+i@��,񃘟����KO1(s�<[�^�IZ�>V���@S|2���ؿ��{��exY�f~�&eұ0X�����~��j=/ͫ-�����G�'���I6�'vl$	��=�߽Pa�SB��(u�6���䆝Ki)s������u�5R_Nj�'{�E��]�B��!�W��Χ%%l)�x�׳a�f��->�B������ƬKSvV��� e{
�7¼A?lH�KJKb��8䶸����߿�4_4�!˝eNr|�|�3n	G�
��R�AC�@<���㌰�Ȫӊ����Ds���a�Ǣ-={��`����H�^���ͱ���_�V�-�GS��E涼h�ޣI<k,Os0	�4�
�7Խ���<�J"�4���˻z�`cA,<l���f�'�am���ّu���=�rQ��n{��ZI�أ�]"o4�~Nb?+�u�
,Bx�N�0zhd���&�]u��"��el�-�^䯱!4���V2n�K���g�d�t�k���ӿ��P��fJ|��\��U��4~o�����tYń��+d��w�R�D����[�)͡]]�n�Oa�Φ����c�g��Qɀ��'=P}|�'i.�Nˆ���(��@�g~t?���7&��h�j���68.�b�N/ݳ�?�aJ����L�KSqJ�~����\<3�#�\����l ����綘㹃�m����O�R�����5!��gVo �q�O �A��X��F�&��Y~��j�Kf�al�`�Dg�a?�_I �u���$����ƻ[�ձJcH����K^�l����^��Bv�<�f}��n�>->�:������Y���7Z��?_���Z�#��~T�b�P��]�%�����4 (���,�)G��x��<��k μ�ǀ#���)��"�&0+��~9 Hg�9����8���x��2��Q�Z|3�m1z�{�R�ّ`�X1���9o5������ñ���#�<�N^n*�W:�.�����ǵO���^|���'H�E`6Yۂk��g
�~���U|����'" �oOTBC(�S���0�Q.^�8�-gM��"����/���kݮ-�q����s�����^�@�7�l-$�����Z#ՙ����W��g�Wa����Q5�Ԝ8#�+
��GP�yL]h��F>0�(R\v��^�ݷ{�D�Ot�8E�dK
zy�x���go��œ(u��EY${y�\�L|/���u������3c�9<N�x�X��Ӿ����O��d;V��%]_��|�u���D����'�,�޵$���3�5�ė�K6�;VYwc_\��ta�'
0�h����(�S2/���=�}����ѾR��ì��d�/'�ЁQY�1���}��%:�&�qs	r����	4�G'���^��`��RX�԰�ܲ�*�䱃N���W�DYGN��(������@���K���~|����O�iɅ �i��i��i��,��;R���Q"޿�w�#��}���;fޫ&�[��lZ���O�'����e�nA~�v�b��/�8�Ǣ�Ðw�CZ����1t�*S�e�jy�_����b�͒�-��O�rA�'�O��Se_�.1��~c7�R��:�70������G.�����W�~��@(�क़���
蚸I��Hp�ѳV���L���ԙ�����J�x�z!}α��͎�s��Zz�1����]��a�Q�d����������P���#]��N��^����^����I$�N{�[��������b��48��TW�yI������'����-�y-� �d��MG���P���X�Nw�.��w# ��f��Ƿ�{������,|ݦ�=Y����-WD�"RC��h$~ꪙ�����58`+�a,�E����I�i+�E�^<��6�E2�ᒑ����|��O�lz���W����(S8scb�3�'V�ڼ���NjtN��'�4ɪ�ܶu�y�}�e-2� I\T�KT�9&2��8P���T }޽�Eem5�B��AS��F�)!G�e[q�I�T�E�kX����mm~X�뢉Mb=s��=1�I�4g߽bz�����t�����.�f�}�
���X��4g2��;G���N����v�U�k8�u�W�zE���O-O�C4Cqv�C��b�C�'H�D,~�v;��� *Iѳ���q�ؘ'�k���93*�P�b��&��W I���t�nG���6�1�<��0�il���&�G0b|��)�u ��Q����������.�T�E���tD{ݼ�$��"�,���^�68oH�ڢH.G�_CC
��`��+{#9r��eސ或o�F�[.��q��V�JXZud��>q����#{�L�T`Fy��+�^�[0�WRF��;E+a��s@�Yc���@_ҽ�f �>Ћ� ڛ����Ԯz�8D3���:�-��3jmR�L���7�S��?3��ؤw�}��iMI��Ii�zǨo�6��/� �x��<����D�7�k6��@A[mT��̆v�[���sR�V���W�BIE�fR2��K�����>O&�{�u�[:��<�`��ŁA}�����1� gՠ �ջt�����7�K�G��%*�SM�~1��P5���[8�d����n �5q�;@L�L�P\ƩZK �I�i�K�8i�;�Lww�H��:��s�������Z'�w�͞f("w�e ����{ ��ؼ:ۮ��\Lh�����MYn�hx�K�u�W��e�8βϓ9�ځ��?u��o���l�Wǌ��:|)`����Ҵ}�:]�]ܸ*�+T��TV�K��e�C��r5�<-�x����e�P�g�x��w�U�w�[�jk��1�����o�XnÚo	M/��E���%x`T��C�o�=�mQ��ʃg�(��RQ�ׇ���^r��L�gU{
R>m���W1`���š�E�.�1'��#-i��sO��oءD�p���_�*_�!�vm�t��k~�Y������{�x���T:;�c���a����c[w�TM8h��r����yY��x�-���G7��G	��53���?�Me�A�j������H��Z8ۣ M�iC�h�ϏƯ���?铏����zX�Q��\�|��*k���8/SS�`zb?c:�}'t!�(�d����Sؙ:�\Z5�-���ۏ4�"W�����5E2���w˳�o���T�u�NQA�P�m@[��Ī�@�yS���t�7�%<>�F�v����[��KZ�[Su�����d����=Ee"^�l�m���c�3X��z����{�:0���BW. �x��$Z
c�#�c\��Υk����Ѩ/�_~�m����_M�/}�߷#wwٕ����$	��+4��D㧪��#�}d��	?l-$�Ukݛ���T����z,��1�ͫsb��N¼�pBgjsT0���-8�1/�\�xǏ���yF�:}V��yIY��´[}�ofOH%�Z��-_�?k��s���À���@쳐��X���L�i�̞#��;�t�!D��[|]��|�)��/�|��/�#s�ķ(0v��ܼ�I�k� ��s�B��8p���q�J�g�븱�H7yo�{���m�{�N�d�����)w�&�<l����3G��q�K��#]'����/���F�#H�S�	|���y;�ퟶ���|f���*ʆ/U��(��H#��Ȣ5@�����նc�������*������&�y@^���Y#	�8|�uьGan2�}��ԍ�z�a%Ѹ4Z�N٭:е��K�}
t>��ٝ���Ǌ�ё-uK ��MQ��}�㴌�}�����=�Uy������܆�[ڵs��ҷ6�"&n?�����J]{w�;�U�|#�Ϡ�?�$�3��FH�b6E=�Z��y���*��5Y`�fD[�CNS5�!�	�ʴ����j�M� �*��$����k��d��� C"�B7wT�6�}=����G�&ո���T���ei� �߻. ����y6�������^E�\��g������]��-��h,�d!	��;�[a���P��ӠV=	2@9�e:(��֞�ԥ���F<lG��<hK�&���tϛ����W]��G$��J���a��z��ETF�|����ҳW�D���r���~���nL�v���r� ���ڣ�<���2�k�m}�Ik�`������z�}/ _��}�5���7�%o���d]�i���E8�&\�d?F�����}0QR������������hXF�1)3��=mo�G{�����}��-,i0���)�P��A��v����}y(Y�
S"���o4d��>���	��T.kpa臢-�
��h���z��i�-��7��ڗ"���|K�7!�ӳ���a�ΧP�j�{�D��7�a	��C�c�bB0DC�������5���Xl=��������p�����n^��>�]�(�U`��l����,X3�����1HM�O��#($>�����$�l�d'��d���^�/��R׬�oGsm`5 k����wmԻ������ϟ_�Ar� _�6-��ύ���&���{����?����>鑏UqJ˒rϽ㒩���nΏ�Go��yv�-��
��|MOϴڔ�N��X�����/l�	}g~s�pe�������- ��K�B��/���Yx�=�Ƃ��z6�ȹD��С�;ۛ9=O��"�+k�c�PSn7-j]陸�S�����(����և��Ҟ�^����w�����tǀ����m��S?w���o�,�^��/���鄲K�m�� )4��1�PQ����EJ�T$%�E%�:����cH	E�N��nZJ@Z@bH�a I���_�����Z,�;�8g�}���2�Bû�b������3+�@v�:J2�Ƭ�0��V A��O�/NXch�N�˻�����m��؛�{<��P)���������
W��O�4Rz'�����Ĳ�*|?aEN,Y�c�r\j=���a#�6���mH�1\��~|&���|�|�LUi�e��PZ�&;�/�~�'#�+2C�}��J%��k�JSA��'[kU����E˥O=�K~�H��nn�ں�7�*3�{k��N�b�[T;�F|&d�ǹJ��_7���ȏ({�X��"X���e�>��m�K�U�J�o��F� [���Q���,�Q��g����s~W�!���>�E.,����S�L$�C� �N�VuQ��6�E���$��W���.J�9���:��	%���N�A�|ؑ�*�٬t~�[�u y�Z�����1�I���Ҕ��')�gy���}CTc����t�	;ѷ�@2:b��er["�2fF}d�8O�
D�	*0艿�s�lR�������&�*�͓ͱ'�*��W(�} �.<�^T[#��1�+�ĩk��)�K#����3l��m��-���]*I�rk��wՍ|>5��5��[����xaTNsu4[r�{~���u��NQ��91�%���Ν̷sm��?N
AI0:aږhV	g-��R�,��G�Z��:�I�D��s�s]����g��O�|Ƴe�9P��(.̥ɽy۠��.I���j,2%��5�;qxLs���*�Fk�rZ���3�2�%t3�h���^��	�֜�D��Y6|�������+�I�|֘v֠��2���^����Zʟ,Q����!�GN
9T��ms�fZ�Zw�=�1��e�YZ%�4M}7jH��~.ϲjL��"D\�Ӑ��ᷚ�b�+��	,اDÄq �idR�޽�rW-d�3�v�������WKSJr,B�d"�??*� ��w��2D�	����bjo��zCY��]��$�C�˓�����OQB-��>;eP�<��%>���]��-#���#��=Z׬F��Ȝ�s�3�3
zS�|A����&� �ٛŅP)���48(	`�cqM���wI�	�1�K��4_�ǜu�m��������v�P��Ѽ��g�n0&�f/������'�1�=7�����̈́�+3�4��	�i%�@y�6����]ňy�m��5�Pj�v�gy�
5�7r����V�G�O����\�쓝m�8����a��nac8\�	��AEw^��'�P9����A4��(�Z.L�T�/�[H�ɖ]Fڲ�D��~�a�����ߦ���!�3���d�`6"�4�X�����j�N��A���9<rr�B�N�Vb��Id!�c9�\<����B�N4P�� �:����w�!�A��U03�G��4
�(&��!�0�9 ����˼�cI&�)pU��\�喾�"ԋ��Ù��������/��X#���O��\������ϲ4wl[t�����Z�8�:����򊍝��d��jźl[�{a:o�Yɓ����/T���[�ᒭ���PV�~WZ�5{:g�핒V<�l��y؎���q��$Yx91��#�����봡36��q�z��a)��P�b��qP7E�O�1��|���ڸ���"�M��zr�J��O0��UV�&	گ����AO���)ٮI:��g9�?��qX;2�| w^oTE���6u�M�\P�f�FjO���N�&^��M|٨ �gs�0��î@�	_���g�^�ݮ�b]��6߷�����̻��Vp\GȘ�Ud������������$�j*A����mϗq\�m:rb��@7���.�ԟ��y��܆�1��Óղ�Z�L�z2�2i#����p��M���J�Y �.�`�OQ�.YjR;�xч�bL���M3ʡ"�n~B�2��R��)��V(�9�:p\m�A�8Ig��l��Đo~��f���T��j^�����*߂��Jl��٪w|×~�r=^4���1��Jj�\%�*`�/Iq�@��o�J������X���>�ri=��Di2���Lݹ�O;8J2��a7��̌鎽F��}�Z�ן����z�����˪��6��!yQW�ѡ^��ά�nK���2�$c�����M5D����7I}��lm��ق4���$s*0L(��z�>�j�C�����uגH�`�#KWZ�R��ړ��,�,f���_�͑�r����wv�a����$Hmuw2���A&O`�gcf}!��AÔ���T��~�X��Z& ��qn^�x����Rk�&\5Ae����!r�`⺂?�i�7��P�$���橲��µ�y�0Ws.N����/̷�O�h���8�%>�o��ç��)dq:K�&|ឺ�n7�ioI���o�E���8�?�P|\~���77|���isvP���Td��l�6<���jX�\!�S�+"�U@pJC��Ug��[�ٓ����۩h�zVY,�Sd&$e�e~��_?N��ۤ����V�g�W���d�>�(8���8��ˤ	�3�N4d&*��p �N��w/��0��[��$�, �k>Zb)��;-oN׎p:��ZvNP�"RwV+����8��q�0Ԛk�K��j�뻣�Q?���e�I�=��oө��0�\$M,�<C��Cp3d�?��t�"�8�a�O����%{��G
�M�[�Q��l����iمX�Y����^VLI)���n��a��x�IL�,�	���km>��>�o]�m�����֞���;����SX$���#�6Ȁ��^���Y�&9G��e%%u����;?	�wmdH<��V�Ot4j�b�
��K�b8I�J0��l��@D�w;�8��ET[�/R"��r�9sr�.�+�7C�uO�FŤ$�6�r+W���M,1��'1�®�UT����#/��/4]���'[��f|������ĜJ5�;�y�W�ae�; p������t{{i��B:��l֖W���*+�#�;��O(:xy�.�W ��2��u����g<��և�f.�6J�-���&����zT���"���ʬ�4�-y�؝U��(x)ى�%����o�=ϟ�.��n�(	�MQ꺶��hTܞj��_��b)�z�|"�ɲ�Ѡl�t�v��|ͧ>ؖ��xp����wLJD۔S`��M��Pf2jTy�>ZI5�5��d<[H�w��3�q�͏P$�Rqm?ܮ"��;�}0���> ���h��z�Bb���/.�����|�3O�3��1�k%H�f�n4��}���I3,v��D�!����DcRև���EI����<U����cˠ	}����QbQ�裍�$4(��8@�>ӣQ�fM�.�#`����a��w-pJ��k�c��A����"]Z_��#Ϫ_��d^[��q�!��r��RyA5�̬�����.!`f�tW����n�Z�� ��݁�N�������?�ղ�,u�MKʼR�m�hQ�՞g����@�����l����͟vs���j�v��_*����v�j��\��f���Z}�a�p�n�S�������x/�l310U������9�J0o�i�[�����c���^.���{��N9���>/rx#�VKP�;A(��u�g������7�P�d�O ���+�`��4��2�� xv��-�؞�Ư�i�x;��m���{ŠYUvi�>�=x�2.g��6�n�n�����6",T���a�����(:�F�q�I:�)ie�d'�����6'��.��u,f�~�<������.�v�������оq��}��Ӫ��0���~S$p�C˥˓܆ER<Zm��2�3�� 'V��W� _��1����f���k,Fv3�o�������a�/j�>���Mx����=�x���HҔK<�p��ݰ����~�����*[�v��|?>��[��U���#w�[p%IBvߕ�t󼺮5=�a�9w�o�L�[ވ�i�\�V]�9��*?7�#���8[�z��7`p�m�x�r �s|[��؇�E�i�D˷2�D@k	l$>����EY�SQ�����)��|I y���f��|�>`,��|wW�0U��׈� $[ˣI����wH֩�vw՞��3�E���^��B���#�;-n'_�Z�KD$�����{����u�u1���r�Yp$)B��˼"D�W�t
+�j�$��'�a�����`����s�$�0��!�P`w�YF�,`��9���U�?��M�p����zT"H\��g���f���\��O���N�2����T6Ӡ�g>���(�G�$|)&$���]��:��8/p���%�W^��b����菟bCwd��L~b�p�q��?e��T�C�e����_x&�"j3q��._��x@��:��)\���f�+��#�BZ�F�g�� ݏ�?�c��44�ug�aNL��=Ӌ�}��r����/h�T�VWV���t�V8�A�n ���X8���k�$�&O�<s1������w�v��F���7�A>��6�]�d��$���)JϬ&���雾��#��jJ�ȑ����� J�w1(� Ȃҹ�r��[JtJ*�ޓ�c��Tа`H���zr�bG������[f��c:�U����%�����4��S�nՌ>�X���y\=��$����Fz+��oo1Mr���0=W�m��)��x�k�&�����H�*�GL(!��EI������6ma�ک|�y�}��,�I��mZ	�Q�,�x�5��e�l�~���0�4c�K}�RB�_Zm}��}�`O�y�rK���%�b�\F=o�L�Z�F��qaޢA���B��()�TƌZٱi2M2qj,��F�
��'f�'����eƼ�S*������� �On/m�w����X��
�*����o�oLj��?��r�H �<�ƒ��>v��,��:h�)M��D��KCb�vM��o+�,I�����D�o%�<�D)�l��2���z�œ��w�I2��ZO��&���l�U��#m��_�H��"){���?�[9L�<��㻎��_����Wz��[�%"߷2 �;���Q�un�$��~�-��Y"�=�� ��r����~}�"�q���V��|��.���>'���ͽ� ����ڛ1��y�#:Cߋ-7YqW�艁M:!w�#�I:�O�Q��s�tޅ�*��Ґ5_�ww�0�D�.rԓb�{�����!s�
ǧ�'m
iz�;`u�)=l��񧶧,�/���UOѼ
�a~����a��1������Y�����C3�(E�Wƙ�r�T����N�˜I��ҟ�H�`ULj���D������GM�z���El�a��F2��Q��6��|��e�Z��N̹0�{f����f�w�O� ��M��s`�<���>�~ Lר�X������w������r�<�Pe�3l7�Ӻ������F��̗�J�r��v�K�[_���m3EZt�%�6Ƹ�Ckw�&�k�����nWL��:.(����,�[�|��lVakQ�]`����`�
O���H	nt��X�C�b15QFȠ$4�p��iK�CJ����Ȓ�������Q�F���W;�*S�Z\�hs��T���LYo��lּ�t��Q�𖍂4Ý���ґͧ��S���r���7V1)R�����{O�8nثv��D�n`�_�)ܳ׃`�l=4.�#Z*�3����s����0F��ܓ=�0�؝����/�v&�}�K)3;�Bq��Ӡ<�+ ��h����;J��$b���˓���[M�N�xtg&s<����j���H�����P��E�ͷW[(	';Y09hcj����@�IP�l�&�g���o�5T�#~�a��崙2o��T���3�޳?�����9A���Y����+f�z�W�5��Rn^?5�ᥚ։��_4��Fj��N�Vڋ{u�����R�H2��n�O\��6EF� ��Tiz>w����11����S��eM˓�-��6��x��ּ�fan��ǀn���#���11�Fa�b�4�����"<\=z'��&�~����a��/,`�>�A�)7L�ڇ�6���b����ɏC�J�͆��4��*u�bӋ�����wQj�GYwa�	$?V�a T1���Y :�r�U�O�0UZ�62 �S3�(���JV��!�d� L@y=���` �%��Ȧ�^e�oL5���UK%b�6Yq�q��\K��֭L{�ԍ�Ls�R�)��W�T��}��˕
�jl�h�m�������ݵ����f�d&� v9���WS�	��|������*��@��?n�{�*���T�Sk�W����4�isT��h�+�0�l���2.`l��H�t��z�5�|�|LBg.�lMs���V�\�j�	���%>c`�
f"/��9W���p�g�� �A�6<���aD̦P�A��u�_�&3�A
�$�F?|�H�NnGn�6�� �7���<�6��:5༠0>��_	�����'�B��C%� hB��5~�r�؛����%�!��eW�_�� b}}cסuFyr�c��,�*]F��m�La��x�����:�;��!�ڗ���p$.�zI�^��a�L̤>KM��������6#�U�K�V����[o��T��rU�EXE�ߑ�Ag=U��<'��z��]�Zm�]�H�>�IN:����t��%�� �p�<4��;Tu9��1�`TzmJ���6��i`��������7���I���;ꉏ���Y/uDCa5F�<�UK�G%��� MZm|�����q�w��ٴ˸�����n��$��3�'' С���!���+��U��<r�T���x��js���j0��<	��0�0�k"�� c�F}�vǉ�倌���-2�����~��w�S���f�Ϋ/�]�������4�\��ff����U+lGc�*�?a�i�k&q���s�9)����4���M�Ta�0� �f�2��B�[��o=1d���jR5dlj���\9���)l@��Ҩ�6$���Z�v�\��v�̀"����Īt�NB�͒�,�vz�>�LоEf��{h�!�&\r��4�|��a�@�� W��BWM�e���e�'�ڄ����c���ϧ����W�١�z]�@/�H��>���ݔ�e��#Ű
,�"�<������w�I�(@<i�#�횐��R�k�m4^�~˫a���w��c�׽s���p����B��e��%�t֟2\�a1y���T��ݩ�ds�M5x��*��G�=��OW���~�HO�S�~���p�z�\��a�Y�����G�Mߠ�0�07��p��E?b���¥9y)�?�E�HɅ�ȁ�����]p�/�o���s��^��c���y%ܲ�r�3�fAQ�|��?Z��R�9��A&�ˮ�i��xn.X��幢Y��A	x��;8V�#��l�3�z �i�&�e�Xr��_y~ф���U"5t����4S��=C��/2:�l�{d:���؞�?4�?ϯ�ez��Q����bcZ�<���T��pS	�hll!�WAr&�c�	��;�_���1�i6S��J{��w|}`��oqD
R�Y�Eq��(e��TR��d_��X憗���#�����6�|^��O���ڞ��		1���������=�����SI<������x!���%e��Oa崯��_1��"�`����zv2�����?����	�zJD>.��2ZM�O��vRHCƽ���"�I�c����\s������
�[�_�ҩ2�t󁍞njg�(�܏O�a��EF��O�MxP��z�}�7�q�����5?�-�R���k����o�)\�V���ly��=~�P�aQ�c���&�<uU�U��f+��l��n��v�9�`!�E�q�Ⱥ�:�8+nBN+3?b'�¿�՗]L:�=��}2��F�|,�rE�ʰ���1�e���i��L,K�<���w�FV������|R���"������/�W�L��LY�K�&�G��,H.��q� |]h�ev�,���2Tȑ�T���C��$��z��H9��Lf�[�!���<�����H͵�l���������:�����ƫ�I�K_��<G2Dr𑋛ȅ]��w�.��/�k���b��иͼ����O�d�Nry���OsT�`��A;Li�U$
�6���o�5��v �8wm�"���q�m�z�M���L��~�o��w#~����>�]�P�ć_˼�M_c=�!\����Z�#=ܞ��h��3�<�ě����f=��b�v�������^����5k��2���0�����ï�$`�� F�3�+N����.pP�E_�Fے����m��\��ao�nN����$u�?_{h���v����+U�(:��C<���E��t�3��`������K<�X|-y:N�j�-G��ɽR�DL:GLv��`�����ΰ��$\Ea�s�p���5z�N�g�������
I)w�oEgJ�"M����k�Xߍz�{)��@ĺ�y�%!��l����i1;�������kB�,j�?k.%��\F7Ń�=�g�PT\�E4��i5q�����{A"�nz �-1EO7.1Et��'L��FP.�"j���[�@^I��S�GsMr�j
;������L��n̳�����ޜ�2s�ޥ�	���a�	�gV����tե���^k�=ޜ�*Ϣ���ld�_zp�b��='*͜F���B!|�i�F���1i�m���1�k�n�c��җa5�o���LI�	�=6^����V;��o]�ٍi"��kӰF��)��Bs8�C�]u�L��9�K���)�yw-�!s`#D����rw������2L�Y����\u �=C�T��ȅΥ�K���2�?iƭ1�H�v2Nr 6���Q��?% P3U��v�+6�dF?`���&��{�ãH���u�8��A(L� �ܚGv��Z����H���?YA̧I�e5%4��s�}��,]���	΍ڈ�w2ة�ša|g#�+5��&�������LJg��8:���n���/�"1�n��*�Ŋa0�lww;��=֤�i?k�a��UK���B�FZnyŎE����E�L��Lӧ���^2E�:�H��R����t��L���"�v�EË���:(��of�YЌ�,�e.:)"��(��n�&�N����t7������n�ǖ�	=G�T1�*pʕ�]�s�jn��@��]���jG�iyu;�gq ��e����n ��T��r�C[�8�؇lb�f�6�tB��j5noY�3�+8���xcuʹ���#^����pn4��M
{w��E_8�4�? ��@ƽ�'��=��d���_����P˕���K��q�&?x�:�I�=��5k[����!�@{�إJ�S�JF��I,�����A�%�o���D����t���P����j`Q�M�Ƹ_��
� #�-@m.a�ED�{U?��Q��m��JB�L=�d9�Z(���
�+:�3e�����Y�M|�W�ޮk�*P�U;����N�Z�׶Eы ���o�HM��ͷ����Ƒ:Ԁ�\7�:=8_�̈́���	�� X�^��Q���_�m�+~��-:���is#)M������0:�J�����T�� ��mSk R�A�/�\�_8g�v=y&��RR��5կ���D��/3'0�/�]Ӷ@���&�`$%O
��ϳ�o�f�
���[R�	��h@B�wɃ{�,�������oH�?�*:T��y9d��糇/�?<7����>�^؉���ZfGg_�t�W����_��!�����Wr'���l�������y�	����!1��:��,e�ю�~w3EHw2�p�ձk�m����'_"�]�� Q�� a&�(@S!���url�Mn�:҆��o�|�X"��u�=g�������u��y�U��>MC���Pq�'�s��	�\���>�ք�:`��ӎ:-i���Ma��z�)���j��>%BA��F�+-��r��4M�=B:�:;ܾNfQ(���BO����DWa��%�	��7: #�8���6;h��!�����;�zF&�ϯ��ܛc8�ѼOp�Z?mh�_���l�J�CE!rU�@�Oc(���Ƕۯb�ޅ9}�뛲R�#Et�>u�&vт��=9�|�Q+��n���-�[\�����E_�Ŕ�g��Wi�d��EV���k�A2��)��L2���#;>��1v��LR��!��N;����<�WW�оi�A��{g4ל���}��K�G�J�T�j."��Cĭ0��L�~�+�E};�Q$چ�nڳۼ� �~�S��sWԛ�v~.�_�L�]}��s���fa�0ػ�U|�
���)�^�A��ea�y��E�6��|�@r�ޘ.��>��fbj}�I�{_��H�>zz�,u?,W^ڇ8���<�;d�gƅ4�6Z[�#�z�V)����]�r�R��5~�le�T�٪A�0W���Y�L��T\D�=;��gyW�̍ޮ�7��2��u�PEI��}=�)�)�`d2�dO��d�j��V��U�����OZƩmȰ��QW?���Ih�ݲ������?��x�*�Oh�,��JEӉEe�����ĕ�&�L����l7�B�|��E��Z8�1��L=�JY�e��cܭ
.a�1.�}D���h��<L�W���ə�@W�U��uyA���i�5T�aN�˃�&�����VG����*w�2b̒��we�-�GÇv�zn�j2�=/�{zWx���5��N�IB�oOf�w�٨�J��	�U���q�Hb�ԃ�!�j�o�.��V����qFv_6"
��?>b���g3~8f u�#F����g��/�=׏=�w# ���i��i��d�l��As������C?��U�:�����~����F�	]��_�\F��y&�Kx2�����3Śi��py-ə��7��Y>�y�1^	yAm��ƹy��EG���Y��Q�/By7b���Zt5��%-��Ӵ��J���[)����y�����������4�M��eJ-耫F6?z������^�v���^�{�L��vm��M���3�ӧG���ʇ��Ȥ�w9$#�*z=�̍���L���o��Fy8��s_V�V6�%��@�=l� �,a���24���������\g6D���y�������ڗ6E�h,�Ψ��&1�}7b.�iOGj��,��PZu;}*����{�<0��=x����!��7��~���Æ�5{n���o��$��ظ��d�vV;�i�M�����hx�n.�i�����5E!zt���D��� �(����"/�n������SNk���ϚvU�bԝ�v>��)B~HC�E�"}%0pYj���Q���a���^}�ٸ����}�|9^��J��׉0��>���;�������Q�n�tCbz�:�[���Wڵ6��,�g�1������i���ʸ��$���n�&�`��:<�^�[�L<O�SY��T��pp>��_�E?l<�����l�?� d�6�.!񓥀�����>H	�������j�7����ǒK�1٪�B?��*�V;}؀]`�|)<�;��3������>~/v�2�+�n�o<c��	p��QVW@��\!aa*�L~#T��4t'¹� ��u�ћnm�yol{��)�#t �dں�F��������7�����r.޷�8���E}�+r+�p���aސ���d
�o%V�[�+s�$�M��#��4��D��������M&�Ha�S`cS�>�_ 
�IK���N���>�$��}�mwQ{��u^��	<��Z��&<�os*74zq�N=��pՠo������9��7����5ɖ���ڳapحH.��|���?=�����v9J ��U�{cV�\�^�4�cC�����ݪ�}+�/���1��I���m����@���Ta�(�`6xb�q� ��)����̄z�/���=	��G��j�`³."��&~����"���J7��߀5Y����8���Xy�A˱��A����N\
xӝDn�dbXT��m�V:3Us�7$�TQ5B��x��<�o�Tb���G��a[�n`�|-����|����V��r���Yu��|�9���w�&e�g�[�0p��9�|�s��_Q4�0�T�О`�WU ��P~�&�~#�bcbm,�A���}����ٓf�a��?փ�Ε4Qp�(�Ь㇊���R�ذ�7���c�r��R�d|a+,�iÚ�����h�l#�¥@��|�@lm��\��Ll'��?"ur�;��E
'��x��X��C�鿡[��ו�ƾ
�a6���z�� Bł[[cb�h0�;�+8�<4�_���1[V#�HW�����\�awf�o;��re[����/�J�lՋB��ҵ\	w{5��E���f��4M�X�c�o�\��'iH'M��p1����@��W(Ŭ.�V�b���Q`([��/�jx�y�嗹�SC���b�=K8���f�ьN��R4
�`���U��NBρv�P�m�z;zUȶ����숏�z>T�=9���8�¼T�2���?��n�'L����Cu��<j����R�l�c����F: 0Ա�F��̍�l M�S��L�7R�Շ1S_��ex��<a����A���GBV�{�����<��ĕ6B�K��-��R��3)�ŷ�۟��,Ƀ�J`.��\#�kz��j���eN|��
έ	yS>�����Κ-�3���gh5��)�9qʛ���������ˑ'`�X�����&MbeMZ�z ���\����lh{�s��MF�*+G7�7������D@���2�g20w�Xod��)�h��b~�Ø�B�Y*�-��2Iڡu��;���Vt���Y�(��@�L�f�����ZpNr��Ç���V�Ig]�jV,��c��~��ޟH=��������U�^4PD�&��d�s�e�o/��3hX����%�ދ}x �bht7J�F��*oɅ��T?���G�K�"ҋb,�R�$j�E����Л�!��Ոi�=�M���YV�ڋ��>�s�W����h�悄��E+6xQ!��}��L�����E�kg�r�;��kE -� W�Dw=a��N��Q��c�!V���Ӓ2�|�la%MF14�0lz�Ј�6�YG���'�H����l�0XHr�m�S�Mj�!��^~��MFf�39���ظ<����g��I�("�A���s�&x�D~t�&	�O IE�������R��b|6J}��Z�V�f�۽Ql܅���/�C�m'�FP��e:et,����V�a\�-
H�rp�A`Q�m�d����(��XD�o$Od5O0U�,���k}Ƀs���sko��99���� ���y�Ǘy���[�ϭ_�zӘ�FC|���c���r��gMl�N�]Pq�RF4��o/�꙱�:
���(pg'�2�BH��x�Ɠ�4���V�n���9h�T4ʉ��w���׎k��!t/�S8�M#����}qAseR�=]�7Ɩ��H#hJ}�i�#;Rk�h�7WB���`Pu�G�J�E|[&���v���ڼ���뫑CIc2�[ZZ������%�����-�r#]�!/���X��j��,Gy��� ���+���	�o`AK|^'�:���g�ﻎՄ��J .v �\��s{�_�����6<#B��8���_�̶jt��E��].�z�Gb��s��凴T!���)�B?�n��H~ֽ�� =�p�B�b�BK��\��%�;��֯ ���Ϧ�B_����_E@mcyJ�fj?"�F1��A�A4��V-�X)�w2���Z]��J&���8�B��X&��z���4H��Sb�&>W'9��+��b
�Y/1��nzsv��ȿ)/�f��Ü��ߥ�ʛ� b	A$�RN�����ۏ��9+5��ԁzj�P��8�Y�LJǠ�)��<�J~<lK�Q6@q	]ua��v�u
����z���>oO��]�?wg����
B�I���b�©1�7�b���f~&O.}��*c(�$ާ!ĩ8i "m7T��K� ��q���Bct��R���D����dJ�p>������;���R�̕_b΅A����y?P,*�O��+��^cË�i(%�m��i�v��H]�Ѵ�"H_7��$Jй;���X�|�Q(������@��Cnk�j�s��L�9O�����3�SG�h�VV�q�E~���T�D��$�B�'��[ �T��G�GWIx�T[$Ƃ��wK�R)~����=~B�A�
��ۨ�����]MS�m̱J��[�ß������s�}aX�vt��F��>�	QS���,���u��g��[�ߝ&od���f��~�W$�L=b(6;
�R�hfQ��ג�b��VvŔ��r��
���Y+�|m��=l�B����e��w��cğ���ɨ��|��Z'�����+���P���Qj jb���+��@�Gu%���7����?�x���l�#���xzC�𣍕W�/G� �;rd8pn����c�����䋩�j�Uy��K&v��������o{�:�{�<�hq���Q,�;��\A����X۟��_M�,�J�����?sVTN��Qd��\���#�%,����db0�T̟>Z�JlH֕�X�&�Ҡ�BE�%��?��	��f��>@-�N�I
��[IFlp���kh�X�f����ۆA�����#d����8���H�T���gEy����c-D�����	w�T�"�agc�`�<�0��j��h�5���<��ˏϜ�kF�ۡe���p,�e�G����I+�yl�k�柑 �����g�����/�s�}��T#��.��GE�O��`��į��e�F��1�֌p"��Nl���7��Dx�w�j+��`��Q覐�l�X]�'�Go(�+o�<����%x�h?���<�YՠMZN�9Š�9�;ܷ8�)�WE�9\��pAu�P|�l���?z�yu��FP���n��ׁ��;XK��OZ��ip�����s��f0��:a����$���{(G��}�u|$�˿҃����{������#h�6֛`-��u�N>~�[Tv���A�t�l%�������E٨rB��ZS�������g�1p��Σ��T����訤�9A�G�N��ȎQ� �#�� �<$��}	ƴ�i�پ۽�3M+�w�"�x���l����|~~��e�:J{sG��4R�du�Հ�~��";����)e�2��Q��@�r}�>uǐ����1w����G=�u���&�<gg2W2��q{[�ß���¹���#�mV�?2��c=�3ɽ��O�
�q����b�6\���]{y�124A%8r	��**���t�S����۾���jTmnm���9}���Ӥ�Ҁ�S���T�K�!}�|[w�t 	�BL�����44��S�Ό<p|�~�
��7�ȟ�����r��HO�E��y7oq�ȳ�N��%�[4*�`ᣳ�he���Akߥg�����`�H^~���<�ʳ�/�f
h����d9����\�3AA ��ڔ P�x`p	��7�9[KNy1厓�<zsp��la��'M�od�>PQE��p��Go/}3Zug��<LOP��zBˣ.�����t؟4k��_�l�4�5
�j�fo�l�
��X�A+b����g_욺�|��ۓҨ�������!�8x�3C+���]�ჽ��U�'L���!���v�ѥL#�_hn �-����xk	.���ʒ�ң�?�w�]^�j�k��.��8����n���i\�_U�P/s��GQN�d@��A�ord��bx ���7a�����+�k�{$��V������K��?�*��2��`W�w*�F�'��Ծ��Y�ϰ,�A}��Y�*���ᾭ��`#��2��eT4s?��(�)K�&#�ͯoo�-5R{m�髥�8���7�8n�F�$�Z�ܪ�T��K	mu�T����]���mk�#��\[6��?#$�ّ���JTm�#�ԄQ�����R�P�:fhG��wR+�|E��a��.�;�:�>�\�����X{	`��b���y��-��d"\H��O0�M@E����!^��z�{s�4�)���ֈ���SNX�u����,:��5�-�� �r���)��6�������J_�1P�}��4�*�zb�@��y>�@1g0^�͛��xh`F\��#���Ja��U�����,Ln�eaiкO���x#qA���ٿP�Ck�8<��5�3��|���j������C���Qn�5��K��u�W���z��~$��fT�.x4~�ߘIF
#� �:�GexF����T�����:_�=�,z�"!oA��U��#�i+?H��X�B���������UA��1	zR�!���.����z�o�z��K]]�bB6�#4o��w��B�W�<���x�'E4Ъ4��y|�1�y�����k����1�b����t���L��)jN��s�|`�}%`�������/�u��X�2��P��TBe�JM�L��'��}�x��TRK��%GY�[�ě�o�09}6c��u�NשG�X̻3�Ul��eV���T���!�����\>�c��d�hZc�6��O���CZF`9T,ɉ>p�S��7G�J�}����R.�j�Y�$��糰U�ކ����L�XY.��0�� Ы�l4����������|G�'���5��ۗ}e��c� 
��;�m�d�n-��` �mK���p?�:����nj�d��5<́��yOv���������-�jn�� �*������;����/WQ��RU��ޫ��H�A�Nh�G�T zE�4i��"B@z/	E��w���~���y2�̞��^{�I(��O=���yixУvk���QXP�ԸWf�?}Lz�b�s�ս�㞾��ob& `�_<��B�j<x���	"{�9�ny�à�s�~JrjM�Ζ���V���+7���\&�/q���D9������mؘ]%$��r~#T?tM@������jN;π��׾��{.?�P�(��դ�#��[W��gd1����㒼0���	���)��T<}_4#���!WB��X��LC�&����O��N*tCh�n7Z:[]\#�y�O��p}�����Re85N�B��ܗ͵�e�,��6�4�I�;���?��.VKq�ݻ��$T,gdD5b�od#?�r��w���V}o�A�Kg%�6����n��O;��3��L���G�H}��~�4�����̉����`o���&h�+"lw<W�߬T�U�#�$���t�� �m5��n�&��rLk(_'�n��{�#>B�'��~CM�����t�5�gX4�OuUҋ�<��y�ڱ:8z�ߜ�4��j�Է�w2[JR����D����<��
���c`�Ľ��ϣ���t�|��	��5�4���BP��w4���{v�'9����s����5Y,��Ui�H��(���v4��p��FC�Ê<����ľ����ܦ����'*�]8?�sEf�x	�_Qmm�Ѕ)�x�f�)H�oz	���9Y�(*�R&* &_����c-�]}��L�x=�|s�x�%͒�I�eIK�=bP�����o�kz���kDWsZY�����"Z�p|׃)�^`�*�a��x�!P0z�n�;�����te�ZW9	����Ҹ)��!���(���ë���u	"�<�Gv�+��si�-�V7���t����cE�w�I�@^c�!�D���Yrb��zkZ��o�W/d�}��k=%��U��dpV��T�M�L��(��pd
���:�� �$��� �b�@'u��__/�L[���� ��D��2���`�����?���)��~0rm��P8d�)h^�Ͷ$�ڎ�o���&2�ٵ<2N�i���,���AF+G�a��gU����S�-m���x���2|\�j;�y�G~a�r�,�G��$<c_���cCC�*���	F��,����e����(;|f������z�h[03��K����k����Fo��L4��2�Wv�Z�����6?�/벷�AE��u���RA�o(m��S��\�%{sT�p%�mH�$����{��X^:[�(r4r�������7S(=�$G�@����������ƥM,�<rbxIG~rv�#=k��+�"���D|2y��X��t��%��4�,b�csEFs���jC������3Q`���Y�Ӊ��3�	������hl$���I��\�PVШ���!�/W��`���O���ݣ����O�7v�t:���D\�dq���t�$�~F����vF�9�c�~��?��l�h�Ŝ�O�t�sR��>�9��as�5,���%zbP|�i���Y1���]�viL��zmV��\�Έ����]ۺ^�Y�@u�lv�q?*8!u��s>�9X	�^+<X(y��I���<0Wr�Q(��Ö�mV�����M,b��c��(�}����ũ�%�k�lv���%!�D?U�4΅Y���r�����5�$������7���U�?g�X�df����;�m;�|}�dz.JA/����B ���9�f��M�O\FJ�w]��L{~+��U�[�
8��h��
c3���\�ޕٱt,T�f��Q{�+�_��DMρ�%����ܬ�x3�]��?�=pV]XX�zT���TF]��$Rj�G���1��[�ͤ)��`�{s�c��_��3�k�����RX����w���]��[`����h"H`�+�����V�u'��բ���A{C���P�!%��9o{Ô�f���>~�5�}"x%�����*�����6s��|�>���^ۤ`!^{e��q����X�������w���F
��]��=���s ǜgD�]p�\�{JfN�`�ڣ�v�B��SVȈ�5��{�{'n{�7e�0^a������ �9>���AG�8�������Щ��:��F�Zp�j��Z�ǵƒ��K�g8��U�Eڰ��P�Z��KF^y�|�w璜�v��nE����))0��L*F)f�
\D���ϭ7ז�������?]Y�jG��]OuY}LL軣7�Q���qM[��|�*���1#y�s�l��of�������/��xs��t�6�}?�4@��]��tDsA�Z����e��I��`W�e${�n׬��pG��5�шKz�?}W�]��9�~u 
}���,:�X&g�JhD�����j�iQT�u������4���V�&e�פ�<�|��=��xV���x��n{��k�z�<:Y
��>��vq"����ߊn9��=�x�xg,�bʍ�ԾKs��@	+�Eb!Z�H �|�� �Sa&j�.�)6��k����s�v�QF�I����c[2Qm���%���.�x���L�Z�������`�Wy�N_sY���K>:�;����;{8o�c�gB�V�`���Mn�/��>�.d����	��i�춇w��0I�(�8�'zi�(LDS�\�t���n��
q�L�x�f[V�r oMoD-f���$�N��wCE��_�=���c���גA��~��"C{�ֶ��x��n�;
�8ݖ�e��е��X��i��P䝋`�gqz�ۗ@ܱy3���+����b���G\	E?j3M��/��ؒ�X�N���M��$H&sj�)��CI������:��J�E�U;KW?}��"N�K<��#DM�9t\�Q6k���yEy�Pѕ����?r�M��t��Di
v\��ʘ:R<vM�Ρ������>>u7����o�%������
3L��������~�����1��m&13��w�s��mI!I�nMD9�a�q'q���Ω�ß�fឤ�p���u�'lTJ�ns� ��/w�9��*�%;��G�NUR��J僎���\�86���jSK�N"�S����Sow��N��2'<����mL g�z����`9�R�]6�w_���������uFF��8�M����������bɴ��i'C����D�ݺ�T��؃oa:��oVE�|
�jiy�����Xj���]� L�6n�&e��5��?J���W��2�\Jn��	�3@c�6M��X<�hz������T�;�R����Y�P�G��j��z^T�⃟�+Wr=������P���Fr�Ȧ�� �
n�st�<?�?v��"��p���R�F��#eV��	mDW�˳Fl5&�
�t��wY����63Ұ�4l�{Q���:,����,�ꘈ[h��O`9p^i���詷�w�Q���;/kW9����?�o��o�-?���Z��YK9
���w�4�%k���ޅ�b쏵-����8�T�}���ؠs*Ǟ��pk`�`c�Bi�Z�(�Q�M�k��|��ڽ�!�ֽhU�� ��G���e�u��F[��sO�����)�O(a?5��"ʑ3,��J�+�����Y�(݉�e��q���3�y����3�Md�	+6��������$`ˋ�����
��_��X�>�T�,�/3��+0���/ �5j�QKK��77 ^�ċ!����d�ib��������>\U�U����z��~~L�q!�$���bX����ȫb|�W.Y��K��l�V�F� � ,��U#h�iN�+�b�I~�8LւX�=��s1�c�Ε�x3P�8��.�����p�ی������ �5�;M��
�*2��LWW��d�9?Ǯ���>hY��2�E�N�H�q~d����y�y�k�K�gE����#b� M��6Y�	��HhsXJ^bwI-*�y�T����G79�� �{� 5y�в�#�-�d�0��c��ݳq��5Z���>I��E�I��Rp1�d�k��?�[�]D9'��$��=P4�E��K�۷�w�����r12�w{��E���r���J&cQ+#'hnȤu�(�[�jS���哓��Io�2,�%��SfK�'�86نĄ�= �9J�a"���>_;�v!��P���K
��O�|a�;��9��l���T����|�%�L8�C��ޤ��1<�"DgسD�T'�$�W��B��z���1���F�����ҎPx�4��/����'!���-r��-�����&���	� 4_<{�*0����ݥ�
�Z��(�|Vj �t�����Z,s�l�1��¡
e�Z���gM<��ߟ��$>b� �8(*�˓_�mHUq�ځ�J2����5��u���T��ng1�Ax�j33����fف�~R�l�x�<70!��z'�5U�ͧY!�T(�T-o���I:i��Q.��g%j/^=��
��K�)��r-6l�B���GU�ϸ85������*���:)Ѹ1`w�6$�Ѻ~���x�Z[?��ʈ���y �����k��s��UG�~��f����F0�a��s7��*8�#\I4��[V'�W�B���BP��qFK���46ӳ��ӗI��v9@�F��Q�K�o��W���&O���B
v6 <�eQ�����~��0_�7�d~�9���]�Ĵ�U�Ѧ��w��}K�������k��2)�^��.!Nz2*	���*&�rl��!�)؟`��B{�#�}PG�8�ݔ�z��e���CRc���}q=U�}�9�)�����6�	��w-�:OV���������l|s�	�|)#t</���k'a�K��f�-DeS44
ٙz�3�L{�<�xn�y�-������"�����h'���������t܄�.j�Jh��[o`~Y9n�T*!+�Gd��8B83`l#�`���l�{���a��o؅'u�5�w�>��Z������5�;M�5*Ю�=�L�3Ԃ�������t���+�=���?�F����%�Wn�8QϢ{���s|�A5�FnI;Iҗ!�����Vn�49F/����X�b*Z��|K����~�N�@S��[靟�~���i_؂�G䧖��`�� �Bu������~�^y�mfT㗈3Q�� �����s��>���AH�a�ǫ-�K�i�n����5�Y�tIzq�0���mt/_�S�T���7�W��I�� �X�t���<(1IDԝ�dZn�߅$5�V��S�^m�!V}�3��o4M��~\��k�p�˿-]�����=�r�$��" ���_JW
p�)G@�3�$�AA�ڂ9���BCbO�t����T.t�{�Z��"����z�P�Icz�Px�ai�}8���^A�ᅺ��N���q�E@����z�х
�@�WooYe�$��$�xD�nߴ\���FZ�d���KVYn��-b$���=HS�iS�n����,����|��	��hKi��d���fX��9�ͥ���x�^%��:��!E�M~��������sx] 2pX~3}��-'8L᝻$U�RuUOuU�9�i�S�ɾ;W��Ia���c�U}˝o�#��]#g��N�W�Xg�ˊhVMv��$R-�]	9w�������] P�^�ɖ��v�9�*͛%���x�砻|d5�k	��v�����ߥ(��3�<:��r�|��_yyS��/�KA"�O����6������f9�fR��n�$ͯb1j\��@��g"sQ�Y�j:Z�Z
a�Ӡ[r����hf�8�6�"�a��|7��K��c�o{�d���s���g۶|N�	�^$PJ�%k-l�NB�� �a�EY÷�1���+a����+ulGɻ���n�}H:���� �I�A�0���W�-4� w�T(qx	T�~cI�Z��j��UCvu|�1�p��셝	Jdꫲ%�4Y��l�}���U��F٤-��|k����ę|�k^9��Qվ��=�g����caX���];��L�:�0��07
<n!�W�Rr{��Oԛ�
�9����J*���N����
��hD��y
��a���qӠ�B�h���N�����؀�����.�"�f����(�~%�FN-*�����������oMB��UH�q/]�?U�n^S���CU:ۇ�V�;��=B�dUXEf��T�"EZg'�nz�N/1��p��0�U�E\�tS��x�����%j����=�W�ɡ���]��)��iܭ�f��d2��8i�Os��D�E�a6�}���u�U2��BS����n&N�6���[�=o��*v�,?:ό��;s�[�2`�F4��l����A��h�t���9r�bS�p�&^s��U�2/��ԌЄ���_R&G�����K����S�xʉ���>�Z�)P]'h����kP��� R�/�BNY�N�W���'-K�M�hb�����h�/i���+�Ԍ?x�� �2�2)��"Z��>���a:���Vj�����&��oSh;W[.���Δ�v�y���.r�͓�sZ��޷W�»�{^�p	r~r�:7�M���.鏱����J2G���Qg<�k��X�fNXv�KJ� N&��y>|5��
t,d� �<s��"��:�Srx�<��t}>5YBB�4X�5Ys����]��C)X���B�;. ���,mǕf�l���"� ��\`&z_]m~�I�P�s�	�f\�P�t��z
����E���xnWH���d��#�����e��*1!o���u+�}"��U/cB�ɣ,2�B��>���5�a��}39�����X�f���ܨ�(��w�OI��3�����Gd�Y���~��!�F���*����BĽ�_ߝ�8��3������G��O�?�F��f��y�6$ ��qvh
�f.��e�B��tab�܂f�UP���ha�g��!q�/���Rw[�@e�w����a}z��q��I7��r���)�DG��f��f��VAWC9>����\�	�죇��g�1᳁�y�[>����:;�E\��u�V���EX�D*�i�"7F�w�y���#��Lvh�銽��NI�z��)ߝxu�]��F��U&U�mcZ/����J�_R"�F��Di��u�*��������˂���9:{�u�~��R��t����=���Ȫ0�{���",�!k��'�܁��4:6[�7�6S���2��'hm��3�^������ޱ�Go�Aċ/ƞ�c��9�`9�*a�y�L��6F?� <�[£�N^�LW`�[l��i��V���\������}S�����%O2%�J��Da��}��OX��^�a",�Gr�Y����.�%�	ǈ#݀�q�?��lNZtYlRH(�oa��Q��&��D)Q4�Ќjggpj=ŋ��w�T���ٙ�Ĕ�}������\�e�v�g���L����"غ�HFV-o�P�e�8=,��}������8���ҋ�ޛ8%t�ړ��.�~�����v������=�_�)����^��f2F��/O	��ge��V����t�%�v�F�I�8��EJ翪eD�$E��Qε������F�^�!�W��bXH�n�?ɹۛ|PФ|�N3S'�1�:^mB�]��D������Kw��+�_R����U9�f�(��џ-�u��K��BC��i�'���������e���59+M?�LxS�
I��%�ُ	����H��ݵ���	��R�K�i�@~r4�Ƈ �ۊu�����^V���'ޢe�>��������P|�B>ȟ8��x���y��ni�{�,��	Y�:ʢ���H�kFr�VG�Z�\}�4ת52�$������9��E�MM;Q���#��>Q:��\4��Cq4��ɗ|���\��,�m�3@�g���La����7�{��h�l��Ğ��M�(l��/�(/Z:-�k� S�MFLsz�_��"n�+�~��iA�H��^�!
X
V��h�%KI)�(����{m��3䝧Z����C���M뜄���(2P_H�������$�x�L������1��!�5;9��&
吨o<X�:J��Z��� ���:"_��Tvv�9g	��I��>�ٝ/���B��g^s{�k�^J���	�c�鞛�q�d10��L��
�>)?)}y�4���l7���97���4���O��"��jt���p9J$�yS�YW�,Z��E)�v��ZD�����4>���s8i&Gj�UЂQ��i���7��v<��D��
9��YU�U¹8��C;�V���.�l��x��9I�N�5���x��L���a�K[	�g���ӵ-[�\�؉^e&r�7�:��dj�>�$�k�9��u��P[�*���L�w��	�w6��}�֟. ro*���F�;R����틆�~�tf�)��Is�����Xs�9���� j�mZb���}��}��́F�%��E�7�AZ^��_�w�@�P~Yc�c��"��x-�W�L��⟃���P\Oy��QcN�1_�1Ꭻ�!_ɐ�e\Pȍ���Y�������J�L�eB>d��З�Y��<'���Q��R�E���RCx�ʘ^��φ;���믦6�g��4Nպw������e���೸��|pP�8M^���4B����?�/P�A|�Z����4{_�JᎽ��U9�:(���Zv���(�o�<(���h"p; ��	pԯ����Q�B��7�gLx/�l�Q�Q�9_+A�?��}C�8��/��XwśR�"��� ���a��Ϛc.J9�>/����Q(�"���!&}wAv����;$��m��YA���1;�����6��p�='e��	D�.S�x2�e�1�滣r�sLô7��[2�e��~ma0��m':# ��t7�r���%�n|�g%�ӛ�+RͼAР@��UϚ�ǌ���T_K����ltL��|�,��<���<�#���/TS�1R�Wf����k�E�\�P=�9٨�;K��^��hp���������a'EЈ�A��;0���ef�M�}��b����$�i��u����yf7{dܿa���R�_MIZQ���^�k�Q��,@����oXk���۝Z>��W�y|�qz'-����QE@�`8@�"w��X��D*h�s1�^}�aL�'�#�<m�o���&�-�F�.�&e��8^�B�T=g�;8��F�=ޔA;�S��,B$)�u�}�%�g'WN���M��ٗt�ܡ���D�M֟���V��j�׵�&owyb�V\&Xu�T������iGe����cɅPXO���f�^�	��M�YZms���2�-R^Ұ@��F't?��X������mۑ}ό-`$)@I����ԝS���M��7��ޛ$�(fm� ��u���=�y�8�} #]@r�%���`x�`%PeNV/�'O ���sOƴn-y��\�I�r��P�i~�aW̲Ȉ���L*W�ќ}�ʬ������FԸ�C�Kɮ��8'kMc�3�/��XWg"�j�r^��5c��q�gX��qU-7� ���"T��,|����*�^��Sy@���k�'�u<q����)l�>�q1�&Q�������b=����>��I�,b8����|�fx�\��ɽ�gO�<�
C�N���ǽ^G1���צ�OP;Hl�A�ǥv����ƻ�h5�h��E�2���
ϸ�Ҟ��f�v���) �x�ʹ]��wx�P)7��:r�5֋�����j��pz2�2�\RN��v4n�%{��>��>n��O�j�͜W�5ڽ�Y�n�M��������	%��h�T٬���E�sŮ�p�"�r0�[�u�7kɻ�r>���wCT+Ww�;S�[��D�zX���	;�����s8浹ö�ɠ_�˳������O	��w��.�~��s��2�9���H����x!z�)6�l4HY�I�#�7�PK   �EX���ɀ  �Z /   images/ba250f07-c285-4988-88a0-9b0d9a82567a.png�XSٺ7�gP(m�QD���fDq@AA��"�tz�x�A)*Mň�4�ޢ�(H��� !�P÷Vt��ʹ����w�93��~ݒ���z�������E]���A�����G�-}r`~�V����b|���/���+h��0��w箠D�-��V}���p��owo���=�F����9��l<�ݽ�T ��/�?]�K���w�Bx�T��Z6�:�~���}h���;7��jwV����c��~x�NR��b���SߴU"q��i�l������%9r�l�C��{����W|g��T�N���eX;�	8�9��K�hd�����t:59c����O���.�źX�b]���}
��#����}���8�)rP a�0��U��E(:S���i�}�$y�MX1c�* ��~%t'l����O�N,��[\�����U$iJj��k_'�Ǡ,3ؿ��SQ/������}ύ�|�B�N뀀��� KmJv�\?�g�-�����ai����ʡV����h��h���bh��3��U��v�!�{�$�#M7�b��d�"���hu)���'�*K>�ؖe�v��f��He"�aKXֱ�������t8ح���ؐ�]�䓧N-�K���"��WH�Lݩ�ڂe����h�X=��l�xWN��fj��sm�{\,fGd�"]]\���9jS��5T��i��Y��h|4V��"�q�C�KZ�{l�/@x|�~a�>�z��1�2��<�a�gk���!
YaKs1-iژ��ҕ�333n�������r�]MMU'�<��P?@���Kجaer^<XND-??n*����ggD�JOO�N�Q�B1�g��`%&F��T$ΥsMc�6�/�<��9�y�xhaa��v�ƪa�@TTtc��J��l�A�0z+0��=�:Sp��/�Ȥ�I0�d�Pt�D�s�����YE/b��yH�ٮl
?��d����RIKx��2IXƗ����v�=<�P!h�>#%n䴫�Õ���[mi�*��]�.�B�R�jS6Ц��ؑ2�9��B&*h�4�,�ԃy⮺2��x`���nm��ay?n��h֨����(��J����:[��2
�BX���) �ād�,��/�}Z�UmT�q��@h��"\wrR��Ä�wf �)QaZ��
3��8s��G��r&"*�8RX=�]3HVdJ`ri�eD�����N����� ��&A�ݩ�H�&Tdp2zpE��|�[e�n6�����[�Sj�"9Tt0��h��!A^���Ʀ�������E�������1QL�CY�a60G7c�S�b�.\�x�K����uz�K���d^�[�qm·3}�Z(d鋣9f}�{$QO�Ƅ���"=<3zZZZ����)e+ �*D|B�P[��^�<���8����-���ź�~���kPPP�l�,`SCO�R/PJ��'"�f�-ޏ����6��h����� B4�$��qz��wʝ@�/@AO%$&iiS:E[� /�ų4kI������#-��R 4jvϧb4!���A�$"�ɘ���^�Uu�Md�*�[�{�5�W)�U����I��1x
%6UA'��
�x'�`�Ӎ2��0�<9�I[�0�����tתZ~B�^ƀ<�x4�\�_,dר���is:�>�&��͔�ᝰ�x��Gc��ݻg��W7���s�h�~钣^PJX�#/�l�ε���xʋ���#�g��"�|���w��Fi�bF>�Đ�,Ƣ�"H���0��� M��&(2g�V��I\-�)�$�1ɖ�V2�9Mr2�c c}�T2��N����	k�.Q�����k��EZ���*���ayC��is��U�dC<� wD6DD��$�H�O�"#?|�x������_��/��m�y�*�rJ�;�>D)������r.577+�N���f�Pz)�況*���wbm�ײ6>q�D���J�f�M�wb%��=߯�$�R�B�/��Oo�U�n��z��tb娥%Q��^��e"��;��^�a�t"�l�_�D^D���jc`iɯ̛k�F��y==��~�#� w���`K�����*�x_N�vb}�S��B �z�����;��3'
�Jg�1V����l�ͧ��&>��lmb���? i�仍��-��t�d?S�<+L2��2^����wv�+���X���Pu8.>�6���J��⯕ �IN=�:@����!H�K��
1���d��s�Ԁbq�&�����J����Z��؇�h��[GGG>�%�p↟���S���o��E��G�����cT�kC��/J��_'78hj���!O�'�����Ƞ���:�
AuXųs����q�
�A�a�dt�����׏�-rG��ۘ�l�������z?Y��\���\��LJJj��:CX����u��eG6�X�O�2ͪt�zuXOt�W�Q�Z��<��]��$ni␎�96~(9�h��sJ)I�b�A��1�}\�G�.'�GJD���d�T�S��״���ol�V`�W�z��^J�rIIWF���ҹƻa�����҂�^���O�VQ���<�1�gE��f��v�+\����Լ
A2��IJ+��O]>��/:�fR�0G<�E�;}��>RZӜ�q�hT?�7���Y��E:_�����;A�0M
B� �̌?�Ehia��Y�N'Ң�>m�ۼ9����ϟ�<'�1趺E�2�����EE���Hv<O*re�!�~�LlZ(����W�)��G���*��n)�&'�Y�tnȒ�:Z�|yWx���,��"��Px��rqw}��g�9Y����'�p^����-�?�����3&V4�(��ŭH]��d��#c~����P�/�k���̦^.ߠ���5�L�	�e���	BN�p���Q:S��XbD�U.i�B���EV��w�[� F�N(��'''�<Am����9�y���Hǎ���q�囇��,����S�S�"�������ɦ�P�T���D[a
�������VJ����E���q߲K9�v��6/,�cu�xWV�Ha�=Db$ʑP�|��O���[<3�Z�����tl�U�c��^Y�����������";{�C"�'�Բa�3��>t����fy�8{�A��#��r�g(�_@"E��5�.^��%�y�'!!(c�eQo���2��𫕾����.˭����j���O�R�Dm���$��vttl]�	D����$Fɣ�6!!��Q�kͩQj+��V��Zx��T����~/,P۱;�l*�1%�J��\B4\�'`�v�X��8M ��2�ǳ���'����MD�fP Er���e722z�K��dGB��Cˠ���3e�҂�U�x0�E��.+mӨ҇a�3Ru��S������swyy����TD������G]}}���U���]y�L�L=	��O�a/���s{jN^d������������{�ҍ�S�&>e�
U�;9��n.��k֤��F�v���E�񥙡���^mrW�C�~
�WP`��=2P!�ؘ����y�ph-�PdL�?�IEE�f��R��p���ϩ}��=k�� ���A��M������|�H� ��1��֤�\�dd)qܝ�E0��ݻ�_���GnB�m !IY��������:tY�Ç[F�d����$48|&���"����j�O8>�v��|��� z�x 7s���OР�o�䑏#�^���		�͈̦aE�V��6�2���qw��W+����6lŶc�uΞ="/R��'�I�vTFF�P�-������x2֖Z�\��M�+�:�X���8@��á�Ik�S�/��'蕪��\�\j&�''��sb@�G�>��|XLt�)�ICڦYF�v�Y�#��B�>�1��_�	sY�CCZD��"���(�ƚ+�8�Fěj$AHR�s�O�Jx�p�Т�h�>~�)���"�������V��tȃ߁"4��h��K���P4J���sG�U�.���k�&i��{yœF����lmllvry�cE��ɍ�+=�����Ĺ4�c�s2羴���֦�鐋

L��%ّ�FŸ}���
������2��d���|nkkCkհ=�ǝ���#�͚�}I��H�C�ꊊ˷["\� ��D��ì���nXt��XT$w�^�T��nbj>��J<*��\�2rˀ,�]��#,?��� V9
d�� �߄o2�2� ��G�-���	ZI��ޙ�^rWC]����K`����J�����4kq7�4"pd
a�iH<8Ԥ����$����$�K��˝B��y��I�?@y�W%0"ڏ"ojaaXȎ�^�r��I#�Ѽ�6�����F;4r�0'�F?���<nQ�. �:�&J;�K:�{lzo���ʁD��\l��$���N�-]�����]�+������T��v��1OG -��b�4��~hQL~�|��U	w6��ύZ��G���@ӞrX�&C`�����d�T�����0!� ��D�`�\��x`����&�nQap(�K TPd�Vq�-��SP�P���K��<
����0����9�I�M���������bC�42��tw��)U�������{�f[�������(���ݺu+���� ��Nx8�N�С��^����9��aaa�o䫹�����~���0��a�/B�����)D(;W��P-��GF:i�WPLL&�c��[S�vEb�S%�	!��#��C�C���̼��V:��̯H{:����7�@[ �?֪-�$�A�O��[��i敿����[	�d��R�ÄZ�p9�ǩ $,���96m�ǥ��p8\�(���K�>��R�xGI�ǎͼ�!�,�;��D��p��������H2���`,\��Ƶ�ֳO�CZ,h%��b����j���Z��NNNPuj�h "��<
��q��{c9a����xΆ� 'Q�0��|��+��ۙ�zR\�ٚLrX���Y8�:��ˤ�ɴ��t��\:�S�������Xp��dL�5x�Gs�r�"�J|�8���t=:�ϟ"�\$/�4����I.6r�Y���y	Զ�d ;33�U�6d��*
F�VD),,�E����d�޲}������"����o�C��d=��aZ���Xz�^�_��j>�h���ɯ ӋTƞO�eG�aM�mѧ�����'��ű��i� �p��Qš\����,��# t���b�g�l�[B$q�֔튎f��8�1��]+3��X
�)�@	�	ڠÄ>�=�(s���3�NS������&o1�Wl|AT�Ժ�{>����`O!�kR�#��i�X4Me}mw�$;O�c@��;�&����@5�uuuՊ�bӞ1�}˂1���6_��O%b��6s����'l�m0�%T".B�P�]�#��́�=�2��j[V��Ƙ�R����J�=�<���+�LMá.���;:�>m������������M���Wj�r��#� ���|�}Po�&s���)�I�+ǫGG_�S����,C�<x@2��,f_*�]Բ���U=;�53g���nx��e����T�R�� �������oBd-���c���Pg<[.?L7�>*V������OHQ��RAd���FB&�Oa����"���LƁ|'�� ؃�b�}6)����M�"�&���a?����ʎ�����}�"�1Pȣ���k����e|!��6|�v����M�)[6��ffee�=����Gcu�"]���xE�����j�&�4(��eN����u��y]�g��Wmk�ik�y>7��	w�ă��2B� �0��'f���D��5[بD�S�O�������
n776��.�b^Y-f>�&W���@&,,>�qUI��,��6?��.�����gkA=5���I4��2{���u"�����gs��B�)�b�@���s(����20�6���V�����@�/��<R$��?�*,4
H��`��Aߣ}د�B�v�5 o�I��K��|�#�G˳��Z)�yW,'�|���BP��`�
�UR�����h;�"�����TS��f���-|x���������D U��n���YA���Q�>6l���0�������N�]��{?�he��B���%�ڠ���� �Y �9����K���(�N>ʈ�69N7	;a�a��֠ٻ�g����Θ>�ø�q�w� ۠��A�U��}�����[f1[:Rj��pW��M�)S����ɷ�R��Ě�mY�<�E>�&s�q���:S��Gr����P�Dߍgp��Ar���C�������@�3�,���N7�DH~7<<.2ر+b! �?��U$í��e�Q����)�}I&�鍽0��̗ɦ�ԫ"�G��ȢRm�Q��"Եʭ������o[GǴ�kֹŭ ��=�,�/[Z^��`�嵠� �1.�V�a]�C��EU�u��q>�L+����)2X�+��S���#��H�}��T_	9� �vy�al��6k �M4���K.�i�����/����w�d@*��l��'���ﻀT����g�:ػ_<]��*��t�_�D���s![�o}O��/e�eZ&~�9*d~4l�Ů|����أ��$�Tc�V�1�_}�l"��577��4�+�4��Ö��$�R��,ӿ�a�4?�M�ޅ⤡�G�N(78䡮k[Գ}�k����.T/���]� �g�RϦ�KW&��r�A�T$]�͆�I}�Vxܨ��ԯ4-{�iW�]���n���?e��2:�M�Wh82o|��<9�8��7=YFK��Z��r�ϙ����33�+���>vDa�0�NXB���f��;��p��K����G��-T$��K��	���~~��[֫�ݵ����9�S�LPe/�����O�ƺ��Jy���/mݼ<~ M�����i3�{�8��O���N<|�P���%��J�>lB^��'�`ݶF�q#0��Hm�_u>����~�P̏��e%�Eˎ��U=���mR��{��*�0�USk.��!�֥�g��ؾ]��T�̱��� �M���@���_������S` @/]�����Q&y_"��9i��S�/�J��khB9��ҍvV��]�o,�<`�ꟙ:�w����t/ڞ�sڄ)�a?���+��uqv��-)��a�.3����ˀ���-l�/Ы���a
.n�(�z��W;��\cl ^�X�Jx�|/�',���0��yv���A�>6Dv�W4֝ug�Yw֝ug�Yw֝ug�Yw֝ug�Yw֝ug�Yw�����UO}I��U$R�lԩ��>f�>����{Q!ʜ����e��� �&ۭ~ؾ+�n�[M���G��Ə�5}�x���_o���{�(=?�}�7W��U������n	|�7�ZB_��~)�A���/����A6o�����=8�p1?`���Sb��E��'p�6���Y�??,��_�D�늎�d��O�thg��K3�W��1���rΊ}ڡ��M_;�t�s��FO��86)hCv#�j�U�f9�Z6�8�S��D����ۜ��U	V���G�^������G�Q��XZx��+��fq�.[��CU/yݕ����� ���󡀌����~A������%���*	�r����΍�&�|�ơ���:�Pχ�ƅ���GYe�����)׉�����5g窎���R��h�V��\g�zOV��c�rG�{ש���Ϙ��R����rp���D��J��inA��B���c����б����?����F�F�� ��n���F5������u�J�އY&�Ȑ	I������S���,S��Y����2>�q�=r��Y�)��C��&�e�/P-��,��Ŋv�"RPv6�O���h)ͱ:xnW�I"�-�ZvFf��y4��x1}S+>QE�҅ں ҡ�L�2}]�*G�*A^�Է~f=[�1��an��h�g(�Ji�����?U�ܪs#Ľ�����膃����Z�]�Ō���_n�����F����R=�1Ztd�9�y�ʳc���x���M��$z�
��񓎐֧��'UD��#��7u����M��y��[����ȡUB����n=�+���Fr)�$���7�4�_W�UP�O����@�e�>�80t՗\d^�0z��M�r�����e�,�ʊ�m����Qc,�(�]77�k�Ւׯ�Jcf#���-�\_��t��o.0��)6������6|B����U�h!��l+�񶄐��k�Y�:��c���o���̲��9	Xy�p��0EB�x��9��]��r�����Cu���.k���Q����ɇ�����fw�j/㸰�����H���OR�n��i笂�Eb���-t*���7�!<��+�mX-�MÝ�zB�C�F�{�&�Ɩ������C��P�,�8JEh��DP�6w���b9ix�>6�Q!2'�]r^��N&H��C�z],��qC�S{�غn�͜1'�W�	��sU�H�uA��>��t���83!Iܚ}�B�~�bB�J�y�S�Bf�=	�����>3��%����^/9�A��_9�`�I󨾥�jU�P��fv�9��	/�ᔅ*�][�����n��S_���!�óX����
����(�	��x-Pp��������t?�/
�K�$[�����-�0�ӯk\$�3}�7��E�K�(Y�50��v�mÛ��̍�0#�4OcA�C�����hQ-!��_��������Ǒ��6|��TC֖Ji�	=����߭>4�@�-��3=)��S�2���*��7�@��\4�U{�vPCX�Z1qRHv�R�T� q$33��G�՚�5��T%��-�+���a�FF���
`<�`f���$]�rr`����o#cc+�dW^N���X��n� $��� 5.T�"��2���a�G��'�r"�����#��6g�.1+�A�r�b0�
*_��!ȹ�U��=�J�z4)|;�:6���mE&�_����+D��YTx+�����fX󺅹�!����Z�5s�A|�(@��p�Ac���Sv��`��[i=�&�o?�ϧ�ʴ���r��v)�uӬ�T7}�\Y����y�h���RjgZ+��+@~��������@��dS�SI��́��;ۀ hg*w =4S�J��3�3g�R�­]�9�A:��br�����s�������c���+��:��Jd�� n��{@��>tf����ò�I�n���a�OUm0�����<8��RZ0-�Jw�ϟ�?��4���8�aذq�-j�Ȇ �7M'j_�RV�4�Qp�SC
D#��!"(mJs�e��JP4��&���u;�*�g�vG�h�^�%Eus� �F�Q�yĴ��L�ta�xz�P(s4���"��P�T�D�Uvve	}�5��n��#_�뢿.��
~��B|u�0�>x�Xh/��1�(�ޫ���i<x���"�̜��*@�]�o�W�7;�)�Nd+?	׼��y�9S�zV�"��
v��@;�=:�&�[�	��AKՏޏ�zM�6�9�廭����e|�2zJp$}��K!���C�:Τ}AG��3p+[�����7q1���B�,�������[2�]�]�K�A���ɍ��C?B����{3;�d6E��y�H�xx�u�B*RmnD��9-���r�\B*K�:n:T��g	��/��&�ڵ��fY���Y�/Z}Q�L�{�� ;��kg�t��k�R�B�hΧ�D ;���ؐ'�J	���͹��7�:z܁��_u�T^�ͽ#�s�|�P�-���T���u��[�9����\BE>}+�<���#��O� �t�N�0D!�Ɔ�XƺIJ�=��������Ρ�ՀX� +b�����W��Be�PT��%gj���	"��zֺ&lb�[ջ�@��.o%�K��>����9jg
����e��.bG�^�Et����\�&�NY�Ԑ;^���
y�YAG�Q�!������ֵ����ߔ��<֯k��B��M�W9p(�L	������߃����>��9U�Z�<�e���s��d6��Jn�S�e�iGHe�3�,~nȍ]���;�um��34�\����p��g߱�.pab[`�����4��'�+�Q#*��!0�*�;���\P<.�v|�d�����e��X��7p%1ǳ�a�m����U��"�A�۹P�Xx��^�v��.\O ^�6��ẖX,�?�©�c�`���1�"`�!��Fw��]�5��窱�^�C?�|��S��4�������^[�7��ߞNn��߷��,��~ ���بD*����)������&\�f�<�甀�`s����Y�?7,���w��W!����?�,�"���Gа�����)���'�����>v������� X ,�2 �i��tt�y��)��	p�< �g��'��`������V9D"]yZ�� �����.�<���2�ߺq����1��l����9�둶kA"����ۯ�|A}�L�~���{�Z�+ӽW���>žu3(��b9�����@�_M�p@ol��v�MNy �>��_@P�v�[Ace>������E�"�C���cٟG�a�&`�1�u��	�ϥ���<�7��ȱ�����/�X ��tMί�f�%���ʃ9f����x��	�yx��9���	M�G��֝���%
~���f�A�����2��m��'�oSAω�}^�7�U��4���OF��`8]���m#�<jXPpJ�;���L����J������������'*��ɘU�ل`U_�U�|vv��qÞ	��ѓ���<���R &u(�.vx4��!��d PM�g�c�P�e����1xԡ��AD�J�_�z���p���e���2?��?��ܠ�r_NkfǢ n�f,4�G�;B�/:��L0�ndl��;�u@ ��ĸ�L��ԅ��X錍��Rݤ�ϢOY��"��0Ɔ?-�.a�
�E/�+H��=�)�ɞ���;+}c��C�L>kE!���h}�������Q��0x�k �-6> ����������<�����qɐ	����'ct�&2�:�#�`B�%Z?ʓ�����$���!Å��Q??:�9�9�F5/��H'����������4=u� ����d�"-=�V��T7�bG �ݠ�)��u��_���f�j!��c��+C`�&G�AV���(�����Z�z�i
�J�c ���H��.��HGG��Б	�>>CV��T)�U��o�}VԊ*g�԰ ���n����+�[��!�7s�-4��׳�)�i��1A|>������>���!�@���m݀a����33����p��2�ܲ�E���`�� a�SVG]�VK�� f�1��B:c"�qӝ����&�x���<I��7c���F
6��)��sr2N������h�6MF2�L�ΐ���xc2Fz��	�Q���yФ�z}�ZS���̅�όG
����b�=��{~�Y>�1�J���t��P-w6���Z��y�``r� ~��l�g��o�nj�w��	�|��X��Ӄ<�w�A�O���ZNg�d���wE�
��/����X&�S�I��EN�Z�f�o�����Dy�n����Q��#���0�w��\�u�F2�������54p��0n�㈫�Lwt�LcR ��ʶ��-EW]�+4��?~Qo.G�l�+2��ΩE`���=��Lt�����w�'+�
w.ԌI���xհ��%��܂���g�\����ꍌ ��}`���^l��`o��q(�����He{{{B�x+s���h��ׯ�H@3��@B�A�P�d^meUQ= ��������X�\�t< �=����:#d4��my���d���*φ�T���_x �?8,t�,��H��2�4`��AFF���jP���mg��j-��gf�����H~�Q$��;9�LHu+_l�r�k��13����ܑğu��h	ٮ萲�������=���!}~!�Q�%(�����L��*�ZQGϋ	~Z��0�����hi#�~mR�UE���*d!c^�;s��Ĕ����	5�
j"�}9�7Yyc.3ջ���=4�Ep+�|o'�P��?3q�gFF�~�bv�t~�h�X�2d�A�]I���H��ۊ�𢁰��h���i�B��.c�;Joe�<Mp�\>�U��'Z��2��3U���\֣�E����uE1l�b�څ�Ќ�@Z�a��� O�L������Y5�������.ΎL�W�8͜�L�_eL���Ѓt�����/8ƻ�'_L��t Tk��W��D�;���s�af��9!R-�喙!�}!����o%N2^��ȹ���.H	I��;f�G�<���C����@,+xX��ć� K���"ݏ$_+�_�7���*�`�S�R�O����\�:�D��y�35�ү���Y Å��}���������I��3���gL�
bw��3n�p$M�SZ�"�6O�0Z�C��'��`����ȨD�I*未�rW*�:g�(oA�aDV�2]���7����
t���x����AQ,s�3��oH�TUQ&�7�%�{��~?�����0��7�S2z�S.c-`ܝ�.�Ʉ�PҬ�M��=+<�_T�����'y�~�ݧ����G��t���R_\W��1�6�3���2P~"�Ĩ��,���\ͥ�������}(�H����/jo�+���UD��]Pvvü�8+�;p�1����r�5���=��m�j�x_ـ���̵,Aj�zNF���V(W�߲YZ(3���9�N5)�r����9�Y�0]��o蕰s�R^6'�=��e�LXA~k��S�2��7O:�b,L�3��-��q/.Tk�͟�u!��]f���ULf�d0�u<�����y�B��=K��[d+��W�s�J~�"W����7��ܧ_��2_"�q�5&fR��u}
���M��ҩc��k)P���k7���?��N���ǲ;�0;_D`���� T�_u ��r������K��E�"`�X,��l4F
�!�&�휌37��zb�K��|���@-7�]��@Q����o �r��`C')��l�?g,  ���w�*tV��̰�Fe,�s�}L�,�X ,  ��`�� ��c�~?����g�R��Ȏl�,+�Ļ�p����D�?�,�?�>�+��,�o_S�`z������`� X ,  ��1LR���X�X ߾�tV8��ڒ�`� �! �+��D���۪k�y���|՟M�����:��� �Q ��~5�~��'�2��Y�?7�o�ަ`� X ,  k��`m1Y , �` U+�n�w۵Z�ܞ�N��p���M���	}4n���usg���w9{����ƈ����������/B������7����C������e� X , ��
�_���x�||�����/����T���YA�v�!yd� X ,  ��`�W �7����Y�7��E0��s%$�r��c�z���>/���ѭ(�gu=d�@� 	���y6�(	�d�'ǫѨ���}�e�G�sr�}�.��p M��m�܅k]�i뎒D�҇��A�o��] ��-kU�&�GB~��a�#�����	��[�ڨ�.#̭��h(� vv�ԏ���GU]~�r�|��w�`��s�/�z�~NW�F�d�}�o�M��[]�H�K����ؽ�߮��<���|C�a������:��?(Yն<ɽ���h��/�)t!��9�2B0%�>d���?�?���1�S��� ��/��4���5]�e�%L�{�,0~��J��V	=ZT�� �F��W��5��%%�/��D��3?yu��B�t�� ]�����M�?.Y��|�s�ptg���:�#����_T�R�m
�f̿�G��Lv��|j��i��_r�e=�
=�[{q+�������~:��a�����9!B�Ȥ���gj��:�_/�%�@�ygƆ�������T�1ier@r���*w�_����߄ m	�����tz�o�ߕ�=u߱2�Ve�����(J�M������:�ٚ[LE�TC�Tٸ9���-��E*x�2<��`�T�ʀ��c4�nX,�l�+�p9��������ز!�s�%�����@�'3���Ū"[u�N�1RP����lBB����r�K����P�w@e�K�����}�+�~�j�^�b����
�8	$o�v��\���ECŴE���8!��Hy�y6ö�(&Q��/�����%��*O/�-���<༩�v�gB�CZO�/�jF��t������A�p�V������ԍS����q�9�@���ў$���}Ce�H|����(:�D�~�3W�D�v5�o�T���7�*�Q�j��jj�W)@�
	��y\�n�F���-���=-R���U�IP[��
&N�k}e+���`���4�ĥn�� �ޑi�����%�ڔ���s������s�b\)���A��˝����Z|�"g���>�H�q���w0"�&1��]�Ǚ-9*ھ>����N��&�b��g�7�{'F��,��:Zx�鲋����$��U���0�����h��p�Kou�v(��-$�V*w����h�kE�U\�Q�ME�hHs�	���2�s�tCX�soNU.aewc�6����j�?���O�a
;�#�s�w'�I��4л9��}<?p��@m�!��4e_@"A�C�R2Uڌ �0g�0Î�./:��)jM�q�%.;Pv�,�^�h~�âK@���[���K��z;��6\��n�+���x��Ɵ�x��s�H1\ P[�i�zR���A�"����8G�S��%;�܂S0JA8j�p��M$�Z�9�� �\�N�t��u���egϟ�$�~�٧ѱp%��Q	�����$�G��&�VP�q�'����^��G�D�ʫ�L��	
ʃ\��5� � '�Gª8�}��o�l\�'Pء>�d3	@�HPK�������⯻��3��䝃�û�� S-�L�%%��$��&�w[_�AE��m�V��_�O�T���`µ��y��Ӣ_�7J�y�Լ_�ݠ��(��R� ��o��!�p�ww�-���fk�.o
�R��V���(H鉢 �h��������J��_������z0P������ɫ���~���� ���ۡw+�yEί�/��FŸ�\RWH�5tV_���3�3�M�_�k3���cr�9�?E%����*��pAraQ��:�b��2#V% ����T*𩎤82���8��+E����[�i��ϝ�J��6RC��V��^��	2���-�n����x��K�f(5��B��AGP����3�څ{�K��Swbr��߉��1���;���Z��I�\+��>~�s�Ҍ���<f�E�/s�V��b�l��̡�c�Рq�E�\,<�+�qf&�w�Ō�fz���@2^�6�k�3d�b�{Ԃ�E5T��U�б�0un�2:Zo���Ѵ�*�e)>"���V!uA���G0�XFW�U�ImW�	�+���L�m�Pa�U^�2'�^��6PQ���� �GX��|�s������<"��w�O
	�&a%ė�A=�c�ݷޥ�y����Iz��AYY�k��ᶃyՍ���+�r?���,ߋ�E����T��#��x�ů����'G
�X�(�z̏�ό�th���P�ε+/��3�ܜ�$�L�O@6�	%9�N��<&�7(cK���#4Z�����(Wq"#HO����P�{�#0� ���m�	�1t�n�v-X������`!�����z�S$-��vR�X�pa&���3���AZkΏ�HeF�K~؎��=����UC���^ieD��ƍ<���� ����K	��xx�ɗ̼��u��?/2����;hE�	K&��A�c��Z���/˹�!������r�^����&�"r�o�j��V���>�w*�g*��k��"K�a<y��el���\9p�|U֋�5?������3:xu�(^�<�W�I�v�yP��o˹v��.s�퓟�^2��u`���#��0�.:��fsl9���m��kA�i)�d�������(��s ����U�nO���=�n�zROM����3J&�Gg���|e�/��]Oe>�E
�-1���&CS;�9�V�2"0�����w�N�5�aa�O�� �2����y��\`M�.��s����8hu���\�a�jr���[�O�N�����X}FK�Pko��ef�_J���lZ���y@���{���咨дw��@��Ǹ=5֝���4/�iG���1$�����������C�@���-����y*@ȑ0�I�F��<@-4�-��0�W;V�?��"�ښ8%��Fg���f,U���� ����
����JOO���aKcc/�t�j5�VZ5l)@��hq�y�a`ьeF��V(��o���Xڝ0NP��Yi�=Cd��k�2��OtW*e������B S������d�����ً��{�q�Ԫ��G��w���Cu-9¢�t���z����Vd��o��Y����A/�0	�ZC�*���Ro�*p��{v�m��?$���"�QZ����<C������VD��&���Ϳ��g������s��P��0۵��]�)����o	�F�o̜f&]l ̩{�Nt'��1�)��Em�{�B�+,�H��dC�|��#è�uχ�x���U��Qv�� ~yQ���;�@ո֦;ʔ`:8;I���*����Pz�4�IT��M���]�B�T���ے�4��>Ú�o�a��1n�^��4��d�]�G��îrۅ!�E�@�0}��i�`k#S+qb ��=�l���`/q�38�ݱWASm��ńV�P���g�/���{� �	�r@r�#�'��-��#)�^~�13�-BOX"	�I��#N �+��"Z5q�l|"G�r���GS1�Ij��d�@��\����
q�L$��Af$iiԕ;�(��熻T[P
÷�I��~X4��	LQ�\�����FA~����/hy���T��	����p>�iE�;/����Z����\��f���7ް`�ɯ�!��a�癅*�I�A��N�D���������<
atX�x��ORz����		�U���wfO��vi��qo��ǉ��gkhq̔s�t�X���1�7OWQ��+bL?S[8Qr؆�q�&�'W`�:^�}��/�TF��8�����'���>s��o�<�2͓�h���v��6j�;�t�P�23�`N���Dc�ت}<� 7�~���)y3A�� �'l�B����{da �|����B��aH��ho���g��(�q3�v�Tw��G}�_b#aWш�3���:����ayb�~���D{scFLad�&f|հ֏���� ����r��dCB�"�E�x�A�K��*a�:0�W���	X�O��-��-ϥ�$��2��w
��#��N_��| N�d���8�	s����	r����2�o��9E����9��Z�b
'��(J8�5Sh����fǞU���?^�����W �<o�ء�"E
��XM�N �$����5P��X%���/wBC�ϳF�A2x��T�N��`�_�Xg�����ʌ��\���Jzŝ<cA�b�j��)f%w��bl� E�Hi�q��n��+se���{�b�/�NK���dٯ�1>$�]�Z�����������g�/|�J0�z���-n��[�-�Sx���蝛���l�WdK�/�D�D�A�P�J���fy�7g�~�12�o���[���h�jn$'|���*�o��l�Pܝ�i���J��g{)��d�E�^[y#;���
��������e ��?nĚ<4}y5�����0���~Zg����`O���_����z�OJ�%i���� T��	�3Y7)�b"Df�������zRu��=�E�n�e{`OV��7%��<�K����6�f,��I�Z��l�9���F
l�9��Fǿ^��ÿ�N=F�����P����r��'4���į����9)EQd)ٓ}	Y��T��HD*��$�2#J��]kiƾ����o���<���:��y�>�羯�}���u��rih�|���hTr���
Pf�9R;��|�|��D2���N�"yQ�����Wb��x�) YsL�+ke~��m�U���G+P�|𧩕��� 6M�>N.W��.�{��P]1h/&_�S@���Lĩ��^�PP�R�$�;��=���>^[��r�yÈ޶H7�M|�eP����ݑ��\,�H Hz����P��IG����S�.7)�P.[�\��7Vb?�ā��,=)�F��@�{Y�SU�u �P���q��v����l��:��G��`Eky�1�<��3B�Lq�O��2��ԃ	iI���b�r���%M���O���"?��U�`0;Aj�MD�k����|�����I��4��=r���Q��0q��wB��m� �C�U?).VS��*�B�JMCfa�X��u�Tb��T�"��P}~CX��Z�G��.�VF-�/[BMD0ﭗN�-�]��Np���v��-��-�o�Ņ �Q0^�s%2�:�tFZI�������˳�?��L�J�9�7Fܞ��b]���n��u�^o�S����}ͦN�b��S!>�Rl�=�P�����9i:Q���;cRݦ�Ey$�\!(0�X
뤦�z�X���R}N٢����'�$� /���z�ˍ :,�_�Ey:�D�����I�3�b����Y�Ŗz��Ȳ�[��%ף��O&#��<}�Z�д�<�Q�%Q�������	7@"�a�����KDa�����f��X�����:� `�#�^��|F8�� ѵ��M�	�D|>}:��NTڰa�Z�m��~�'�;�����%��� �O�	؅�) m�ܥ�y�j�T�o��LIN�"�#�z�.���u��"��a%$��%�1H�$a1�-�����'	��W>�}��[V/�hioo����r|ڀ�E �FuX���N�;)�sw�-���s�2�J
˦MKP���Ѹ	���C�VC�����a��p���dFVV�s���* ��_V�.�P�v���Q����>,��W��nS�fDإfO+�~��Ovb�??���?=N��H���5ky?_.R҂���8qk�V�)�G�����fU �5C:^�5���� �z*�B�b�:� D�Ch*Ya�]M������L��V��:3ľ��� ��A���1�t5�)Ÿ*D�bJj��-U�Mm4ky��}Ĩ`��f`�kC��#��v9x�����p/򉈷^����R	@eAo�cw޹�rz�w������A�au�~'Q���:{ȼ�n^>c�!v��I�G_�*�7�;=�*�*�!��X���7�rY�Z�O+���H ��#�VBRt4�Z�Ă{b��X��2�X�v im�����1B,W�L{s�������}�}�<E������\臝�c��:�8Y�y�0HY!L�|�l�����M(mHT��K?H��]��9{uh�#���1 &Z����z��)���`�aH�6k�C��-�ȷ#�?$`a���;L�}�ܚU��F-SXZ�dFD�ev����:����L܀�_��)���3�I��\�6n�)�Qp���HM�܆Љe��ϳp�ӽ��i�^ީt���-zS+bC�]�5eo_���J���M3�-�l-\�lR������<V�r���>J�6̶'��'tD�Љ��7 6���>��%b,���A X�$(<�EEGc�z?��_��6o!���+O��-�X=E5����M��E��z�w���6��=k��y�ϡ�QF���/��=�=~H�=}�!#�Pe97�����U=pN��4q�H�J�����j �3@1����{t45����
0���}S36�)�W�Cg4�k�.GF�h͋�kU7�c(Q:�r!+r��h�buj��A}��.>�h'��ј0����Beq^/�H9���4-++�o�ĺ�
�&�/��5Hɹ�i����>-(��M�q>�-//�JNnㆉ�g`:N)�S]��y��@���i�Q��T��"�k�_/��8x�MeoZ��IN�=��c��hU3��I��o5�l��o()���%�e\���͒1))�K�M�p��R.wQ��&�vFqh���s�̩��u�;/���F�$j1U�bxpv������D�i��Ql�ֆ��Q (���5��G��:�g,�;?�X�LW(A�Rrr���P~G�I��
�������;4�9y̥�sUS�
�� �W�W�:��0�l��)�h�D,������H�e ���D�_�q�&�y��oM>�GQ;=sE�päp�V$���d��)�2P@���ȶCۢ�M�i����&�VX�<�_����Ah��3>cw�Ea�49}�bnn��dK��=}����6������غ�f@�=a?�0���Xu�TXeʆ�2��f�@֮p/��ܜ��	�dy=P{���:�Gt#M��Z���e���QS�\x{�����S�N��8�d+r_�_e>���
����/�ܧ��C�%��}��ORm�H~
p�<�x��l�h?-����uE�_$U���[	N�5��$$'� �t�la�a��X ��Ca&}b7�
���헕ɒ�Ep���~c͡G�C�4ojm�*��)�ul���(���z�ů۳����n<�ݱ�X����������J�y�G#uLa�g�.=?<�R��)�ͱ{z�QL3�\*�=��G��)&��:�'��r����Z>������y��� t!�B����fP���x�'}�%X�3�;:�����U�;��,j��#�Z.i�H��B|$+��`�6R0v��;H�1V��|�ތ��|t�@9WҚ��Ȭd�N�IN��c �����VU�dMM2��ܮ���BvVc�%�0�`� ?��ˀ���^�{�ײ�Y�N�����X����9�r���@n[����*��bt� ��I麳�ǰ�,�.&�0���/&�6�%ːl@� ����R��pv߈*��� 9�6��|�����Ħȃ�?���A"&:)m :�D�H�ғ�<�	�8�7�ӷy���L�gԁ���N���.�n�!�PA�8׉���������&O�UA���fl9
�?^|z�RJ���O��'R���K/�W�����)EM͖�E��ؓ���bq��<����-҉��,�L��$��/����D+7mڔ>�\���88g�:C.P�P���|�p��P�He��8�ͫ��&�7��õt���l��o���QdA������{������T��pˊ 4���R���bX�1|0t-������?�ߥM�3NW\ N�:��?c��T�s���IpG��w��SCƐ���|V.ѣ�p�O0\a87��r{��<��n�>�t���-mW
ky������o��AFJT��|^�g���0<����+�����C��R�^����mE����:N*N�⒦&����Ђ�}��8Mz�;����Fi���w%��ӪQ����HE��b�������O9�3vuur՝�8X��kr�NWY���0;|�4}��<��|X_.n'��ߊ����J�V�H�bkHJ��P���M7x�)ϗw�ȱwi3�F6��̔	ס��Z��I?�Y(4��3]�����YX��dd�F+�'�[V��V<D�P��̽��?����G���b�Gg���� �b`gZel�q�L�Z�r�F2`��@O1�6J������B�׳(��f�Rí�Ɵ�)��3�882��-�h��q{��[*C�ut���'�B�?����f&~���X�,p��TZl:����H@�T��gƂ�&�St�*��Vu��E�@���k?~Qv���;T�8�>���������l������d���Ҩ�����[�Y#_NUfxNT���F��0�;���*^��}@�b��4���.^~�G����&K� �q�Jy�%EN'��� �hS	i���3ci�����$+my�YVjBOO�QP�0e���uqJv��u��_�\���Ӛ5�����2u
��Y2�;�{�; �l�7�2J ���R�+t�I��oJ�����@ "��t@g������㦋������=}U��,___+�bؓ�>Ѓ��.���kUYC��U�s��MAJ�{#�փ�"��n�%�?5�;���ϡ���H�z.�����Y�#�E �P�R��p箂[�|TDRl4���S�D����>)Ncݿ�^�Q5�r��M�`W��p3@ �A~�_��h$��yIv��=`�8�Ë�d\j���3f䯌�H� ��VH�f^��U04���>����}?�)���cʮ���u�,��G��04*v�m�f���eJl�����"�k	Y��/�j]����{0R>�������^���D�ʗ������X��8<8���k�2����/�����]���ٍOW7�%�%&'?QVB��Y��1g����r���y{�&'�;	( T*�+��V��hk϶_^}!p�O������Ō���u�b�he�-��Ã�6�N�O'f�a�n��>�����ǯqy�ww�eN�銧@G��k'w�ɮ?�@��=p:_k�T�n��j��ȿ`q�../,A@�2��4$��ku�i����f4X��	�q���]a;m(���aO�k#m�4׻w�����v�/� 7Jo'?=�ZFG�O��������ɋsa�&�`s�&z�Ζ�ڸ[�)�\WEO�A8���s{���}�� �G��|��c{�U���s�. u�����'�9O3Ex/�C��6�С�@~���.W1�͛�/�.(�f��,k�^�>r@�X�xQ�@������L��4c�@�?��k��Q�����D�&ŧ*V�]L��[UV"����Ǳ�����m�x��BTЀ�D�h��OWu�M��{�a�T���32"�y�?�Y�J�/��SJw�� z�D�i�Wc�\�鯥m��2`P�f֞��`�M[7�Aw�i50��~	�� _3����T_��Dn����HϠ����,��!h�V�nlt����U�*���8?
�����̻<�����
��{c;D;?_.�@�x���t�D.0����;P~���5��4��2�l�u���w�w�ۤ7(��#��}I?���@f�P�c�dzk�*ѱ�P�͘s~���y8}�{�Ʋ�f�oNo?��Ao��M}�I��v�K��rڍ5|�w�?;�������ˣ�b՝k��7��K<=^sA�8b���Ro���{-N� �&q���B��N~A�ǣ�5%�D�/��m��7�tu�Z�6:�y����%�v�+	��^��MN8N5`��v���D����#D�]�gR�ԇW.�"�m�d�S���x��Y��l"tjB�\Gj�Vu1y� ��G�~�{��|y$�t��P�%�������-ӡ�<�����\��d�= �g>��	����Q�.:�92�����1��/��e%�*�j���6���z�?�x�?'Q�l!�Q!N��G��aF�œ@�e�R�-��$��c�	�M���N�<FL��Ad��S0s��P�m�"����3m^���c�P��=<<�M����>Ȑ�;::f�D�ީ�|	"79pbK�D@b�J���b2��65��;�ѻ9'�� �� o�vVbE�G�#o�!��o�;
�ƿ��\C"���=}�0����,��/�[��5s�m-"�/z-�g�-�w���K��J	�ԩ�mBW�
8�;[�O&%8���m^�>��,_sxZ��f �=����%�����7�b�SXz�~07-��Z������L���N$�U��o�'(	���8%�. d;\b����������J��[vg`�+&����-��z\��$։OĨ�i7HFX ��f<�<��u�����녒�{c�l{nU=�M�u�R��_�i�o��r&B}��b��)!--���hX�E i����{c"��r3v���~3�<{�X��ɨ!�qΛ;��$���
�7�o�NB��T��,�d]����������vj���+���w�<���vkekS%�	mr|�5֨g�o�kz��ٹu�NP�v"GR�o��Ԃƛ�"ռS�����
cn�	���s8���3���]��o+w�V�QTcc2b�)$I������eH��W�Po��-�� rІG%�^=�z�����v�>~��;�ޒ��B�R��D�v_�13��?����G	yoC����6h��s�쾡��^�56m�hX.�6���c.&#ڍ�&8z50$dD�-,(C*6����uޜGhe�3s����V�K��r�cuW�G�H������)��֗���L	��堯�h�4�T�$gz�-�%D�NG�b��E�������()�j�c�]mpdeFX�i���d�u��j�=�]�$ث�hktW;H�:f��'�;���Vŝ�v�G�б�P�n~:�s�[�����r���.'���S3���%��m�Ytjt�W�wWAנ|�T���x]g��ԛ�}����,�����O��-�UT�N'�Q���%���RRVL��Z��-�r'�.�m���?�C��� J���9K�ߚ5��`�?kN�À<��Xo��}Z�'�1uFP���5}׮]�!b��T�S,�TrN�}���rB��0vr�w�9���Ђ�}�:NΔZ����
�]����?][���m]����a����n�dv�)�:2�\�-��84���k:��N�x�y���y����u�~H��z՜�|��D5@����׾Ԟ}�~oq�%[.�������q޼�MkkkB�ćQ�Wet��LHSpw3g��l��!RW*j]�0�Φ�Ԟ��U�"H�$ ���:�72I
{t��2�V?��1(ޒ!y��C�p��<UX��Dy��$(�uu�kH�kV���s���ۑ7���t�$Q��~%]��~�+�)�����@���yG��f��V��Z`qA�o���l�&�S��	�����0.΅z����e�c<H�������$k�m�:�@��<�������F�bx����������8��_��cև�����<򁥪fgg�ԫ:�PB	�׭�'@^�[�'5�u]-� ��������v�{J|��`���q���%J��g�0ۧY�s�a om��)Hٴi�7pz��~��ޥ�Bn2�$ۈ��<�s����7�2r4_X�B`~q)d���B�`?:�[��������Nݢu��>�ꨠǷ؎�L�ďO�:śL^Ov��SU����P-3��*�q����5����H �:]����
�Pu��
� l��-���^������)`]oMu�>b����~���_πQR��LuU���	�dr�)������}�Ҥ��b����l��`8����uaΪ�b����aee��7V<"r�I�(*�����>���o�cMml��8��v�� o2��RA�e+Q�_P���1����;�Kb����� f�+])!�Iř��t%��p�}`鹿�)$(��"Z�� ���ZT���
�ؕ��;���7�嚢SP'\�
	6qq�VJ�r���7)���⏩��W����\[����1&U����g}�q���7���r��u�����|1
�S�a�-��=�e2�\�h�
m;�$��p����[9��"�Ս�XJ��ssq�u���sfm���}:��x�{2Ȃ�/_���.)Z����H(z�P����Mڐ��O0�*v�H�/	ޖ���p���"{#���z=a1�W�_�;T��B؆i���0��:^��M��%q�01%"ۅ8�����bd|��#�#��i��oR U��ˣ�z����i�I\�=^�]-Z��ʫ��V�ᵠ�hK_t�kV$y�P͓�?��Z4�bw�ƷR�!k��ԍ6��Xn���fB�p���Wmlx{��[���ץ�r{��8��g@�L�QW��2c7�;w����uVV�y�C��:p���¢	�ɍw����F�<�)4����E�g?����� T��?R�-W�ډ�eQ�a�n�DH� ���W��+���3}`�Pu��PQ�j	���]�%}|3~����\q({"G���%GB"��	�ѣ�ǎ�Dɚp����gP�j�%����o+ ��՛�4;��ʷ7�wvzU��VT���să���нڈ��M<~�9f�]�"˙�*z��GD��ԗ,��n;�t�֣��ѷ��Ft�UEV�&ŀ����|1�����u�;�yc��84�
H�ן��5Dx
^͚+�:��`1���)f��3��Vyx�A�"4�99x��'� 3Q���R�e�|k�C��✈K'�˛\|��,��H�S0�!�y����](^	yf��Z,�R@c��9�s!�st�(���qO���z)y�J��֪%�~�e5������&�%��Jy�#B��H��% ἅ�K,8���3�N�UE���],���V`�܈�fxG#�U.��|�k_�ﻍ�Ŵ^�\��u$eQ�mմF:��8T���wG��P�H�xx�G! p�`��f`��v�o�+L�o?T��#����	f^��%ɟ蒘�b���:�s��=~���y���q��7H<�3��CWD�( ձ�1T*q]�s7{{e��(�\(���k�06�*S]$�}�z����o���_Q��������Hvv9]Qj��3�(	�vb��f�ӯ0��P˼Q=y���#��B����`E��׉���a���"��^�a�eĈMm�2�߽{'��v��H�z�6|u�0~6����7'�PO& f�͉�S����4�xM�?$��6�H̱օ�$3̾�<�0յ��H�.�(�(�n>�׽Ie��[���模IIg���A�yt��k����W�;�j��[%���ߝ,��\��y���a�1�%Gvg��� M�G
�u�����5Y��;*&?w�P��/Qkq�.%�<g����wE��aˀlpU@�R�$v��9����f�(�e�wo�Pa���7�a��ꗯ�-W��oס������S之A�����j�.�P%�i�"����RjozJ�v��0���zކB��#�?9�0R�Pl����c�w�����̒[��ّ����e��E��u>\�F#|t]@mW��(lƑ��c.uޘ)�i�h��K��Ϥ���%�b�T����؊��k�H�^v�������G�J�fO�WU�V;U��1Rq�E�a` 7~�/���KEq��d�4��#����(��ޑm2b��j�0�:L9rԎ��66!P��b��T���Iڃ��xP<y��X$��m�U�DS�׍�w]o8��0��e��
e0� ��|�S�EJ�x�v��O�[ن�c�?L�XFi�7��#�`�u�1 �:�[�OW[�OW�溳?-��ި��d0�I �tXNz}I��*	q�����>����?$x	�z5�"�=����Զ?s̷艟��G�26Ө�a��/1�Ņ0�\`��i�U����U�M�|�J����5t("�U���*p(l���+ߝ�ï�WP��VI
b����L5���\y>J*��O��� R��U!�<��2�6��ǝD�&�JO���VX�H�b�F���-�.�䭛L�]xјn��{�7D2�-���s3�G[�D�o�������X^�ΛSà�$y��?�5�Cv�_P���ޭD���F\����
[A�����.�t��b��d�c(��\̲��Jp9暝�-<ۥ~6�}c���n�k�&.)r���}1?d�z2�:+���r"��'@ۡ�虦`C�x����OC�!�A������{�y�p_�2'���ʎ��0�%g�J'z�� ½��X�*����<�)��~�#G�r�T۔6}�:� ��Ě��_�z�B �� ��ߦ�Qae�g�T=^�4�T�������?gO�Ȍ�����L�d�]�������f�p�{��]�j�/�T����=��
fpl'o�A�~R��lu�j�oZ�̲%�����/ q��+\4�Ț����H��j��c�}c�ϡ�=�/ὑ����1�:�����<�D\�$����ҥY�+�y�F-�	!�x�Ӄl��
�0�N�TB�"��Dא����I ��9#���P<��6���s
��Mtg�r9���׷�"�n���Af$�ɓ'i��)�,Bg'(�k�=�h7��F��x�yz;Ea��U��V8�H[����� �q��Ju���B����1p��NP�Ł+-�ս^+v\.��_Y�إ�p$>	�a�'j�y�C��8��{B)!�� ���]*�pM��*+���XF�w�Y�r�0�p���`n��<�*ԧ��k���ض�B��7o�0���Vu�}5߀�O��4l�3���{�F��X�z~��e�sXOs~�S&v��6�<k)ܱn ��<쎐�Y��z�I��_�mU���K���j�]�j����	!fvE ��mj��m��ߩ	�qv.�n�D�Zy-�F�! ��@<����Ň���c�{��q,�\>��|Ȯؽ�U�}���@��Ŕ�{B���'�3kGlD t܄��ٖ}u�;����(^Fb�d�;�G�y������^޹���R��<���������Dǰ�<�v��_�D#���D�F�:?=#0���^9��Λ%��rI�|�-�^���Nu[�����`�uި�L�Aѝa��q��p�hq�<��D Nx{a�n#k^-�CN��'���Ӥ�w _"SX��7�I]ʂ���m�9�(����)9'��޹s���T��E6Fs2���-, �=x9����B����>�����q
s������Kqa����_�'�z�t��9!ov���P���h�By�Jǭ�o0mm�9�s������#�U≝n�b��$e8߭<�)��9-�6̺���k9��nn��k��-��v�/�|2��A2</����0H6Al2�D��a��P⏶ȣ%��]��g�_� z�k�/�XKhQ�m[C��=��o9����_Vyh @BzO���̹Y8s���s��&�'0L�ci���6C��W����B:��$��Ή��آ+���˘q	p�|7�M�9ߧ Z�;n�?�hY�hHފDB+�p�'KT��~���p�o�,ME���C���IF�@�����r\�����@�Hs�����%�P���f�����	"/����!�ՠ�v=:$(�9q�#a֙u�߇����4z���zeFl��iG���a]�c0���1�-�bʜ�1�۳\�[s
���Ȝ����z�9Xz>)�����
Գ�c��nI��~)�`7��љ�K�����5�:���'��<d6vF���bx�F=��� ��I!�Ο���]j˔,Ti�J+a6s��puT~�n���v��(;3�^�Ϲ����M���Q�@>=�P�˺�
5��
~p�Vfu�y�n
>j�kfz�%�V��f�#u�����rʻ�S����t�;~F�CX�t��Ny��N i��(@V�L}��t�$�
#��z���塓��(~��wyB;���Ll0f
pB�c�6-~�A��t�t���3���:�ر�yK��-|��JC�+�h2B���l����-qk�g���?|5��ߗ�(����FfEKÙ[�9�o������a%@ E�L.,~�����o�N8��i�ph'�i�I�`��]&��y�D.� V�|,�04���Й_��rG�7R�K��w�G��i�'Ȭ;���rz����4���3�m��j��d!s^�l\{.�W���5�$�s����M�X���r���cv�ŢЪ�fƘ�{�C�^W*w���N�xl{�;%��Ֆ�_���x�B�h�\������3��.��eAB�KJj"Ү����(���I�Ӟş�0��$$?B�@�Z���0.����@�;�Yy&�%�Ӡ��ϖxX���̅(���\{]/G��o��Z>��!i ��@B\]���J�7l	b�h7�'O[%BN����F,�U�y
�c�5�͢t-h�"\�ƕ̥�Т;���z.��[�Gf�A�vl��|��~��&�E�yy��?�9��p]�i0̻�r=+\��n��z��n�M9aJ�\.�xg�!��:	7��`�㺋��yO�J���^�ҫ׭s�P�6�ה3/�T����@*��.��t-Vg}��c{j�ut�:
�ez9�����p�i$�t}��b�&|�]�ϲD�N�-��s�cMM-R�y�s�k��u�~F 'f��\Oy�Y���QƻY Ū���򙹺m�1�A�X�]�8�8�p��i�^��w�������K���u�g�Iy{�{��}D�1Z��q�bM�m@ ���]���Q�#@χ`P�6ס���P������M�s�ӆ�pF���~|�y��3)��q�#|���ܰ�PH��g���j��|bdϲ�@���E���v@*\^T�$�>��y�L��IW���6���xcW-:�,���9��x"g�)�����{�Y��<(*:zo�L�=Lt�1�ͥAR�c����QxE�>�D��6��؅��*�����F\��a4����K�"q&�ಒb<4��Y�(W���(�$���7��s�3D�T�Y!�Ӵ��Xn����n�-ֆ��t?�V���}�:�\a�X�a~�16]�d��?�aI��C;�-��u��\�T,�wf�J��-��ޓ��4Ϸ�+C�[t�MS�0�_˶1�QI�e �r�Q8��?����8=�rr�G�����R/����fUߦ�k������Bj�v����M.��bQ��L��Ǉp/�֧�0�� ����r��K�d�8�x��8�|�܊]n)�M(��	���7�g�}'�,�����A��^ۭ�39��9�z{�q� ���V�||��s�/Dn�(�%-�6����aj���G�R��Y���-T��x9�O�Ԛ�ȧ��=��˷�f��H����TZߎ4<���Ә������j��@��{�m��5��1{Xdĭ��V/-f}Js���5�K+
;n��sU~������R`�&�ݞ����'��t��zQ\�rň�[BB�{`ͣ{xyq���lAU��3�&��Y���/���v>Y�i���wAܱ��ޜ�)�C�#��A�z����Sn��8{v�7��.�=ݵ��K�r$��E�[`�R��V[$������I��f�9�{�m:�Ǧ�a3�����:�q�x��ͪ�9�m/��
���
�M6�=/c�I�7s�{ʁ0w �K�� �9Lz}42YK��E/����8-�F��O���}L�ၲ���8�_�&��)廳o�X�ȣWm:��~C����St�h�O@�/��m��~�b�� �4�ͩ���/|Ý,�}�����Ɏ�F���;��r���ag�J�S�O��J�_�R��� �p�o�҉禧a��4ІA�@���z���^S�o�ʇQ��?���ܥ�g����ƃ�ǆy�=߿��7�Gvn%��׻J(�{�0�뤾��g8+�ȵ��,��|\����W@�,�U�e��<V5M)�];A��t�,��Z��n�L�R��~��܂ȁ8�fvs_}w2��h*`o��K�����ș{s�J���;~�
A�d�x��(H�~,�� ;���P� _�ts�OaQ�v0��-��d�)K�1���W�0J�3���$w������&��_z��]+�T#��a	�����4�H��0��r����K��N��g^ɷg��wS��jm>�=gC�3z�*ʊnvQ�U�|��jN�9:��q5[�k�6���ͭ�M�YR��p'5o�k��S����{'ϰпA��l�����o���ZN��\�ʎ}�S)�%���I�����'KMf�d���w���ձ���� d2�2!��=�Sb�Pݻ�:uu�ȣ�6tˬV���_B��j�p���znA<�Y]g3�� �'~o0f�?�E��~ z����*�i���Q�!�YW�.���mF?eA���Afdhf�n�fq�u�V]�դ�0��K���uE���ض��E���-�?���l�a���&<�g]6����:Q���i_�>����w���w���˜HF!^WGJ�)ySНc�8��1��Rwye�4���i��Z��.�e�p�qn6��t���n��$����[[�.���.�c_�E��#��Wh�l���W�x�o;�Y�C��������Ͽ�?�pc벑_�|�7���=������_�PK   �EX,��2ϙ �� /   images/d4f65665-9cd5-4bc8-bf69-d8b87beba5de.pngT�T���?� !��-  ҭ� !ݍt7�TR�[JJ�����Mw�;��s�����8.`��o|bf�O9qT"T888�O������P���?e}A���"J(�?���g������Z`_O�̔�CBǏj��6Ǝ}{#8�lfm�`�ok�lco�x @�
N��{%���������qr�ky��Ew����~F������Rƾ��M��JFN���edxT�R̭K�b
[�-O���*bna�[Om�ϡ)S��:���DG��O����¼�j��zϯaN�oX/V��P|{���Q��B�F�x����:+��}����y8���y�<���p�>�ӈ\;΅�������w ��󯋯����T}˼��2�X)N�!�t>H��Ʌ'���Щ��'(�
H�O~PÑ#&�G�~�3�p�k��Tث@\'�������A��u�օ�2�!�C��:�X�4�a2�^zb����(����&��˵�v�h!�J��4��H�ȯOi�7f�g���!�;���b�i�Q�d�Ә�3,I���OΟ^!N�Y"��'��)��w�S� �{�a)��/���$������!T�`9�>��(i����i��ٗ��}-��P,(!�a�ͬˮ��f��o<����B]�$U������%O4|�I��7�	����[�W�+��"-��]���HJr<A��7\��#Ŀ��ӿ�`�G�O:}qv>9�����_��f7=.[y�X�Z���n����?S�i��z�n���JW��G4�u}����慴�JG��(j���#V9������꺉�+ra���Բ�z|�t�h����Ry3͉�>� e?�w�Ӻ�N�<!���Շ�<�A^���}�!\��w����;���~	�opW��p!�v�#p:4-��ӊF����?�Ӣ>ԛ��D~�M�x���xD8�
}%��/���|�=�9������͍O�Xg�h�����P%����X���9n���2���8��س_�Y|���2�G��x�C)Oa#�8�:���;U����i�;����3cWd���p���X����H�����|��ζ���ݗ/_nO�W�,q)��K�}�~�"\��\���c�f>���������M��������ޞ����L�Qa��kf�|�`��I�S�}�
C�:'48�'LQ��iii�����$�[����u�Q�SR�'GGG�
U"#"��eRpsǮ�	{I�B�E&�����r�X�˗��&-��������	fS�mk�#��$��D >x!�jѼ�Scc�������O]?W����y����O����ؓy��S

_�*��اSN�Ӽz(�* �ޕ��ϑv��1�`VVV�����9���ȐҫI���������甒�D-))i��|���揆��~��5��v��e<@�A��l�uC��+Dȿ������7�*�������sp&��W���Ե�������u��rY��?EhB��O�� �ٍ
�]{⁉���I������#���vg�Xv��)O9SR��J>5M@n�J*��?~��������L���|��D�j�J�y#7;{d����˜Қ����)�n���j6jxXng�P*�^���HfffF��%��d�~g�.����'�6��Ń��-���l���~M�d}/����ä���L�ts�Z[G�G�M��)���@���x(�J�/�|��8TMDMd�y�#t4�l��j����9��� �gh(l�Ps��L1��B,����,�%E���'6�ß��<ί���t���x�5�J��4�@_e����VX�_,�-56t�pgmo�:�����_�O����+�E<W���p��;Zi�����v��<���Tշ��ew���<�8�!bm��&`I|N���j��#�>U>Z�e?�?�,�����>�Df�(�v=�D'`��^�}��y��렣�c�(-��|7�ʧϟ��4�l����Ǳ�m�qa|N䢦�빒����YMLLj�"����t�����&�����)��b�!��;�d�|%�m>�P���S���^|�L%D�\(i�����a�#IPLxxː�c �t�kΒ�K���R�]к��.&�4��J���B���H�Ӽ�v&и��������?8.��)3����;Ι��<����.(-A_�'�,���/����D������]�YYY%�mH�r:�ԢC��}�[Ue2���)"b�e?2&�q?Ad�e���3�̀�������*_)
�`^�7�Q�2d8k��� �  �-���X_�	��Ғ�t���`R���w�D?nƖ�����D��/� ���B��sYQ��B����9��?9G�W�� ��C��2_m7^����P�����ݯ*Ш��MyC*��
��� O� �#��&�Xy$�������e���'SK����z�-Exx�d׋��J˞��>�<�ǩ����%�{�p�-ET�/��%�I�p@9d��X�Y��aԩ�s�<�#''�y�. p�<�O�#�ae��\�,TlZC@S'��>m߱�!Z�Եdf�(u�����k"�$q{����i��D����V��Dn����g�1dbb⬵�7 6������a[�ཪ�>:>��rq�~��^ݿ��ׯ?��oE��-�[442��$=Xj���eUW�ٳg�QxR�;cc(
7=3�������������/���h��P��-ֻhV�$�2�{�*��0kK�NY�����SY�s���Z���sT1荢Û�ab
p��y��8��K�Ĵ_�[ZZ
gko�:2��"���&���Px�9K*6[�ƞ���ͅ�;Q�J_����QV�Fp��:�fC��iԃ^4���hL�_ B��$ ����+������@��h�G��6D--����7�������=���i��I��sU�Ѡ��S�L�>]mg�@��o=$xIb�p�>tڊ�r4&+�{-�oUs�G�����d���4�9;sL�UReѥ��(.�Д�RX9<�t����WZ�+އq�-+c(�q:^~k5�@)���!�gL�.��rQ��I���1ږ��:��١sU�3h�D! ��s6Mv���222�mW�		c&B%U��EDDrU��83�3Ū�������rdM�*�F���v&�ˌ���
l�K��"ie�O\���� �������ly��?�
#��
 o ��"�&k�����}�f�pXL�:�~����$�(�!�wf��qL�5��9�Bw�(fe��fȡ8BX�t��s|z�v�d��؂422R�Ç����[��?|� ��~+s� �8�/��l������8��r�{+ZUg(�DEE��/�"���`<���{$���l�m�H
�#5L�!�^�� XR���&� x�8��NԄ&��A�`k��`��CY��)��<�����~3�4�Ws5�*4��r0{���L��f2Y�^]��Yu�{0��� �\��7Z��@����B$��PS7ݴB�J�=�5vkb����nщ8��n���.�l���U�'WWW��`t<�?����ޫ.lL�zS���uo)}-+c_YYq<\L���s�u�윜������Ȅ��S�W�O-��� ��t��%p��'6��w�3΀�����{�;�pwu�r�淈?���R�$�L�9YYl ���^}A�NEn�ZE+��v��R�l��_H $!!qوVu�-�
�_������������/6�(X�;��>O��(�}ڪu=�Q̖^�;lduE�BDG�'�����:�
*�����E�'��`�ݛ.G�O,��� �����t��]j��2�'_�]�	���v�]� ŷ�Pm������<@F���U7\���@�ŅG�����|����mԛ����J]���`s�NRwF@��{�3���;	��_�+j_���:W�ߵ��� 5�:Y��(]K�L��گ�,y�2�FLL���{b�j�����6�!,P%�������#�X��l}��~wq��B��E�d0n��?&����*�"C�N��a��ι}q��"��P���0<)�s���������C�o[gg��r����ݏ�B4@���U�9B.��h�H��A���"�wf��!��
t @"��z�YL۽�7puQ�
�-"��>� 'JeƟn,�m�OJ�Q�u���x����l~!��ܹk��T^+��ɮ���P\\ܝ��s�oUY�A��Va�7���iww7`��3tE�ORC���D?%�^�d�:{�B3��D��B�����l�g��b�Ь��r�Ȟ.�V9 ���j3�7����>���}s��|e����G�z_��똪�9����Z�ַ\KUu0��n�u��ʕK����h&���H`|���5
;��pum�=r�k������x��-bUm���m�	o���-s����ߔ�3���6�Ӳ6N+ )CE����'Bq����(��ng��!��@r���t
�q���Ӑϡ��07��n�����s��G�Ȭ��XS���q>.� �I��Ԩ;t��ʥNqq��Cc��e���.9��^�ï>�ZLa�5�G��՗?�?�'8Xt�$�B��r��td:h1���F� ��T-��q'�xx�0����?\ߵwt��QfP��gg xso�]ߑ^+�T{q���R����tO��0��ȗ@�N�����$^�8���.!דש^7t�tc\\�w�.�EX��t[�~M��:)E|�oުȄ|��s0���@���]��N�d�������r��t�ێu&o@�@B�sZ�P2JQ�,��Ւhi0��Ä7�wmW-P{ˬ-�w ��a�	Mlhh`�틥L1���,5`�agW�{q��30��uGU$���v�]�F�-��B��0:Y���o�vV�+[Lr!�R6���sU6,'���� � ~�qD���gi%�B�+�
�׶Mu_;�on��+;?�_}[��%�L�9 �P�e�����b���"���H���\�Fe��,s#�2&�qUcc.��j<�X6H��=&TVz�^�Pe��B5[:^��x@����������5lZ-�R�D	�	����w�Y~p��þ��M���3�4ħwק�I��!��	��2%A����>~���%ɽ��r~x�Ų�<���U�'��*щ���:��d�f�1{�T�ޓ��[f�|iQ����yC��"ø�&����)|K��a��%����i�˙�����TO���[!�%p�m���X^�&`���l�ߦ$'cL��*��YN�:?�꩖���0 �\�� n_�A���x�;�K<<�c���HBa/P�3qb�hO�U�u������ɰ�������O�l8̿C�r[[X�&��=W�}�kq����L.\�=���с��/L1D������ �e&�د������	���!�\����y� eT�:���ۇ=ݳ�����+������Ka�����v��uG���l�Ȑ�!��ω�����ū�91([�+1�54@�P+��jU;F*�O� ��t2y(�)�T�z��/�dD���n��&�ba�7C%�i��:h�/�z�M�]]] �������((�ŵz:$LK�u��DL����~���>݉amo]/�c��[�/+����>�*SBj�ռ^,���t�2���K��l���[jZz��,<�X�Ö���@T�	y2���l��d�?O%�m�>�t�b�����B�
��飖���b��'���=�4��:G�K�/z��=6sZZw�]�l���?�O��w�_���g��]=�ԭ��	]a��L�����|lg��RO$-��,���=.b|�td!A.�r$�Z���#�0�a�Y�~��g�������Ps�����NF�80�ߗ�T]8r����y�� *>� �e�]�:O����<�?���Ӎ�"E�P���ܜ����cT���Z����Pt�vY�4�7�pf$�M��蔮rO��іTz�*���X��uC4
E&{�\���
���|��b[������`�^ל�s��d]�`��F�8$�!������Jl��2���n4�f���+�r>k6��N H	�igK�U�����Z��:0�H�*�y�
�1+-�*d�Nt1���L�MbZ���*H�
%��zͼ�_�*Po��������#�����\�`�da����	�l6�H0���[�^f;U9,\�,� JF�{�%baщ�}��-�fc.WG��xxg�
�4�Me[�d��Le�o��$5��v��(�QZf8Qf�������)]����baF�6Oʢ1�I��P'�9��������rs�_�.!tk��S���-��;X�?��0���!���<�z���� U���Q�{&�۷��3o��,MS2��`���B&���v�s� Y��^��*��^�?����ײd�Q�`�D�\���"�傓��#41�x��Q@�[A�j�[�=5��|��K[H�Q�l�'����]N��5GL2��?y���}��AĲ��b[� .�G_�눥ߡ�!V�!����L	N���;awK�/.�
�a��̮�Z����mi�`S�v2�����1�>�0�c�#wG�_lvt�*+*6`u�%���ё�822^ڱ��)rB��Ƹ�&}�Aw��X��B?k4½���M�9Ud����p��d���h�.@��008͓��,񘵺Ϡc=���'B��K��ҕo��8���7�2���Ȩs��M�������?�C���.rBV=8:::�����^}O |�z�YFuh�k,�xt~n�0���ַ߿_�����::¹�vG�߄�*�rW�ڔ��?嶆��g"�Dp�U����7���-B%Yy�����@*JK+�b��Q�}f�B���5�}���3º�2_��F�� �l?��D��3e&�|�oL�R&nK���)B���c"R�6L9H��_�_�P�~|lu�E�уר7����]����ENs�d���G1�w��q2��q镖�R��A�����X(I��)P�|�y�s*<|��ޘU�ҟ�9?A�	����:�m������ё0I���� ��jii
r�\E�Q��r^����z9� V��Y%�2Y�ݫP��X�&��/�U�7@S�繥F��N�$�T�w
`O����݌�:i�9���P�@M��撘�z�H��H[�1�������:j�лԲ��2:A������b��_W���&l7�l{�5-�G�dV���g�`�d���l/yVF��oS*�Z��Xt�����53�rR�2 ߺ�:�,,dB@B�����ɯ�9u$ ��j�b$6�h� r04\��ǁ�������::^�H�nxP�:��FjV���>"8>>r�ǐЭt1� lG��*��r�Q8s͓���F��s徺��K����������t���sĕ�cc��ȥ�C���&�a9d��"%8����|��8�7o~�z?z{{�uU�y{����mA�.��򷂏ݜ�7��1�k�%	/��yS=����:��:D0���F!��͢ X�>(�`^(�?2����{8�Z��g�*�V��dǢӴ0J���p����3R��r�$��S��ђ#8��H �6��V��U�R�]�������Z��R�1�?*��G0?�3�3�V�H  ��ws}B؟�P�T��G�/5M�v]�Hǅ2��������4�9,bE'Oh��\݀�[9@2�����۾H���&;av=Yf5[ζ��F�0[<����߶g�In,��m�A�GGr|��w���n��B����h�G����:-3�
"||q��:�|�oQ`��g��� t�ֵ�0�Ɯ�&,�P��n���-���>Q����c�VH���q���B�wj4��0�_�~EO�����?�-n�ߝd��d��F�B�V�����Z��/W-��ww��Ŭ=�v[��t�5d���ְR��n����3���q���8���Vm�AB��H�T�#n,Gv������|)7]!o{��JBB������H�q���?�EZ5��\�B���/���ݡ<��oH;����z�Л����f���荞�&P����vZ��;�� �97��Y��s{WD���k��F#h����i��W||���.̥ś����dffR��H���ZgJ���������ԓ+t��c�)$�(��uw����I��Ӟ�t�5.�:��.�^�G胚�,_7����k��m�%r�f*`�ι���~��v��<�7��/�VmZ�""5٨Ç����G�+�pF���Z��+E&"r���y +��M^�j��-��6�ٟ�aL�|�G����r����iܼ��i`�������D����,i�@�8���͙��ٶ��.���D�+L������q��B�ϩ��u���u^�o��r���V�x�\o�d��`!|��m��&d��E.@�M�h������D��V��m$kTZ�'���}/�^��;��bh0:T?j|\����{p�j7�-A��C	�T�.֟���4M�!:[>ѯI�� ���T&R��i��ԿT�5���:��N1����TTA!s��?8�amo1���b3�C�r��V�mK�m�

0ll5�����_�k�7xl�}@X��M[�ڜ�+A�͕Eӹ�ŧ�Ԥ�F��n�+�JKj
��|MM=�.�<Y�m1����U�Uq�PG�����e���̚�Z���3D�re��lR뫫�
�%��~��?Wi��?�}w,��mS�P��52Es�!{i{3 � ˁj�d[���!i%%��	+���H�(/�@?`�.}JY?�����uh���޷q�����ɛ������z>�]GO^o���\C�8R��l��m�~�RR��egg'�$ �<
x�׽	F�.�p�dt�#,=������'i?͑	�!3��Z��ک�VZ�_��z]Sk�9O\���y�٫�G���TH�����B³��9� ���'$�cD�U��x����&��	�i*�l�B��Jjh+���0�"#;>7=H~�$����0����D_���;X� ��`��P}M�|�G�B�>�r��y�	C##��sU�nN�r�ʑIF?p75ۙ��q|����D/i˺��W����m�筳��6F����u0�0Y��۸9�g�wvcCZ�n�L��aU��:RA�N�B��� <K���6��P��m���A��;vy��<BY��y�)�YZLs�"�yˬ�I���H�B㾋�K�doCo|5���*[z'(�ʚ6y��3l�m�ꃥ뫫����B���@)E�������S��Q$���+����[��n~~~����E�bk0����1U|q�F��ى�8���>��m��5��%eeLg7��Ұ� m1X����u�e����h����zn%C\��0j!`&������"�N��z�W�����Jo#o�s׸r�EH:^�LL̿�K�ts ɦ{rP��7�m�@˫Z���s�haznnu?k.��bM�S
�X*b�3�*�c-��q�Tgp�;d�@�s	��⥊h�ց��a���RV}�y�߰���p*p�����D�#��'�FpIt}��=��`�ֺ+��lw*���@����nk�Yó��_q���<�#�h����tҧRy�^]��:���L�
�ex��ys�&zC��#t,���>_%��,R�.�_��|�5�>���4�Ӈ�ŵ�Bd�.�q�9L�����}���hP���k~��9p��o,x^o(M�!�N"����raǗ;ۏ^c�����!�&>��Z��_J� ����p+f�a8�M��.-7R�I��ŕ:���s�VG�RQ�����\�O�BK������j�3`e?��9Kax��wBI��?)�w �+�)�� ;��,���o1~I  ��u��r��8�����;�u2Y��qԂ̧=W`��@̹}���*����9�Ώ�}�Z��B�w�y�F�������
��I�C>�������t;�I�x�ͤq�OR�w�OhD���+-g���=|<�����bb+X1�Sݻ,��)V�q����6a��n]L�?��M�8���=?��0aԪ����ʢ�Ӫ��g��>�궜�C�3p�G�������<ke��wq:�)�JJ�G5%6����X��tz�u�GL	 ��A'����Ź�f���<is{��p�ɛs3A:K�x�j�H�7�$N2��h���¬o0��R3���nxxgˌ�ZD�\�������ov���ML� K��~H��Elv��y
Y��/����(��ʹr�����G)�kj*9����و�D)11�����F�D@�̺���T��c(�Ѩ,,,�����#�����...i*��WGa����}<<<w[��b�aST�"j���t���BBB���&&�����k�$"i��VC�!�Y6�C��m�߮/��9��;eld4�����2び�T�y+ ���%^��	ٹ8
��,G�o�3�b�%���g��ي�+�\���]k�ҍ��HH��Kn�D�>%��^v}�m@��R}�XW����6�����o��#��T���	��Jq<�#�����n��}��d$5[��oO�wYW�u_������$]�B�+((h�E�?LA��8�,�8tm'as��v&�����uV����C'�(�e
H$��
0,l�7rH�7�I
L���@�d4���:�@��׻F*���vἮV�S2������R�.�����9�DC:0!�#_5*�W��ւ���aw��� �-�*?�h�H�6\�	��{���f��������MO��C�a1��yE��$��a�B�t5��V�s��'����g��-Vv��s�?�������ۙ8�0� |��Pp�m��`u'��9ךk�w�̣"o���2�^��;P�?~�h�i�٢���M>7�k���Vbd6{[b?�/x55d�9Y9ق��݁}���67u3k���5{��U��b3&��&�%-W���� �$wv��tz6�EK��$VrqE[ZZ�ᛞS���c�؇���>��4):>�m��[ %%���!_YYqbsؔ6����Sn���������.�PWW����b��NII���O6si�G�����b��Y��ܲP�C �}S{@�5WeC|��)Ka����E��*]�z��\t=T1��^[k���ˠ�cQ�Q����G���7��
H Ce�)�����;`9fF���F>ȁ�p��(�~�*1΀�B&����z��a�����ɂ�6,a��0�D�zdw����ǚ@E�m���N`v�C�_{=l��V�e;���ݟO9	m�&����a>�FC7-��t].�JJ"�m�*?�G���*�L��I�'��L$>`�`��^�]��H��ľ���ۏ3����W���U�.���U�w2rwwRG����RH!cf�K�0�8���y�'���S`%'-B�����=o�C�~��q������z��w8�����)��O� �d�����/P�D;߿�;]y�N�!>�]�[�h�d��SZ7�臮0,_�W�f���KK�{N�

����*d��YR�Q�t\My"�Ʌ+����j�=��i�א�</ ��qt�۞���m���{�»�� ����njп��@`@^���EA���[�Ğ�  ��^�mhxȭ���X��!�>����dr���7;U�V�<����l_�E����̖I6��ȁm���l��G��l2|���R�$p�W֟*�:Sfm�ucgk��P�r{Y������[���oK��Tiii��)��A�ZG��i	��ܒI�v�v��v69u����ɡé�=#���1�ͽO��oN�4��w�?%%|����1+'ւI׆�rUaH!OO/5��h�H���8$44[���9�V�@6̂����]HHA~o3C3��gS���Y�ft0x�v��8V}x��3���	��v���L��D�޵�~�㰌�)�E�����M�s�]>O�9ޭ��=����~���].���O��'�{l�#����x����#4�	5lll�*�mmm�[��K����|�KA<�F�;�<��$�4�����&��b�$0�!���N ��u�������H�@�"$"[ �t<ϕAn(S�FaWo �MT��XZZ�V�?[�	¢�䵰�V��,d=σǤ����X����ՠ A���j���g/�6A��%<"���E�24Q�f�������<lz�i��))�L�X��Z��a���� � �r�ׯ�_��P�O�^�p�[̝�N%XM���L5�P~�%l2�6�癝�dV�-K����H�,�؆TN���݀��e���Ǉ.@�g	� ?=�'T���˽qCSCz� E�x��Fx�9e��~�Y���x���xn�@%�WF*_Zʺ�%x]ꬲTr��!�l��5��`�L��~�;�~t1w�GݕӴ��?�S��Z!��?c9�b��ȠZ�j9�
 5{��n���̪Fͯ-~ȏ[�*W��$�A�֟�2���g����Υ(f�������~�l�����@K�/���?��F�@~9���Q}��>l�D��ᏆX�G̉��y���щ1�u�b��R�gx��\���l�q�:�A�.�[SS�T�T�xy ���u�Q�os��rg����a���>�XW�9�O��L��<~��+h[��]�[�u����\�Ax�Ƣ�]b��7?��t��3�*:�B�� w���L���%Ld'�_12e���L\�V�
2e��x���^6�7r��F3Hݍ"�Y;�yym-sʳ+�<�c���1����7��KM�r�@Jxx�������z�Y*�B�*T �e�B�z�LY߭��ɉcY�F��C�'2�cWG�z� �s�&�&/���_�xk�ɽ��'�Hv��7��Ц������i\�n�z�q'��"�V3A~��-��0��ްyE{g���<��b���9}O�+�zC}���իW������b�I`����Rw=���.��������so�)57��˗/?IH�LMŖ����=��(�j��9����������6�K.M��_d���#�ub��;d���b��
��� �˗"��ڨ�w�-���]R,��x��9P
��?��;�����)���Q#a�D%ذ\+b��uw,�@>�}�C+���7�����g�!9��=f�U��������0��~H��Y���{>�KW����u=�NNn�zI�^ܼkieu��Z;>!A�֖v�M��3�K�f��w��K�����6��#a��N	� qXN�����/>=�]P�]�0�ƺ!{�[���qe��<e�VV�(�꘹�g�9ϸ�ĵ����|5�>�B���w����qsN~�4 Kn!އ����m�'kJ[���@4q��^�ف|����p���CK+�$�Jy�����w,��SQ��\y7�S�T!��)����H�2�l�0s�vPf&����`��]LR��?������@}��6z��6�s�3s�ˌ��/�`�wǦ�M�/}|�S5��R������&��.�V:E  �U�:�r�fc�i��`7^�6-��*{sU���������n�:���� 4l���RGG�F�����K"�JlS�2_�� n����	1+����b���zc?88���G�,I܆~�u`_��"҈p�x�ꔝp��WT��{�F/�l��	�;�+��_@j�)���I�^���5A��"v��f��3�%�p�.��R<u�~�7R�c�����ˈ�q�v�G��uh��N��ZZn�X��pg�FZRzX.�Ex˜:�f�V#"Ȇ��-/�Q�eL�)��!Vz[�MՒz񝕕�*��_ھqa��76��74�ĒL��G�R#������T����g�a�e=�:�R�����0H��j�����~rUU�:�������'��o��Ccu�~2iV|�(�̊�Y���J{f�3N���zƌ�)��	H�qw�ii
�Y���6����r�>�ǆ�@��Z�e��:��͘3�i����������_gg�$�=Z��wrڸ�>�~� ���x�s���ӿ�U���e r�1����=ai�+���j�FI����4s�Mz'!g�o��k�j�t���Gf!���\|�kJ]���
2�߅��ZZ������{�4�=v��V�>ǂla1İ��1�tt%~�b�������-�^��h�,0�q?n���<��L�.�v�h�l�ö~p0����>�[��:�
yµh-�޶寫�iۻh_���$
.1$w$�4���OpG#�'�MO��]�IJ��\��� ��d "c�4w�]jk��؟�4�}ALL<�īh��2��i�aTO�J�t�]a�mY(��۷4�m}}�9[��333���PN��F/. �1
��\���mS܏�;��&���B,0/i>'<�"�pצ���KuukK�___Y�{0%�ȆU�+��9Br�^������ M@_�x�_.y� ��;켊����Ϲ��$#�����.����Ӆ���u�EșC��mp@�OR�{V��M�F���������P� ��+��N�f1Fs�c2$F$�gC�l�{/�@?իf7iԵ߬5� �A �)W�Q)mT���z�J��{:�i�l� ��3"~

_ E��P��1zƺ��N�;s��X�?�9�7Sv�\).&vr1g��=�Q�1M��,oo�t��r�[5�7�ܓM���;٪�z�k�����-�������!���_޹w7��0\\�L�+�8r[�"�6b�c��n?N�;��J���K��Ý+"v����o����9�/�k]a��̞�}8�ΰ����w�۵�S��g�R׍�^�n�?ַ��Ӝ_ݮO6�3e9�k�� ��d}Q@b�jA!�V��#H	����le�o]�+U
5^�o�Bq��~�Z-� Nz��K��KJ�wp0t�/vW�Y��P"�ùB�fXh���T��M�c�#T�oܝ�
<6��uo{I&��'�o�� �D��� ��T�Szq1� &}�X8-����C�����ݥi���雵ΐ�ݔ�`� ,r���?��ÅT��5��o9c��u����� �UO�	n���7=K��Z�.��~���B��ޅ���hjT<��e@��O��w��ە֦�'��DD��Ě8�^V��-RȤ
��8�lx�t��V����ys�c_1k!ք�*����2:Aڔ�o�v��9��ھcUa5�e�-��~��@�x�F,��XҶ�;;;���k�����������zp���s��/yDg�o}� �өw	Yeyh�9O]��lv��	4w;��:�x&vN�!Y�L�h���5��ysd"�����乩Z���/���K�`^9eJ|���0��l�.�:�"#B�GgQ*+t�ᐶ@1Gf�QG��+�d�Y������V��ۛ�{{4�%>�f�Zn5�'�:�mв�>w!g;1��2��S�.���Ƥ$��K}0j�������L�K��'���#�;�'�$�|_�������_0�i��&�W5�d$�9ї�D+�y_�Ӑ0W�y��d-Lxr{�>$�9��i>�]�7�x����)�%�ہm��uQǳ1,-rA������ |�P�.����(�	��Q},�p�@h��������X{P��6�.*!+�rT{C��=�	-c|��\y�8~^1�k|è�8g�QW�+��os�/94@�$x3�%�P�go�yw_�V�	D�[�,ܝAx� N���(ځ�O�f\.l3�[�4�z������t.�%mR2i�OU��,��Z!�������X��k��a�J�-)|��\�5��Q��ro��=�/A+�6\�Mutd5+'����\�r)<�uu���` z���=i��ņ>�����+b,,��(���"��/_F<_��35gn$���K��W�5C��<���������b��}��&m$�i �QC8�hw��6��w�	���@��7�=�ŧ@:�-n*�[�Q�`�mL��Os��|��<���y%�Y{����Ew,���es@]��_6�US!Wu(`��;ݾ������2.�+��n�ts�9�[Y���g�dy���L�m΄N����A6z�����B��#�*5��F���Ϣ�A��%���;:�ߊJ���=�.=��z��-ּ�ŕ"�.��
jt�l@~�-�>-U/���z�k��5���222Ҝ�Ruw�ۖ3���i+��P8�iR(����K4�У%;n��RS����#x�$>}z��_���*���f�F�� a�U����֭��@/��é��D�m��&m�������|��<arRR����x�a�vP��������Wei�Ҭu�Z�͙���&ao3��&o�4)���/�T��5q�c�t��8HMy����UΏY��+�i�����]&:��nh#]O�9���b�"%�A�W)N�ܥ�Q��F|�6kP��b�p_,î�ҁ��-�?'�rq��PJH]]]���9��IQ��s5�<� C"���^e&C�g�-��w��J�=�����59�K	U��G�uQ��f�j���}�m�]��*|}Mʌ��)ڧ�v(��.]!Ī��M�yJ�M�u�?��1���t �l  
�_׺�p:ng��#i>�!^��30]�~U�-uԄ�<=##�x�����k��Դ����; ���Icr���׍1K�9%��h;F;���Yt�!9�)�X���%U�������c	d�N^k�Y�N���_U���{j��lΙ?����$��B8�3K.9;�2��$ؓQ�
�r�}��M�d�[|�>��9�ԫ!E��p���/�Ɂ�x^k���s�@����#��/� d�acc���xw"UA-���ί�F��I0gy�_[�H�XP�>h��ߢ��wOT���;� �i��WZ�h)(�8l��8isss�9|u?���q��?��ً//���a���9=ZeԪ����E(D��|�S����N�ػ]�og'̇�\;���B�v>s���3y�ƻ.�S��E����.wQ5���%������:iVY�y�,O�̢(��
�&�p��b����lc������f��c|�U6K���T�y�q11 �V@��#�=�x��R�U�e)Û��*,����IHI�m�jj���76(�蠩�#��m��Q_���"R�tI7H7HH��tHw7()��-%-��%���]�l����G����̺cf����%������d�ܶ0���o��yGFG�����,%]4���"�:�w'WW���QL��	FFF��g�I{���Պu���zc�5ud����3%�S�-�kT'���ۀ
�'��~�珞����9N�A�2�7
O��
�8����Ohѳ^���Ը-�B���!1#����/��o��M��j{�/�o��E�h���a�p��u�${"��_#sA�y�����!���Cu`ݛ��ix������K��L�{X���c���|Z�����+�����6ȗ2�Ĺ\9��23�E�j;i��P�Mp�Ex[V�u�9_�_Q<c�2D���D���`�����'��?0� X�\��|�_R�'��� ����r�ڥohH���s����ݠ�qPSS�����@���*R�U�
|,~�]��D!��,]L�F�1�F���n��w9ss:CC�h����^��&�av���������pd@ �x���-v�*l���� h��k6�_r�GIcc�Z�
��5���)D�����W��E�g��TV��0R�, ����W}�3�W;c�N���iZ��L�T�7=���I�{{[��Qߌ���{,�����5]�7�-���oj:++K��뱶���䈍*������ԗl��*��Q�Io�Z�z��:�R����M�D!%��{g�،�LD�=�s�0�>a�p��bo�ꏈ�ڰ�y"�X���/r�r�*t�7�[����q]o�F[N~� P�v`����XQj���NWP�auss��亾�J�k�N�Jho�O���{s����5�p���h �W���Q��Ah$
f��	��6�e�Ė�<z�ƽyR�UU�����#��as0���y&����#���T[�L�m�0�Ӎ���ga�����F��J/766²䣥)s��>?p��5@�����5�
������|[��״��ҕ�"Ϩc�K�f��p^��hJga$�$�g���L�Q�ݵ���;���C��F���#��|�P���ڗ��W9z���^�R�%*LU���Kk��頍��Zî����X����ߗ�a�.�c�.;cy%�����.�v	���	F4lx����o��1(0���z
196���o��8mo�'\ ��es�����@[2+�̓�������=��t��x����*!w3wJ||^�&�p�=B�M@H@=.����8���p^�����Lf�y�{�ny��:5��C~vԹdG��`�J�/�̇\U���E:x
�����n�ѶP9��_ccc��JF���9���P?�ֶ�R�.������}W:�	���V_���2'[���p��m��Ж6J8��� |S�Pď�������ԡi���#e8x�T	��!@'�����ܝ����t�)lUx�L1t�Z������Y�hq����5�&5���)�%�./)Q��|�;��k��8p�4-Q���#��� Gk=�<$N6O���>��0��?ԞZ��0�+wDd����?�����de==˘W���[F�#MI��ҿ[�����T�E�:DP;���������sZA�}_�jW$�����`r�ޞ����ǃ�n��g��;p񟍒��ؼn��m� �� �Q��a��϶�O���uA)f1�Tn���$�s;����r@��k��H����==r,�^gƻУ�4���,d��� ��z�<圣�B�h�CS�,i���O�0D���O�>-1"���@`�g�X�8��Mt�ވN�ST�P��qxh���^�����UVoғ�h���ki��56ڌtK3o��7�R�(���|��l��1�� Y�fW"��[��IAM�bXq��)�r�Y����3:�vho����w��Z�R���V�+�$��-��>d�7\��lsz����W��É�4���x��e������לL��߼1����Ehii�fQ����s�r�G��#GS�a��Y4G>���/�hG0����3x�U0������oG�O­����_J��h$`�._���	z��s�S(��烿f�[��t8<n�i{yq�Y�i{�!��9=x�5[�<�"
�?���-uӉ.1�C\[^n�Ք����J0�H�A�j�z����y|�Ѝ��v"�4��P��S�� j�A���';ׂr�#l���X%vZ���t�Zm.qSU%%b�)g.����h�lE�nZ$��믴'vƼ�V�"�~.��S���P�Zg��'�Vv%���F��D�xm'ꍎn��B�d�*���[���nn~8��ӫkė��8P�	

n�T�g�o u`N����S��ҙ����8��^�ʒ��N��s��2�X�{X�ΰ�O/����U|��9R-l*��[uܪpq �իmI�D8��
��(#���F��փS�x�Z�k7�IEF66������.s8���X!�6V���9���YLL��r/���ⅅ��ձL_tY]�ƖXߢ�uѴjj�Kp32�}L�`�M��Z͔/��;	T����Q�ɉ���RIe������k>:1�eHLq6����O�������g0Okp�<�PS�c�æi���*Mc�>��'`�_����sHI�5�^�Ϡ��򃜅~B�܁�$�B=�A�T��3���Q��jg'���[�~�}/"�zwk=e��<.WζG���B�&�tuS6�R���K>�<�\l$��3.y���WГ��`.Ls���HH�5<��o2x������Zj�
�p�B軓�/	B�S|��@���t,gp���ܨ�����ЊMvv�z�%^���S������	77y��P��͘&����'�[2ܬ�3�Ԡ��3
��a�z/DJ(�hG|�L9�$ߚ d��Õ��|$���G�B)u��QZ�7+�Z�b��J߭��6����Iou������K�u��~��^�/(,d1�Ǖ]��L���2��F;���
�Q<yww:��>�w�7�$M��i*t�j�����(z��k�1
�M�Eh�*|��_��w� G~�d��B<���͸�<�ȍd�iU���tƱyQOH�僿����a$�;K����X�S/~�2����s��e��C��Q�}���L鄶�������p�;h�
�)��I̛�| p�o/��}���}E�i\޼��$��G.���"W�4�w��x�M����?�nl`�8����w,�R�iV���n�M�$Bͮ�]���Nw�.Թ�����oU��B^[����5�w�Y��i6Zq%I�LLLS��qs��.=G,�*�+�x9����}��#S_���s�	F؝��Q
��)�D.+d=:g�5/��<����2��"�{>)�mO�8�[Z2@�pvkIII�)k������2�y�"���yW"2:?w||�+��_<*u3�ۋ$�q��W3������U�����jذ5��VUquF�D��^�SR �K���&����*Jo w;��������α-�.t�K�0J��k���_��ߦ�7U�m�������vw}�S��N�V�G#�b��b�jy����8�G7�``�z���H�Jdߏ`P�f�r�*��?���/����D(��:�����y�3�4;{N!r[@�����7'��9%�D�ы�r,�z���e;��h�e6���n�g�u�����f���|.FG.d�������Qop�@����i�]��od���M4b��2�%�7���gj�s�BV(G���
��+��+��c@9�Dt��I3� [ �<C�{S&�N��$ ��A!h���,u9�#���*�*�(�����r�}�} �����~c>F��%�}��i����M�m�t��~t���;����Duk,����P�I�^�
�����Y���ssi,�_�>���zl�
�ϡj�#~��DkB!�ԡ3O%dj��g��dt�=`^���>� _~����k A��L���8�G\�ob�Q�~�6�[V^�n��չ���٭-�)G��/�~Ϝm=��Nl�-B��l�O��/�/%��s�n��GF�*���;�?�R���o�0Kg�444:`3�c���_G������j#�O��m_WC�r���Bv��+:B�B����`���$@b��T�~B U-P��tt�{o^�6���C0���r� ���::��3���=�����q�Q��y0��bDoI�Q��}�P��/�N��C[c�jh߿/������{�a��_ݢ���l2/Ĥs����Q�H�R'H��R*Щ��ļ�|'k F�3hs3���@�����t)]�E<��~�P��(�'�}�`�P����s�i��>��xxD�g���WF� �W�l���*R��斖/�w�\6�'�$d�?�dw�O5Y�n��C�ͭ0onZUN������1�i�\f�*���A�h�L�4�j���e]�σ�v��	�cM�S��yyya����H�K����D�G�ddj��E�[�s�p��rř�?���	�=��� ʗ�t�S1荦�����{�w�3N?萯Z��M2,V��Kd$0(a_�"���}l�G�>p*���A�ח�..] �J�����״�,��+��掎w���;�mק�
�b�⪹�Ҁmp1�k��j�*��#{�|	R-�$eb���	u|���ߠ��K��ɨuki�3��4`1��%) ]�P����b�.��W�nf��q��R/
���`�����B$�7��S�\��w_�$2K,�,���eT	[��Y�6��#�c��L!��e���lj�z�Oisvq��|������8�h���{4�k��O�m��u�g�d`���\j6���G���z�/�sa_��Ю��q�@Q���.f�뒧BW�ŧɞoB͇B�_���fGJ�>�b��<��u��.�/�L���7Ʌ��i���S:� �`�q�52:
��YV�;���,�R���K�?"&:^p[Z���J��h@@ ��R��'�LN;*` �)�������N.nZ?���tuu���k|#��E�����Τ�n�
>4X �[n2_q�����d�<���kco����^��Vgf�����8�kV���5�}��W�/7�k�J	Q)�I���Ҋ(�[/zE�O�ܑ\��iGDt�����u��74g��bb`�=��	���RJV{m�����=&M���	�'q�v�Lau�Jy*�>,A�oV����u]�Q�����|����70N�A$�


��౏��E'xt��g�n�p���=��^#��Ħкb?�zH�ry���:U���@b��"�M|��u��-�]CC#i#>11�����.9px�#�[l��e��@��r� ��3��6�� �׹t�ND����XA!hA�Qx�0d����q������	��/ii�Ǌt~����S�9SaK���r��!�B�$�0���IZ�v��{o���۟�vEJxz��'q�)qӑ_���K�@�_#"���F��Gm�V񣥧��,"�)V���)�U>]�*D��W�b��a�ޱ�u�:�T{]�������)�a���.d�����Go�����-��C�v2��/]�`�H|T�~}I�:��R����<7;��S����f�:;��"��;�.AYM�`t���1��4�½���G�����N����?����(�{<�d]�S�|2�T�WNӗ�RZ��x6��
�?�����Y3n��IIIG��Mm==R���_`��^8;�S?�;U�����o�kd���J��nL�F�s Ϫ9���.����jź�uΌ�I<~qq�s�n���j@�uڵ�%�wE�z�0��"�@a�70�U\�u�*/5[ec��9ւ���7��D{�ߺ@t�L�����|�5G0Tƍa�fP���4o�7�F�%���!Y�\�v���j0t`�v�hii���xazoƾ�W�~.��w-��1���p���S��!���rł��h^B~�o�疖�G�A$���ô�� &�Pɝ������"����p��vBq��4��������j�(y�����H��GѮ��ӗ�^m��dj��j�QQ��}��e�s�z��Dfܐi�<7�d��c�6:*��L��撊�<g
��k4�}���y���H�����VQKE��������a}�����ng�>>�X��q����_�ɀ{[NV��N�Z7�T'���x�$E�'�"i�	`j���0�����3596
<7Zqr�l���ީ�����p|�IqS��%���B�!�����l9vv�4pm��W�x��7*h£��O�����8dO���?ܹ9�M��� ��b�*�~R�i�~Pks�ǯ�VVf�A�D�L����8����JR��Ϳ?��-5�`��y�F�z� ���o�����[gh�"��'�z�P�kmc	7y�I���{cu�mWp�x�nw�A�
])��/��AF}��
�FVRRb׍D�\o��M�=L,�d�8O�-c_��-n���=��z �\�DH!�t�¢6��ic$��Ԫ�@�l����� eH��NI^�&6!��QK}����@�#ٱ�L�9Uh�pe�����~��n�e��n�%��x�Av%E�.��M��DN���щ�ھ6��H��U��-'�@�/�<ޒ@6.��@���@^c�g:25Y�7���^�ٙc���PQ�����5 ��ϫ�۞���ƪ��y�]�u�PSS�_��uu����^'�^fG�a1!ķaee���[o�T���H��<��}
		Idw���>l����r9�er(�����^ر'�糕�>�6���jM4_8��a_�
P�]�{`���ja�0�&����y8s��t�����?�p�Y�
���������c��g3��.�[�\7<����v�e u�P:�&/m����g�샧����kt��������|�m���0���Í	!D"Y.7gf��Ǥ�GkDʴh��U�:b��ͧ�F���V�i���{()+k(H��)\rDEE��.����G:{-���`��GO/���T�F.�Lq���T"=�v'�'���w3&�����7T��g��͉ԌEy������+i�I�m�|r��zP[�����>l�K��"111/s�BZL���RZ�m�/�|�M<��YXq{;X�NJ"��W�49��� �(N�e���:���;�x��3�@4�DG�)))PQ7bư�8��W #R��LӪ���)`�H��x�:  �9�v�ETHi	�f7��"pBP�>[Dbb�Z�(p+��^����n��C~&{�B�e��(��X�u���ֆ���G�eݞ.d���Zj�flm�����o��;�:��<	%�
�8d�2�j��X��.�w���^np�'��{&9��U0������48��D[�I���mA��3�Z��Lঋ��8W2HI���#sK��wE�ui9��d���&�,�z" ˡ���	����gp�P\�N9ڟ% �n��D�5��?��¾}C�X���M��z�W�r�Mu-��o�KSKB""�;��x6x�TZ��m�P�����`�E�@�˛`W>��8y���-9++���`�����1$q6���g�Y�䟞�r4z�������SF6�K>?���,�nq���@E�ޟ&%JWc� ,�#��&�v0�K\>��N;66�����]C$�j�&���i$m%i�ݲ��������*'x��ꇛ�FeXޡِ�)������ >����$��\�j����e�+���ޫ�'�ƾR����&JL_����9���(o���YEY[or"���Pת\͊��Py��ݑ��;;feu��cy�9�㿯v��C���&
JYm����KPcd��.g�l�lll@���N9[���s���������DMI����� ����@�����~���pf��p�i2��]������f~LʂU�p���V��We���҆�ْ/:é�R��
��59��T���a�;��L �߇���F�.�����4��L��C�	*����K)�v���G$���"30HKs�X�C�*���r��s�6kP0?�Ĵ˽��U��b������²a�|X���fw�V�Μ��AfnRNlllz����WnwW,$BLθ����0���O2���*�y]��C��$A@�e���v9L�b��z_����Y:ZC]=�C���= �%S�
���u�O��?�y	�ǘ��F:כ���H��[T�?P1Jx�2FIV��V�)/�s�gG�!��Y����b(_�{��t��"�X�]��e�Z#19CzV�� �FF��W�5��w=J/�$%%?��,�U�x��-����Ft���J�i9�f�b ����"i�r{^4����#��jgx�UQ? �7 ��X�kjj�*ʈ	��!��OO��&�����"�|R7����*�����5�>77���J�)�e{�ePu��b���|Sy��o���i�+ȅ�j/���KJKi]�>@��8]�鮬��$ �㶶6�
�#��Q���_��e�}����;L��A6�b|K!��cF�j�YoC9���t�:,u��/ǅ��88]��&&��B��ʊ?uL�4��i.C<��,��V�����bZ�r8�$�W0��#���kS������S�^�I���d>�=��7o�Cu��ye�1B;�m��V���b�ק��ӄ%$ v}��*�i���TH�o�W+>���L�)6���''gIU�D8>t����C�*ʬ>;]h>�����A5O���W[���D���i=b��Ϸ��};H���U�
�
T�����C>�f���T�4�.���W&w��g�LW�+wu���i�&��=괙$���'&@��		�.���\]�w���1����	\R����ڗ,�8�	/����t��u���vV>s�M�G���n$&q!��Mc�1�����Dw2a �����$:~t:>v�i�$����;,$��謙����B���=oW�2-����l2o�h"���g��3z��?&CP� �a!_����i�/10|Ǚ:<i��ĩ0W��må����v=&c�k�< ��:� "".3Q����b���7��b��jm}=�(d�����k�D?��$�c�u�761?:��t�d^,�N��j�,II��պ�,���~)�ȇ����Z����^]W������bkg�fR��}w���3Z�c���QJ�z���vQ.3��i[�9��&�vsR6��4xa�;;��=��j�e�Ck�~[ �: �˱t�g|�:5�:_�5�Y�d��Gb����+��/��o1r��d��oə�"}�T�����{�BGb��\)����i{�8�������%.ƃIy��r,ЮQ
���,$Dr@P �9�A�e��8��\P��7_�3_��.'����I'�n����{�)w���i�|޷���X"�#��K L[E
x�)��>�ZB=2f�B-����`k�X��)@d_�7����>f�[L��<���~@w�ƕi>�0hG��i��HT�x���}1����/p�2Y쿋GU}֥]���n����J��27)%$휄�(�n8	�� ��k��/ǳhmx���lҥ��O
mCs[E��`���7Z���%���\���1��0�<;�*W/���VCo0Uh���*f&&貚��k�RQ�X�������x������.//����[{6Un�	UU�4���R��d?M���鬤����|w���X[���"�|�H��[�y#ɹ�qSR��������N
��th>l|4ԃ�yo����t������PE�*0X�}�X�P�C���D���C�q=(����o�z��:99)������[s$u���w}}�Za^�6�Y�������+|)c�j�5�����_��D����).빷���7w�y|�9>'a��+.�Y:�o��_����uN�@��GL<	�U�3��e���\�D�~Q4��������񗆆a�g^
�����EQ*�����e�/�0lk���Ps)��2��p��}	���Lb���1yxxj�g��r�p�˼A���z�'�j�Y����qu��}���J��'��?F���~YY�P͗k�x�����2�������>PB�g;������������&���v'��&*��t0���I��}t�{�V ���	H �)���09%�H��$�w?1]re����4��̷�� s�]�HK�a��D"�e��	��f�C��U��p$�Q���KoZp�܅����K:}��<3��N�SEE�=� �W�q�},����@����'j"#�,V%��]?#��Ѭ�u���W,L8�Rt*LK��*ڀ$������kQh	$��B���E�s 6����z6�l>����l	�0�SD��-ƛ�� 8k�n5�����e�����j��<zw�z ��,o�P�R��K�;SAo����j �Lys���"Z���T�.N����j�f�@�W������X�B$�2�a4�Ȼc5���ʱ���(�����s�������y��v��|������E�~�)��.����w�lN�Hߢo��-�͒����퀱1�F���~9��w��� ^Ѯw}	�"�����{{w����/����魵�!����̌�ᐱ�Ǣ�]SHk]�oζ���!
FDE5h��.y4���t��	|ܾ϶ꜭ�P7=>�YZY�m⏋F���rs��ݵc��:�}~s@�k,�N��@R̢��ӻO�(��M\���:����Z'�թ���嵵v�N����ҟ?�	�|<)���E�~Y��ݢ�����{���]Dϣq��L/z+&z�_G�X�J�Ä� �K#��d��6��͹����	�;�Z��
T�
���;}�lE��������*H|:_�4��B-�)�&'|���*�;n�Z�m�T��<76��j��������T�||/b߽{G�� �����$ /b 4+�\xxy��~��B��N�e����X��5�G p0Q6�R#���V���"bm]4á��3\a�-�Q�T'
l�|u9 I��������cÝ�ԶԳ;K)�v�Z݌]~�!�d(��_����!��˥}WW���Z� >��0a5[� "��i�u���4�)�nJy_@�����ߜ��۳�좀`&(9Y�f�����.]D2ਧ!w��C]6�/%�ˤ�_�����5�hy�T�Nಌ��d��'�
���%�2���z x���#,��q`h(�ܿ�jɊ�%ӌ�8���#�<M
� �@D�M�oc'�8S��j2�쬃E�〴P���	X�}F��,&
�l���l/�Yj�%
 �@K%�3�f���S�G�ff=շ�-��9Hc���՘e9�,�l΄�eϖ����2-e1�O���g@ޱ8�C^
�T���IIa����HKf)S��������P���'HA���t�RTӈ�BJA�Ei���y�%>�9Ԥ+�8J�"��&�I���h�m�j����h�jj�7-�pe���x��z>������{�'�/���a�ԍ>�s�ä�]��{���b�x��d0�֥ި�g��%�&E.�3��V�*���j����;���/hKQS��Z�y�t饠c􅷢��u�Lm�&H���Yf�:����A9�)0Ҝ���%i\��zVe=�R�.�y.���L/��akÝ��f���~�V�zWG�v��/%ĹX�1L�y*m���;�B3�9��3���m3�S4���K`&�t�2ޅ.mm�8K��7���؛Ό���v	4��	D;Q��C�PI.SΤ��@�,zu]s�W�-��R��6�����+��3�Bm=�����ܞWo��?k���99u�t���.��չ�E�����[>8@���G�200�[�ׄ����q�Pi9�:E3�Ӄ(���JD~�B�c%�~C^�@��1�jdD�� ��H �d`�ą]�����1o�TSЎ��7KS�J��ѧ5��.�[�猹�ut��D���Ù�|G��2�.�^|�pV�r��/v]�Z��>Х�Ro���.xa��p%3���$��C�K�]�7�{^���5�ڴ��Rb����Uu}�:W�P��}��x���g{&bjJ���U
0i����-����38��N�Ȁ�!�����ѯm�T� ��z���Z��~N��#&.i�����]�t�JA��e&C�@B�ry �<��L�d5j�w�����2>��ӕd�Ks���?ee,�a��m�[�_� ���i���k~P"{b>n;*��������K�A��ۨ7F:k�/O�z �il�`|�~q��&H�lF	9]m��8�⼾к�����p�y�ꄜ9��_���# ��yCu������_s�]�<EC/�?*��IQ� �
�]���W�����������bR߈��)H8HC=�a����z��654�%  �������<==ˌ�8�ٟE���O��s�� ��q��.MQ���S�n=hǬ��C�**��DA����`��c���]4}h�~i飮\gyl���ǽ�RXXx�1%G�C.�;bA��
Y�+K������r��,c��k����D������(U����Js9f�kq��cE:ZV��P���; ,O�[q����VK=.=��%ۑ��#��B_�vm���k�V"�z�$<��,@.�㿱r,�<<,����W�i? =t����vyx���\5>�5�3n�r�
�[�ͬ��Fi�;TM���<ejhٗ����h�����(��s�ߪŅ
�U�\٬f���Vр� �;r�Y#ۓ5)F�K���_>G���j�{c���h���R�m��Et�a������]�>im�" =������M���}m5���Z�-��<�6#Հ��~U]\L8���:��_pşl������ij�3�������̸w������͠�ry]A�Ͻ�\�m@�P�Doc�� &h�YQ�3�(xS��"�V _��u�t"�p���d����x0����9�� ��:�烂���y>)�l	����vee�/��Ǒ�t��%.��W���g[�D�\y���$�`���Ǳ���L�PPQ&�@' ���$ ܢٲ�R�痈6@�oq����4�pp�M�TZ�BB$���IŔo���p���Nn�=��)�}礽�S@����>s�aM���W��nci�\�	U�p[#�a(g.u�Q�"T���-������t)��DvL;�D��aSW"�M;�;j�)(wC d% ���lllӅz�N����3@+#A�*++��}21!gfF���s�9���� [���[���niF�=BY1������	^��ED	\6t~C�~�\on����K����װ�W{I����B��7S}���f*�BU5[P���cb`$X�؎O�e��`���⦳�'P�E�Wid��5r��lF쑪l�L=Q����Pmx�!uhb�˖p�����[M�t�t#��$��ˡ����0P��gY�Չ��<���)X=(j=X��g\𠠓d#���Z���Z(P���d�s�;���^c������=��xW4 B�fg���JJЍ���������>}
-2qso�ɚ�ѦxW��6rtZ3FJC�'�^�@"�(��D�nvv,�X����j�#�h����Z��(���+�!IɏD..���?~~���ٛ�L��0M�R:�u�P�ds��Ğ�F�I��;))�V�<�g��jϔ�\�U^>D�&rj��p�-�}�Ol��V�q�&664}�����
Ssv�,�kzXH�OH�p;�����븕v�~	��֑���0��twWr���,v+bsM>z{��uW�{/�۔b�K2uoL�o�Z�
�R5�������A����8P���	[q�ZJ9�'�����!�vh�����o��h�5Y,s�a$�	>}���7h�wt� ���Y^R��4��0�&��iii�����z�ݼζ�C�Q�|ɱae� .>�S���O`��\*�_�1r`�6�=�F���<��0��R�C�ݯ4d�����8�m]8��Kj?��Q,[[�#%co����7����c�Uǻ,�g:�p_��1���A�����LMI�/M����au�*�q!����z�� ��\v:z�^�O��ǆ�\L*�����@Ͱ��|�UX���f�
I�F���I���Np��T�}�p$.���F������r(3bMJ��'֍1�T����y!#3'ɩ@d^1D��}}s�^7o`�V�*b���z5�bS1�ޠ������a��9�����\�a#���ɓ'�����B�c��O
=���888�M�k�@�����4�h��ZK� X&�T' %�0��!22&��Eʳ�c�6���3
�j�ʢ�	���Od �1ne����$�T���YJ	��w��nU��%���v�.����,���t^��韕6�ՠL��c�(�
��5y- �|Zq��I���� �+�^������������s�2�F���s��7�BBB�]�IpI
�LW\��Q���*��%����ն)���2���#�'J#|bjdb��m�O�(Y�eeeUWHL���ɔ:��BqID\>���S!�K�N��	�Ya��I;��.�$�C�<��d�9}�L�o)�6��`���5� �2��:^�� ��5s{������PCB�R8h��z�{p?����l<��c����ӳq1�v��񀲩d-��QQʊ��̘���+�d |�;8���mk��%��.�Ͻ�;r30(��q�FK�ct��yE=QE��2�?^����)^ww��'�t��P�ж}K�>�^c;u�g��L�wr��(��V�b����L�
������Ѕ����`��yټ�TR���VLA�����U�))-�D����cP�0�K�����7N��J�Ummq�v�|���z/�(��~�vTX�bC�q'�f��v�z�6堪*.��YQ�m�����Q/��\� �(*?�_�2�r�j�B�Û]j|ɕ�_��!դp:0?]���o��!�L��L�mpd���Pd�=���&��K�X�kY��>,�U���CoE�S��"�*�k"����-���	R���hEDEI�Kr����]ϛ�������[���'��p���!;�����!8M��]Ʒ�,���,�FF�;����̞��X�d�A tE�$/R��rڭ��)Y?��}57����*e�l^`���F׸W�B���(�`E�Sc�حB�R�|�~����p��iwb��p�T�ɡ�C�_b��*VWG��~~PGeB>�05L���E2��y��y�Rƙ�%���"��n�K��Q�Aʹ��>'��7YYY��T�rm��b���Z��5���L�Λl�<�;;���紞˭\aJ��$�~�kcc�e7i�]��`�KL��*��KL$��ED�fh>^�r�gm�f�j(��L�kށ3؇���������M�ɹOɬ�4��*M��`�š�P���!�`O�U'Gw�,@���7�0E�D^/�=��� �}oc�|{��|������%����� �{^�.�K�;N�۔Ę� �c�}!H�_}����U����w>��LD��,����qX`?��=W�[ɒ)��/�T�g��r<r*i�C���<��{�)Dͦ�p2�G�����YIkR����o9�V�c�6_$k-��"F��i�ʀ(�t�������? �\��*JJ���A� v���Z&'q ���� ˈ�eM�ƭ��	�7�
��������(�>��b��!DDD�d*��w���\���0I����z���/�Jf_ ��T�sr�L���ʙ=a�r�Z;�K��� Б�*��wZ�ri9�r�m~��ٹ*0U��z!����N"�r �:���w;E*�mz��thm �̝���U���:��J;"�f9��;1�g@m<�U��sC�mmh�Y[[{Mt���o���b��ބ!"���xC�^mDsȞY<j���+�����w�1�6ӫ�y*�eT�&T{ʯ9H��E�j������� st�|Q:�m�}z@����X�����`N#���l�-_�`h�qiyy;x�,a�]>�.�i �c��V�ۂ$ee}��O�]�9V�Kŋ�Ǵ�Hf)	/�KS�����u�	M_�˧%�2�p
�DI_cIS�D���b��$5�R�R� H��4��>W9'�t7((�!ewm��h���~����ga��v)�}������Nz��j��i���=
��̜]>4O���!آR�K�{M{I�*]}ڜ�����Tb�G�!��
B�-sfb�8!!!t������K��/��w�w������'4x��WQ�������p�	�MZ�*}.>i��h[�=
�3D;��dx+���|Y$h�T�F�)�8В�����	LNN6�N�Eh����~�3h���ZSg8�T�������k�<�@�g{c������',��NO���bڅ!��]���jn��q�̭�uC�.�,��9m�߮Y�$HcƋi�t����Ng��������	�v��u���B3U6�͗IyGA��87/�}�-�`����0[3�P[�d���"�ۚ�ŗ�[��`*���5s�0�k0��8����ba5И^��>ŕ�'��oF�Ō��7d�]}���j�٧��.¡��ގ�ܦ>�섀Y�:U
����훝�֟(�H�r;����r�}�ߤ���sZ$l�PR����1���)!�h�a�R�7<<<I��<�64�4K)����ؔ����^�}wG��mL�\�v��|3J�ǩ������'0�S%�P{X؋�O���>�'P1-���_*VWW��Ce���ݿ�h���9��Qc ��N-���f}��B���We8�)R�c�Յ>�������f��N���e	"E98$ �����Xp���(y�����A1�X����X���~�ݝgr���v�o��Ţ��|��/�[�P%�BJݖ�q�Y�����zS#	 ��ά,-?��p3��-.,H7�:���xe�p�	F�6��,��X�"�;[�f���-,�x��1��F{���(<�?�;ut��TWR�CO�@G+�>=�>�\�R;���УZ�@DB�?�g����fz$����{��@���k��!��
�
��������{ѠRe��7S��u��z�����F��3�����a�������݂B�g�Cr/B����.��4�+�'gf����T�AÞy�-����ڸ]�r��5���,F�%O���-=������D����3���^�T��ZM�&&f�٨x����ι������5#[mb��X�VG�_h�I���Ko6�ظ�r�������:�������颅1�.i��CZI��i��TJZ:�����N��s|����sfv�5���FFYY+��Q�[� m���&m��g��E�0��V�����A	k��Jԟ:��;�g������=�Gg�hE���7Gm�H]�� Wyä������\*�'O�wW�4�Do�$��\T323m�H�o�ɕ�V�����$
�h:<�,�6>������2��6��A�HnRQ�|.�����on���yT�Л^���Tޤ�Gb6��s����X������_s/�:�|2� �U1Acs�  �I��po/�|���ߴ�mO�����Q�RQL�Wf蹊��x�8rX�J��F"�û)�ˇ�17Z66L222�y���]����ҿ�~zFm⤴RR���Ls�*b����a�]&�n)��i}ec�l�f������0&��E���3Ts�]��+��q���X��%m����2_M�Օ�T[�"�� z
G\#ټ��s�@����*�;
�����R~95x�'��RN @["8\3��w ���O>jsR�n���۷x�o;����
c��۸).Ab���Wv�1Ȳ_i�vOv�s��uh��i��K֤�ux��ۻ�b�=MS�Z/ֻ(졔j�9**�7�%�5����&��|�����Ny�]��X������E�k�-�gʸ/�"��H���ڏ�P@K�� ~6k��N�ɱ��V���z�iT��ܫ��(�������<>��������j9���¨h���A����z�_&��.aB��E�QI����T���ߪ���4bk8�w9�~�aξ
buK|⺫���^Vޜ�!>8�zϪ��z����U@�H����4�����7Q[C)v�s�
�Ǥ����q}|��riS�{����i�Z;99�!l�*���˵�ʞ�V��<��r�V�PV��e�M(� �D�����bmѰ9y��g���i��y��eH@���'�|��?���S�H�lmG���Ax�>>x���������qx"
����&�l�T��a��eh��V]e3?5;u�{�f	�E.� *���h��1QI��t.���1���^�,AT)�O�PEU�{?��L�=��%����=��+a�"qŽ�ݏ�{�r��%�8���{a9Ӣ��C1� `	�(I���}&����h"E�Zʥq���ʢ�E:J�mr��`jf��9�=Qf���!iyņ�̧/�ZZ����3nhcc<��׀��EB�p�b�c`���2M7%0����\T���f�ʋ&-�u��^nn�'�X�"x�y�f�
3��E�6=I�9��H�LV#!�g5hG\T�<�˷�|g��P�(�Pf���-�W3���3]s��m��]<2���/���)3n���6���#44f6q���(J::���d��K�H�FIǤ��+�O����7�����`�+�vI/��GY��)9��Q\�������{��Ë����W���r%""�wVV�#)g��ܑxn�oW����}<��m�������G��J�2���kgB���#CBt}���UG���N�\[]Ͻ�/J"n��Jh����H�A�=9~]�O`NNO1���K�����㔒�i�$�0{��	
j8���Y�i]{V��m,�M�c2����Z��A&�l��S&&&p���[�_9�L��Ņ7��ȈG�
�#�Q?I*��\��y���xN�����,�UQj�$`��O`jjj�C�nT�թ���0̢`�	,L���NNN>=l�=�� ������k�xdr�T�n��_������bT)�l_,ZM��u*�^�����Q�q��w�?W���ؑ�����3��؍�ȣԢ9y�6TͧY L#I6��fѶʋ_\\X;8(ٿ����ܞ�J�%ڑ�TSU���Ԩ��d�`Qb�\���]��b�o�,�j���艇@n-��舤��@��/�',,��<>�E1$�����Q�i"ߕ�l��9��}�	���Z
B�PF��Ǐ�ħPoQ�����.��edD��c����
�_`���R�')̦�ڜ�P!�0eX
����z����v!��Г#6������``�k,ë��䉀u1���ln��;�݆�t��x����	֤DHFy7���Ϫ�.���.��	��פ��f=���H�8�wy�������������5��[�
��Q��	ѡ�<� ZM.m�eҋ��Q5k�UTT�ߵ-Ԏ����s��� �x��r�ʢn�\~�^Dpr8��1�'�,U(VK|�m��q#T3yw�:u���_�UG���W�Sݧ�x]3���%Ja��
�{�t"ɥtH�<o��3�ÅU���q�<�xD��M�z2�O�]�{�\�:.���me�f�磃 ��e�A���3T�ҿ����j�X�R��=�i��"�q �g���K��92�s=�n������ 5V�d%7����=J���]C���o9���e�?o}/�v@�%�.�rE!&/ҞT�l$���FF�����D�㡜HL�L����-��PP1�A/RVM���x e7���\�xݧ��ߨ�V>HH4��ߜ[$ܺ:9L{�������2_�����;k̉�_�������@3e�.�1�֤7H�<\RqyI�����QI���ٙg�ݴ���H���{n��֧ ,[��ޗ����n���;;ӊ�eGR�+S� !QQnn<��Å:@�^,�x �����v��|�A쒨�Zϣ���}�e�gM���H���3���J�O8ah���+ߧ�XXX�g^�5�'|�
~�WB�j:1�3R[���l�C���nh����RV
A�h�Z��%8�t��ݩ�|���ΗR	�r ,m�FC/��)}��5vG����2�N����ҿ�o��`4��x.D����5,Y$���8q		Hx��_4���ce1�	�R������{�C�| ��#�C��Q�-��n���F�?R���v��4���a[6Ϫ��dͫh��|oMC�v������Nz�͠%��O�nK`7=������C~ɟ��5�UA2u�6�	�VO��m�G^�N��Ν<880�W�<3."�۰e�s�_�U� ��ϯ�,wg)7���vsOOn����f Ү�QTgDJF��;Y�=��J����6Rcg�)���@B�(L�'F�Df�����:�S�u	��t�DL��~��%������$K�RK^!m����;6�%�}�0��ѡ�Ⓓ�7L&�=��ر�Ĭ"�l���䵰�|L�4K)n�%�_�~�{l#�%�8���D��?&�u�@���:M�t��R�d���Z�۟���^-=>P(�R>{��0	V�w}.t�Y�>�_n(6P}�䳞��֜y� 9�m��(_�����W|$�Ut�J�71))aMͤr��b�go�ȭܒ���֭o��������֕��fբƾ��yZ>|M���u�����k.�=|�h\��o���kF)�׃&V*����բ�^7Fl_�h�D�î��=��l��k��m�g�췇?�&��ʃ�Y�;��3���˪S;�@wA6k����m$1�r�����.��|A�i����[��W��K����a�1�2���'�:3����$�OpI*�M�xs�5��9�����s��������zSAĤ�3|��?X^�Ą������H�K>*��hߒd����[�e�h���L /�XJM���Jo�\��ֵ��ϯ~��6We�"��*�U���t��ղ�땚��S,z�W�;;��A.� �B=++dHf��cS����\S�_5O-oii J���f�x`q���p����[������g���U�0Mrg榦�,�ȑ���a���+����7f��?>���N��#⑗�����绠�7v��y�z�C���I���u��E,r�v���ܭ:�L�Ï�K^�pb���2[M⬭�]��n@���H�q"�P8�:_:D#�j�+���Z�]<=]�7,r��_���j�%���́D����h�nt��ƶ>��s򽈥q�Su���uk�.!t�d��eoLw��+�Qn�Oa��UƂ���>99�� +���9��A|�		i{43h��C��2_���2?[z��eD)����a�祿J�<�vz����:�h(���?E7+��! !=�����������v�������!F�>�c9�8,FG��M��P}1T�����)��y��d���Ț?����L�0B��2��"q"v�7g��/���#Iq�:5�,��$Hz��~���Xn�Nrc�O;�*�n�WZ��)�B@D����Փk�z�h���4b��)-%�\�)�+��9+[*V�Ϟ����� ;�� ���s����������J��=慎OX�Ԋ�~��$f�;�Q���@X}��)/��GHvʓRS	*�u|��U�5O��h]�"��Z���w�����4y{����J�FHHXu���ݘSV:�ړ;�j�2Gk>�=A����������55�B��⊄��J��o�������Mm
�l؍W�H���j^��G]h#���b���'&㿓������ۼ�9�$�����P{m?���"}�@ �����Ƈj)*�@���V��5]�1��'r�/�� �U]e:==��ow�v��w���{Wg��|F����x�j[[��B$�,48`��N��x^��p�xz8��$������F_�g�Y��fYm�P ��%$�Eðf7ů�bi6Yu�ذ4w�����ށ}��2�{�K�wvZ�-*�����	�۝U
�c��M�� �L!>��x�=B@�n�y��WW��+�f;caūѕ���z��O����4�zEBp�ز*+�w�s�'4���vt�KNvĘ�	��*PT�Դ�P�i�����t,��W/7y���bZ�{r-�va0�3���]P`YA�E@_��q8hx0��ʉw@XXW$E+���ԙ�jJR,�&�i�0���t�<ckA` �ɼbҽ��vT�ݑ���ڠ����)|t�8'/4F��@��qL�{P�s�T��I՛�� Ѱ���
I�z�٦�x/?���^��WT+�T���L$��HyoC�Όw{y����|w��8���m��z�so�
ą��z����B���f�J"�Z���q/�n��%=T#j�FI5WKV��i9'4��j	��W �Bzzz�� n�ViEEHI׍���M�+-ް��Xy�� dɇ��L��{��F�׋��	�p�����/5z@G�HJ�����<��/��Ȅ�J***��\�+�_�Q��V�W���v!] :�wF=;�K�WV��x=�WUm�+ ���V�lp��
#��|���8�)�}us���Ҡ��ꏣ#�$~/?RR�ԯ��6�M!�4?>\��@b�%����_j[5�eR������U4r��)�j{zz
 k7�=�xy������7V��biaJі��-À�'!��LT,�����'Gg�����M`'F}����`���.����gMW��9k��~�X�k�[��M���ueF�q4E�.�Rn:����^��Y�!?�,�u����(,�Ra�qN �����G̼\�lk �%`6ǫ����^Uq���都ܞ.I،�;���-/����6���{�� `��
[sS����8!Иm����\�\tv�mEC-T 9Y���`����-���=�o/6������]�� X-''�n٣�(8�_�p��#٤���:S�{r:��w95����#���������Y@Z����7o~�g�����b�%�Ӯ][n}g'�������=�؀�� p�ˠ��|e;=Yi9�|p@�2>�i�O��e�K&��p;�]�X5\�������2<9YXJ�I|I:*�*��7�������~-U�W ���8U(R~3]U�G��OyT[P��^���9<�wFv�?[��b�l-'�~�:�H釳[�2�a���m���_4cr2�_�ϔ��݂��7<r�$7�SH}�7��d�k��~���u����|���#ނ�j��|TP���ޜ�`15:* R!�˔����v��HMB ���� �dff�q9P���cbyg��r����y�����U{� �G������H���w����kV@�x��ԉ��붧����Y�BL�t峳�/�iB����ҩs�sܟ%S.%���`ϒ��b<�#�$��e���r������[����I�N�iiio��4��B�?����홖{����������t���������PCk�������z����������&&ffŸ�|������:��3�=��F(�����¢�g���K/�~�e9��n�eA��tQd��$�l�j�Y��pP��a��<+V0y+DJ�L��q�E�`p�������`}����0T���w$���4�\�� �_`��H���=���*	4� #;����
*y3%��SIel�pG{�s��=%��� ��n�4+�c�h��д�?��C�U�v��ќ�˾$f�%��Y�������=�e#���.����|w� �����0W�P�b��R�_>�M�FaL���ҽ���7^^^&�E��5p�$���~��C-Ԫ�A\$K��d[C)�!z��_�)�?���?�(�+���V(My��`�	i�A�P�1͚9���[H�0�Z��������0k6�1�kJbs?��1��caF���uĐ�0�>�T����I��|5�&@j�嬘�y;���(1xN�����E��Q���n>Ƥ�ݹ��{&ɥ̔����DF^ej͘�d�j�1;�|HK���ڟ0�\�Ol@I��,^}tS>Td�v5E
�W���K�i�* ��ќ�u@��f+-��.zONO���p��b���ŀ�)�{\�͘�eIE{���[_�5>���`�f���$����h��
4�R������d�ܴ�^�X��I��`n���v����� �
{w1g�oz:���^Ol\eYY�J�?NJI�aO��#��wO�����>&�[.�� r}��,���x�Zm�:,t�V��\c|Ɯ��i��B��%�C:h�I�Q�ǲ�u\� Eo��$�/a��\%����H�,����kH"��c5Re�g��Oѧ�*M�Ds@�R���&����j�g� ����F��h��6��ϟ?�:�����)o�Xܭ���	6_��v�H[�E(��W����ׄ������a�����5v8��x��y�._��GW~���c�ohX�ަ,���r�m���5�0 a5z�`�$�y�>2�!}�;�.~E����@�ۡϴ8Zn�%m��TPA]ZZ�6%�oc�?H2��h{u�Ġ��?ʍ6�wp�/,�P+�3Պt��ŞZ�Pfm-����5��m�����V�2ʰ��A�$"�h3ssᐑ�(�m6��O��8��R����y_�OVrsu]��[J:��ҥ�|��<%H�z��\�?�-H������p��>��+aa�GKZj��d^7�	U�ut� �.��`Oa2�T������a�����G���ŋ�� ��O].��p�����;Fqu{�67�x8�v�=��5sҰ���]4�j©���X�ʧ���H^��
ⅴ� 
� ��?�_��$#�[b���w=+ '7�G�f�<�98S�W펳����������qx�4��� q��b����y�)+�Q��+��;v�K��v�\NNU�-OW�Z��l��#V+�K�S�Sx����o�`� ��SH�403�HC����^��hX����?��P"~m�L��̜�W
�� c~���M 9k�]lG'�(M<F]�_�gg�WWW?L2Y���k쌡�}Css�`��߾}s��a��6��'MO���)���b@c� ��`����=G�� �w/y'��	MJ�bF�ۙȇ�Ym���G��vss�0����Jwdy�џ�8Cc��hT
uﮎ���������j=�_.���@���7>��؟}냒6�p�E$�৩�%\h��t�'�fԏ��J��"l��.m�-� �I�����y=k�=���W.aM74�###՞���ᇲ��4�B�n������R`����X��u�xт�f��#�IGu�[��i�����yl�[��k�Z{�t&`�E'����b���Â��j���5��v8Ccc�������f�3#�6��Sq��_�x͛Y
MG�2q.���M�:�(�����Dk��#"�#p鎤	�����(�� �q!��ofp�_PB�9Wn�̰����?�̯��D��gW��u'y�����U�G8�#�aڹ��u�;;���'@Eꟓpqq�3���D�9/�f������فg``(�Z�~O<D��d���RW���ݲ���v�?�B
�L>7�d��/CӱG�eɄюO
�}�n����yۤ�
& �'RK�Cjz����J�_`�Z�:�  Co���؊||��y+W"�"�u��9(+�c..�W��z����l k�N��ƪ�DkM���g���/�e
:�~	����E�Ǟ�"���6!c�����Ǧ��(]��%������B�C��qO���)�r��HGGN��P�����z�٪G�c~���oQ__�,��ɺX��T<�{%EE�|tt�VK���NzO����`-±cx��o��[�? ؁q4����s�1xhbv�ӡOQV^/Ā��O��N� 1�H��R�/��d����V�D}U)�~l��pp`c57l�\������1�a��	��@¦uEN&è���c,[F7��`��4�z�;��]�q��5s��(�*�oc)k�����s����{&����c�Bg���`�*��	��X��/�����+@#e �����_X`��]$����V(�r���(�EM�:�z�ڷ�� �[C�W�UK�8�/|}}������a�A'!F���.��j�s�������cv��*/Mi[��0�5� aA~��کF��;]i�u�9�me����'�,�9���Fs`�&���o�fM��7����۳5��)3��-�W}�m�L�r���Δ��s;b�&ɿN�b��G�UdU�Oc�|+m��5�<���$g�!^�	`�����0"������2�[A0��w�
9p���s"^~�&��*��j	Έ}�4��O]N֭Ȑە~��R��|U2Y!@�?���������tu}�ܽ{@�}�05U�b��v����1�&=6 l������ ���><R#	�e�����j���M`��9s���@�G�*�.��UUUU�&�͖IQ����,�ym��~���[����s[ ��p���ELI�jqq`D=�.%��5N��B�~������RD�����G��#t�=���H79C�337ăr�;���l!�RM�lb�}@ob���
��݄�[xu�a�1�5�,U�����5�����4 ��؟���������;�#sy� <Y�r����.���{S��+�{o�ޅ�r!FK��󁅤ɲ�̫�!�� �V����}�u��x0)������� ���s��}x(��.z")HHI������
�CG���$N(���h����7���$�y�G��\��[��"�0�����q�����|��//�������)��F��EBV�:;E�<zE����kOw�:�>?�a����0��7��>��.��$%z���d��x��eϏ�?�R6��1.�F��^��Վ��J��ͳ���~,ϫ��≉�4Ӆ�vYȯ��i�����p���p�V<���������H�gzM�7Rr���^*k*���$��_��w��s��/E�r~�(o쬛X�ɄH%�/���J�s�)^P;��d���a㺄�s��ɉ/|H�q����a]I�U^���l/5�+�Q�\����w�� Y����;�N�ui��ݻw�C*�:Q3�\�L,fJ}G�bw>�g��́ ��;�s�f+����ʆS��������q������?l�N���9 �ed�]�؆��� ��|��G܏4�C[����..�i���ip}��s:,��w�)��UR����	�>�6��igG���{�JWM f��g��30DB~23���`o�
�"WC"��ay	L�a5�r_J������揎2?'hx���Ф<�[ڼ
M02!�j:ȹ��5Pk��\�*���{�ʞA��ܲ^�������o�绹knA^�X�A):�e:[���s��4���a�70��F���dIƷ��
��e����E���G �G=ܜ��:1�'������udI%.��y����f^��ͪP���Ma,���G_�n�q����>���%�¬��:�.�إOb"�d��E�+���=&&�j�],��/tŖ���K
J��,`!���>(��O!q����s��w0�bg�\*����e����Ήh���ٛ����)&J���?j��ˤ�>6r����[�D�T{ݟc�0�&�H�qc�v�{�C +C���ћw�������W�!ɔq��49�5wWG�bfi�b[y{�%Zꖖ��9@���u������Î�m$>C `-ol��ORz�WG��޶����:�d�ZT����S�@�}8��Ǵ��+��^��{|l,,h�'p�NH�PC�U��v[��h��� ����ܦU�:#�C8 G��n p4]�a|�ߕ��f�����}2+frR�����H�����֜�ܚ��Ԁ$�=Aߥ6�g{����\\bb�|��`�M��3�`��lkT�MP��^�|	]����؟� D���(���w[d�&�{����ყ��[�#��u{���<X���+�P_*4J
�����1�@{tt�/�1�-�'��g�qԙp�`��%n{ߢ���/Ui�.�&R�WO./�9�j�����[Z��M����A,��}?�Zmu+���CY��S�`^�h�j���&4$� �������"���`Lk���Eݙw�� v�����\����A(Ā-#ud����|bNe�?� ��Ja,yP������"�B�˅/3�--�2o�h��;�Ud�������D�hL2x{h�J�H6���7S�B��.��;���E@�g�LΓ��e�*��9�O�V5K�Q����K.�n����i�pJ&ޔ�>̮�����������^:Ж��[&�iFRr�^Km��|z�:�ƈʻ�� t&����<nW�|ޛ.�si��^����.��W����5�]"��X�a�)M\W��E��	������B��擯+++��T߽����[���T�6�"0K�o- �tYD�[RQ�QwU@TA�W
��q)@H�D߷��Lr�[Z����ҙk���ۮ輻YR�:2��X#;�/X'�2�r��q��B�~�o�~(u_�]��:�E�=� �&g%~)^�ד�i�fJg��2��J1��b����T ��\�U�.q1���K�C3���St/��2��"9��E�{��_��J6q(��� �$���.���������K�֙�򸨧�&��y�X�.]�w� ��,� F�U��L����oX����H�}{|a�5��3���R4q�̈�@Bkh��ZW��	,�%77��Bmt����8��ץ�S���P�h��"_NEF���ņHg�Śzff&������P2/1vw��s\���{U�ŵ�lF��IE�ɓ'��eYH�,6�G��?�dO,k�Ḳ�%C�~�s�&��a�jeFp/���alO�fX��9"�F��<|~�g=Vcd��l�����9��]����"�|�����S�8&��e��cS������<�]�t�	LUĀ�����}e x�����Ag��a�ru~ho�OS�VlL���YB���r����j1L�NS' �W�~_fJ_ !!�P��P>�744�1Dvx�����4E���F�1^׳�W�c��<D���617�`q����0� ���01�\j���D��I�a(((T��(U_\�ϥC.b��aÈ��ƻ�ڞ566
�Y���{]�5�x��-UAB�@͠�E;ĝ�R�%��9+��<,vd8S����2o�k\2�x�	4~�M�-���ۃ�:
S�'���>|��&����
P�o�u�t��ӓ��K{=��M�݃�o�����\��PQ%�&˟dk%��L���4�J��[���]u���'r������X�<�d��`e[�00��*�q�TY�)�z�LC��b���x�K�D_����W��y�?��ER�Pk����|��U����|�fNA)���|N������Eg����ǡ�ph�,$q$'���~v�ӠG]Q��\�t��4����4�ښ�:�a��n΢����gl��SNγ?�r� 6�)3f9 ��|���=��&�b��Y-Wv����Ѯ��*��k"����=O����"� .�\�؂������e��x�ݒp8���_蒓���_'m� ��r�^�j\��d��(`j���j.�x�8��-�0�����f��`y9�� ȶ?���r8�����Ѩ���ҙ^��{�)b��E�TKhO���t�@C�HI��^����C&	��J_�DYǏ���"KKK�*��K.?����S�aӣ����6!�t��J���B
T�����~����<�2�����Lܩ�޼^˕�f҄ﭿ�F�I����a1z���rw�(<<��r���3bj��aM"&H~����,��,22UnE=_� z5��Xi���}
���	�?�R\̈��'G�����(�~�c#q��q;ꣲ?>1�,�$K�;Kdtu�P����N�+��4�,�ײ���E2'�:�ܦ�,a�ᰒ�$f����<��������0��en� E"�j�[j7�愥��� �������ͼ�ik$Be-�&�����q2���� ���K��@�����^����˘Hh�ٹ��̠6i}W �C�F��/n�:'cV�/_��&.٭����n�<a�3A]^�؀��OBn�L
��C�Y��߿�xkݲ�B����0m���q���|� �^i����z�/��
�h��=����a"@\YY).)ɵ�ߙ�w>Z��M[��+7U�����s������&���L��X1������Jѿ4.Qu�

ʿcѪ�B�T����@E 2/�{�nJ}���f�@������ Ůj,�F#\]�E����b����������g? V}v�v}>�1�,�_�kq��ܛ�!�#��Ή���!�B�Q�nz�;hC�B�4*?���@;��\;��@0���w� O������ݾ�H�߉�
��z��*A �F�|j�TS�{����?��^;W|܋<=��6�%�ɶ�>�o���/`�U����� �٥0.A�H� 𦕍��b/��Z�<���W��IϽ��$CՂ�SF�I������z�>p���br�� ]ҽ=͕��LCjH_�j��?���ޞ�����j�:^�SV�tB�tc1i�s�HR�r��i. ^�����*��)'>L��C��E�:��vbo�NŐ�HTTT��ns�I���J�Tِ��5�*��/�_��y>�c2U��kN!����uU����������|��%�������4�S$_m����x�N1࡟hHH��m~��:^� ��r�<]�H�9F�(S�ў-��1N-NN�ѩ�7z���g�������é��ѩ.��*uOfgqو]��
0�c���x�կ�l[�]mX����%�}f���N�8�����+B?a*��Xl`�o��1�rIϗ�}���=(x2w�3����N���ӧfw��,�����h��i��F'��9�w�Ѵ�"Rq���p����7y�ȉ��d
��~��jffa!��"����8����`bW��Վ�	fGii�h���յ�����\x��Hzu�/�{`����4p�1<��ν�����,,4?�`��_�+%����qbiltT@R�N����]�@��rS��~���+����t�8~##����s��/
������(Yٟ��'4�9�6��d��Z�߇t磢0`t�������R�:������*�������q����.�퓓���."���n*��%j�  "b`��u91ܛ��<F=U����_�S/N*H���--D�|��a]G+���l�H��8�oXT���%[�(^�A���)(�[r�.�v����
�����P��"��ߒ� q�#�0�w�q���gP��*��Z����Xڴ�ò��a��G��\�ƶP�d«5�C�G�51a.z��Rį�v�'��|
	d��>�����e�Paj��^�������|�G]볪��,,�3)�G���/X`�+�Y��%��|왻La0�1�k�r�k"���^Ԅ�2t�y���b�g>�{��F�6K�-�X���o����*zz�o�I�����N��Y��j;;�'�J m�y�;·�(�U��$G�EDT�`4C��l{���;�`s?���4lx-gY!b��	~�`����2����
�c}A�1 �4<��+���M�����Q��...)h���zz�JKKu�c� I�4��_m���I ����Ժ~o�b}}�����r_�ɉ-$v�+uW=g�6������x����D��V�^u[3ʚ���������۷'�UVK" ɩ�S��*���jii$&�9<!&:��s+�0k6pBC�\�ۡ�l5�����e�-.�_��ޜ��Ѳ㦐JJJ��AN����++�X@f�:_0��t�>���V��S�дu���Ϸ��Ae���6bT��<Ag23�>��~/k�C��aYMt���m=����p�k��{�#L���.<�'���l	��ΌB����pb��a��V����q���Lxy"qI�����|{}�K��_c�������/mo�
��BY�+��l#�V��T���I#p� ��?P5�T";�$�&
�JW>�A;K	 ����������3�����:֙BJ`�������EDD�����,�@T����6�>�,� 8!a��������%�����5�iH��}�g|����n�2sp���b�)3�.���)���XV�ݯ�I��.�C'��z����2#6p���˕,�ܥ���������x�
���3���$B��Z���@d3N�ز~����BJ�2#SR[<���c�А�.���k""�F����7�-�-�L���B��:�	11�����$�m}*D*�&=��G�#璌��z�K�/H!"F]���DǞ�=
���+���JM���y�=��z�Ʉf�Ui���tWZ}��c���	Z�Ȗ�iTf��*PQUgT��rz
%�D>;::��E}�MEf�uMM��_z9Bs䙣M���V���χ!�ْ.�����>OOϣ�3��e,��A܎�é����66��\��8 $X]_���
U���_"�G鋡�$�jOȮ�~#F(��CsU)ת~�ԝC�F<ْ{}}��*i���+�l��<��V�J� ���{�~4�]ZLuw =xz�Ĕbd�^%�'^R�p�F�!2U1qa�X˾Cf� ����-��Ɋ��O���W)G-�E�ݤ�o��H�����7s�Z����|HW��+���g��ɱ�s���	��꼇nMh�j��H�?��F���P���������PU=ɨ�����v��ܸ;��p��,ԡ�kB��6��}��);�p��Y^�Փ� )?Z��"ʏ=S	��2����b�L
��^BT''288���Z����ZkOLMs@�>NRJ
�2é���5����9�[�-g�CH�����0tyY���q�a���Rc�p��N����	�J���ss���0U_ {];�cff �y�� ��|�eq����|xt�;�5�AA�11~*E�+����v��j,�����		�a���� t���C�~sw||a�`�"^�;;;ۓ�,!\��(7y��i�����u�^Z͖S�:�$���<�|xl������P @�{����=�`�����BG��K�������r�~/MM�B��P��T$��UVVZ;8X�_�ρ����R���~�����tO �~����ʁ��z'Ջ��Eb�<oY��i��K�sX+�4��*�F?�ؿ������,ғ�·ufT6��=>jfaf�k�[E�mo������.��@Я�$�.@|p�Pqp��voy�pN��$� 8�DdP�������e��������t�i?��� �yY�(-E͛���h�U��1U]L�X�66��'_ۨ��eU8�"X��$��l�M'OH�@�ҲT�  `�К�:r���"��W�χq��#4r��j�H��W���(#�.��P�m�T"��p���O��f �����O���a����:�E�796�?�����^�pn�.���^f�ܛ�LN�scc#�0��}<���g�m �6u>�&Rlb�Q��׶sS�7ѧ�3�K��s�&$�LM����`���,0c�Γ�U�O"vmk��N�����[dt�/0�ŁR����0����5�-F����ǲ�T+|$���K�`	(j�p"Æ��\�������`b*m���MjA5�h����&'�@H�;UuB����W����?c�oh�����	��`������l�.iC���_��n>
�����tдw�:_>�uW��<�BU�z��@��P?��4�ZE��}	P���q.�zz>^,�������m^!��9�-_���XMyۑ7S������ނCF-�n�UVfA�x'���BBB�w��gGIl��ǧ��/�fizZ�~wQMM�x�=�8诧��c(��t5T�+�'aҙ74$���3D��)��j�L�_ְ_׺ ���[��;��ZAw���J�`�8+�����ш�P;�2�k.�&7:ӔZrn�p���U��|{A�^a&+��?���$$$B��������uNȼ�g�ܬԃ���%��kI2ĩ�g������#K, "t ���;'C� ���V����?{XC?puu�".�Y{���+W����[C±/GFG�.��T���|+.?�����Wh���R�PjlKÄ�|Y���p�(�[i8' KPp����NQR�`�R��N�Y:�3��� ��!�ul� @k��8�4��������̔�13���&�s�����34Ե���1������^��t2w����v���*PUF��6G��O��!w�@g8�(�x��r�1�`�_[j.���t
��a]�����˅�4e����m���E��n�=���&Q.]E���C#�;==����'����[��èþ+~}.@{��?�RS�A�{Ѝ���!��+\R)3�u!"��;��^B~���_��:��YY�P�@���8�Է��HZ��d>9��������î5��Lv�؜��E���[�����;����_�V��!!!��B�&����+Q6)3�ٛB���3YG��~�M}~�o�(ǹ��z=�����c8�e�էjn�A:)\o����%;g��Tm���VPX=۰�����K������1O��H/�JQܛ-����FGEB��T^�PSC���� �D�T�znH_������
���us���%���K�MM2[)����c�*p����p�IH|<9��b`����ǲ�f��2V�U����>�ս8|��-w�NKh���Fr�z:�Wx89I���G�ku������o��2��(���@�&���>�by}wW��TS W���F��M��7?�L�^͸�-k�e����[(�XU�(==}i�,Gfk�ӫ��I>���b�r�3���U�s����K(%t辥E*z�4v`���؄�usf��roK�j����+�U#C����zK�Fu��*�x]M��"��A�����ݳ��͵�����Bc;\�%-M�x&�HΜy/�w��!'��4�o6���o ���w ��ۜW��� ��mz��WɐX�S��M*���EN��p��1�0Q}�e�aGGG��t�cbDCh4�݈1��Ʈy��k�ĉ_ƐD讎W9FFEA�;*�89q˽�z	\e�!{	^����8���(�����{*��ss��~��]!�ir��T{�DTTK�yY����5ѽ����,�u!P.�z��`���� p8�t��+��a�0�L��O"K�	7�����MAA������޽��J�Cf�{W�`�>�5���gK��Outb�T2t�Z��!��4ݨ����� ���!TlX�z�LSZ��ۤF��j�����q%ٱ,�qe*��]l��Wc}m�X/C(���E3�Ѐ�;:x�ӝ��h��K�� �@$f�v�� �|11Z�I�ϟg�`!�5�J�c������Q)�J����4t�2�.M��|A�R16���c�P/�ө1|2^^B�3��lk�W+-��`0�:�t��Ձ���W�������x��5�lW��W�Kݛ����K�g��|/I��N�-��FFF�=߿T�^0�v����M�U@F+W��i���T&mG��X�P.��u ߓ^\�[�PzC�<Ѝ��B��������,v�2����a�WC"B2?�-OLLi���2��1��LB�����`S�㠰A�r�c����"ss�v�,�9�q

��v�c�\d�ܣ?���̨9N~ޣ�~�{��֔s>|� ��L����F�WYY�����j�ɿE��Uz�X�7U,:5�S- �ٍ��_!�{�i((�)�m/J����G)���޾m�!~��M�T]?;{{`6.HHH�.���˦��E%$�lP�4ޛ5n��|A�73^ǩ[<<<�=�թ�8\p�l����NѸ�1!S�UmhXO�*0^~�O�A�Q�K����>�a�G 6A@�g����ä|3��)���`�h�o�)��zN�g�N�V<�[������ݺy^$���t �`H6չ��Ғ��b��a��A�|mFs�.����ۂ�T=I!`�d�@�\c�����a��N�^��^�!�;j��� t�.���f��۠�v�� yږ^����wų�mm��_ m���|3��T���')�[7o����tz�5����O�����N�
3��I�h�_�&��c�<�N�i.�S=�"3�5��i�������.@����7�����Ǟ��wD�B�6��#ge��ߣ��(�{d[��3SK++_������xf�IG@E\�Ssl��7��2[����_6\)����󽗋�.-8�2��AP������xL��k��wHxT�P��)Q.+��q'����0j���%�X+�kj<r�<�J2�t����V��3�����Rɺ�w��t��L���ю(�Ǣ����{�ބk�D��{�\$]!��;oM�S�fZ�'1��f���N/ǀʁ�Gy��K=�ttս�'"7yx���oQ�����wva]p��� ]�>�R��!�a��b���/��CR��+MJ}�g��|$?B�n�L��=���:&����+艚2@X�݁ف�7h����_�I�/��W_��>Z��H%?;ٻ����D��!"���am��ª���s�1�W薏p:1}���5՜���.䔗k�������N �z+���r�-���!�{@�����F��Q��t#vf�:.�Ļ�{���9���D|����v&���o1- ���ЛV̪��[�l�;ly��^��,-��ފg�k9S\
)sf���Yo��D&}�4���g���U�	yb?��n���pLxd�&K}�4���)�gw[YRG�P��߰7�͖��&FN͸�Ƃw��ry�?�{1Ńת��ΟѲ�U豙N�����衎��W�5g�_�����s)�X�ϕ�z!��'�~�W��)}���cR}0Bb[?*>^Ǩ��8=��2�w��:.;[ú�#g�N�P��i��rr�5)@P���,��V���&b�a�2�(��De�F=���Ī��"	����#��1׾U�/�+��!�l�;6@26��������V|��<CEi���V����v��2eӾl�x����#%f�N愥����1�ә^�Za���/�7��*��E�=�2^�Z�G�,�2Ud���sZ�,����0ȹH	L���ܱ�W1��F)&���z�N��,l��UT�wJ\(��.�>��\M�el���PӫQ����޷��ٚz�s�N�-���$2����p;��ٞ���u��fF��/�t/��,u��� ��f�����3RbL�;^a�C�P�����p!�q"u����Un�fa?Y����a3 ��Mk�p�Ť
vk�k�- �C�%�kyd�j�������*+3sB4+++Qԫt�ǧ9-��J��NDUakJ�?�7�WP����Ww���322�`7"�q����;%!y[�� z�o3]i��R�iN���^2H��h��&�Ǭ}�+����	c؀��5f�Ƹ��0�PX���]峝�����3hВ߫�(m8��^[�AMָ�d���/J(;d%}���0I�s�Ja�E�Ɂ܌7(ޣMN����z�w���OI�`~���M�X�R���'~�����P�k!��5��VM ��}V��?=hcY]��� ێ!��%"V[5�g�;�(����:k��ı��n{Ԟ�E���!�&`�����ߝ�~1���5�0���r���P��t"�}�K�	�|L�v���0(ˍ�o�S�)3��A���tZ\�B�Y���:4�s�+sy��+PV�샩���,�:�H��8�S�붃�A|���e��K���{�i_�	&=����7:��2�(8�~{�9 �}P*������|�ֿ:����*4>�j�{�]8Y�x���{�P������+"4�nMۭܱ1�����acX��rJ�{՗�!�|��1W��OK#GeG�ǽ��,��2#ٸ��=�*�K�\�]�P]I?������@A�2di����-��o�P�*�� ��;��/O�2����=����D͉H�lbz�ϧ��c'�	�YS^�⇹e�O�z�����r��_�,YO�}5���ݔ�rk�J��jy���U����u�Z%������=�b�!�M�ص�o������h���{��q��%m{�YuLIO��A�e��i��;��Y���ח������%��'IUX��Ai��k尬�t'
������$L��{bRb��i
���e�߰�?|�6�QN0t	�s�1�ȰS7�U�s_�ԫ�lR��A����挌�y�cqhmR�+�1@F]��o��=&7�_�Ht=����cum�E5�&����4W1и��צM��"z�?FG�O�x/3�m|#�#�ӒM7)�k��=�����&���>j����0�@z,ի`ws���X��5x+���G�:r��$9�]�畢:����=�$S�P�� A�sHWMy#R���::�
&������>Y��/V�X�Ji��54�,� +��N^�z���we�\d%�������6����Cxv6�r�a`�j���~��|U`�W�C�����Cu�9QX=���O��՛t�����R�j؎1�ݐ��ɱ���ͷ]���[Ӧ��VhŨ�w��;��bzQEb!q5+���߷���1���C�����>c=��+��OA\XȽ� ���,�<y��p�PX!�t�~��pύ�b����n.����;����ȪR�
�-���XP�ݩ���-�f|C�E�H\�N��1	 ╾ً�Q9`&��Z��;(�}��-j:�N3f��͆]h�F�>�|�N��	�P�T�Zב��7�dY��i�W�oY����{��}����X�Rb�ؿ�IF���;>6>^�M�I�ƫ���k�4��m�+���Y�
�|6q  č|7���gj��,��vP��!�`�?���T��	���[���S34L���v�4��'o���aT��o�z���_����s���92�·xI ���9���i9qLB�FSJ�i����ϰqp�(Xׄ)viR|Y�q�&tg�5���^%	������ӥC|����ʺ��~"F�=|���.���;$N�U�d������'�3���a�Vu�:&%U���AFK��=����>�P
��&]�����nu�b�İ�b���R��y���G^Ó���&X�N"�}���-��DK+�%�SJUt�5;�ߔ��&+��c�"��MƊ
�p�mw�/!�}���gDM�ￕ4�4��2tȵv������Q�I�����"W� �^<��t����( ��p��@���2�a���r��Bl>^�����˯��F|8 D7�Oep�/R��t�z5����8�C����y`�DX����'>0{���1�@C�<����`��`���U����:�9���d{�,r��Ț�x@�e�N�P��o����xU/�u�	�ȶ+����z����N�4�rV�����f�?Zh�JL̗���P6m|9^bF ���ӕ�bGm�i�Fs����s����40	n�b{V���U��s���8=I󩜶��	��-�<Q�1U��7����AEӳ�@X+'�id?Qk����BX/
����xm���$�՜�^N5��|�L"ӈ,���ť�E'���|���g�Fz�鈉���j�uD�1�}�������e0��9�)�C\�>�:_�v����&'��;���ƮN5��d�c�5�6�(�ss�7�����ܟ)o{��A-��Y�?p��@D��|�q���_p�u�%#v�;=Y����M8J�m��6`�-�]���r���ʪ l���\0Xe7 ݇��_j��ɭ�
��)��Ґcu��D�ZZ���N���@��L��>(4n��N�#g/���_	�����k��[yČrVߣ��
ge �!_��zm-��Z<��a
0i����P���XstcDDl�
���i*����G�<�?Lm<//���*�2���.C��t�<���dm��p��2۽{x���b�+}Ll,�ߡ�r���~9��3A	z��t����h��YߓHd��0�����K|nKO�l5Ҷ�i��:�.�����yXӪ��iT��D��O�j{:Vf��sZVV�A}�h���� 3��b32�sתr�,4���i���j�����khkg'{+@9���rn�8W��6(EH�`jW��XM��#���P|	s;	أ���ьlll��D��q y��ya@��.��_�����)�lwz��T�Q���߅���;����� ��Z�X?� �ˎ�lL���\vӞ����=���/����{Y���M#�n�Ȩ5�>��`��+q�;��C����������1���
��1��N��*��	腺�yVWWm�&������1��4 �������\,�i���^�)Ϲ�/I{�x�B,
�O-ѿ�q�);� �eA�j:.U-��*F6q��K2R��<���.�wT���փ�3�XÒ����gʄq��7�!�{�VXӱ~Cn���~�u�~�[^�JJ>d�rR3FβB�
p���!�G��P�Y���+;	�`P�ͷ����n�S�+a�V$W1�c �MN�m�j�)��BԖ�JP��7�	���):�]�^F���%��3���A�����0����+t��)�0d��q^<��>->���S�O�y@4O:�^�=��~��X�Lh0vCǆ��uo�M:��޲��5�m�P�E��Pqvv]c=888.b�p����vG3��]���N!&�v��T<R�,�C�y�J{#.s�@�B�X�ć�.����c�5��b��՞�e̯P����$�'���N�N�t��R:@Z !��˲��t��kn�0�,��k;@�[�Ko�jii�Ø�e�&^���ݦ 'ςP��5~�z˵3(��T�
���Q�4�� ܮ��*a�>����������ʤ�0�ձJÐ]G�չ��A�_n��Ozw	����bZ��&�Q����r�����Qj� r��D ��P�B�e0W�4 w��$p�h
}8��N (��lrg�2{��0�L_CE�,;WGkj�����c����U;Ϲ;�Do���ȼF��gdHM�n�C�{s��fe�P[>���� ���9f �B!t��_����=Z�KT��%��+���	���Z�J�vg$c�0Ebnc��M��[��5���Z�--M��Ct�℄���s}=��&>&�9�~1%�mO"���#T2���R����3���R�tN�{�e�[�P��|}��@̻�3�N�o����D��w���q���B�Z�;i��Γ9�+b, D����IɆt�&��U��ra���@��a�o7�yge���vG��}��d���8�,����	H(���߿_ ���Iv	�]dT�o;\����%���y!��(��`uﱳ#O*��_^����)����b����"4W�ݳN�
�o��_]�Иn�C�p��4f���[v,w�n��%��A���J�߅��#�fl�&�Ձ6��V�_���)X���D}l<�p8����TPFf�y�(-��_�ڣG/�f�~��{\\�C	�?be��}�6��B�+��d�Y��W#B�ܗ.Ô����p�����DA!ڔ*,44�u6j`9n�AP*S^yy��*3���7o.�DJ�Q��s�VS�]����F�{�Y�N�Q��j���jC��߿ﱰt��I���e��9I6��?���ω���5����eH]�����p�П}I8�N@hd�Z1ݲ�m�F��@e����Sq��d���.��;j½7�ӣ�m�J =�[���P�#�r�g9���P)d`���q���ϸ��m6W?���KL�.�7��n�5E%}8�	�<��,��D��mc����'�����b+�+TV�j��˘|B����'�}܋���c����l%�tn��ۓ�_׊ ׃�i�"(����U	#��r5��:����[�6��@���Mlel��\K����5�h�Q��d-`8�Ǐ��hA��s��B8@�o�0�n��� �T(� ���>wIp�GI���x;Wa�+*��Ho7GG���%,+_�jF�T(��>>�d[���}Ď��+��l�nH5O^����=D#`�� ��Ӊ�.<!��@C*ٵW,���M�Iԫx�6tDa��hj!�Eoj!0sC>'=���h�Ѩ��	e�ݬ<�&W���*a7Lq˱�py@Jm�RLu�3q�.-�����e�f�����݉I��UR���s����?�����n )���Y���sq���ӧ�c��*��L�70#ۀ��x�|,9qn��XِBB*�Cu�lu\����X�kP�ZЍ#M8�ƞ�_��O�x� Q���ҌVS�^�CN'���#�EL�-��p�,!�	U;���V�������ׯ��d�3��Y�vuVN�-�%��	4�XYyyvFFiׅ�uk�����_ġ�on��{O��P;t}�<��@�!�j���>k�|���{O�w���bgc��{�W�غ&|��'�>6��+���/O�g��� �6~W%�j慤՗Q;﵆=�[O`hM�xL��G27c�n��m=��FQ!��Y��� ��[�&�=y�hG�A֤"�%44�?ɱ1ϵwǮq�^ �*�߮j|�	��%jQ�/��˙%f��4�G�V�g�vVr��Be�;?qsKF�軹գ�!Հ���.J[�{"�d;~A��5>)����\d�Y���ƥ(<�]��]������&=��74;�����0�JMͿ��`�9�ۓ"�s��͊1������GU�@8����tL
�����?2a�OY/��Hb��i�͟����M'������7��:x�����TV��;�:L^���"�͎��D,N��{z��¹ý�bN��{""㽡�}.�����
��n��7'�}P���J��
�dᕂ2jl��ڙ�k�V��[U��PZ`�T"K��S<R���-�4�JtΨt�.�B�qm�8��c����C��^ѭ�(Q��
K}�ƀW���v�^"�E��6aD&A�Cb��1Η�����3����
����.����z��ȓ�n6�m�`�� |��tV :��4m���@�3*����N/�[���-n:���,�R�m/T�,##&�r�=���U�Q�����pg��V'�w�_w�VI#&����Z�7&�r��|��,���Rd���n�������:����I�.����5!�{,�.8��s�R���M��-9�����qU �}�=��n���c���51���׃輗���@8�nv��L��֠ڑYJ��UG�]n������878����Q��Hcg`��:����(om:��ӌ�"�}Pr���|<�*��<&��^�:c��uyQ�f���ƶ����aO
JVA�g)%x�hkkڗ���U\�I�d`�z�����澯�?�Az�x���A�Ie@F���1��6+@�[Xd�����3��cL�*�n��@j�c�)��ʨhiW�h$]���*��lUz�ii�)�(�َG���;�w�~���{u�8�L��u
�v��K(H�3>��k�Tf�z���;��d]U�HQ�����î^�J-& dEf#�G}[���RGK��+���2AU~Om��֪E|���6烱
,��x:幡�|��FgQC��6���s�p�Nm,_���*����(s�����������m�B�)���27 ��u�Y~�_z��b:FW�6=� ך��[��n�;�3�J�^xx\myr�K	��ܰD'G_:�(���I�د �~F�aPY�Q����l�����2
(Qj���0��}8�󽧑��|81v�x���v�ǉq����Utv>IIDNw���2�y���3�o���!�z[گ��H:��$�ݭ\Zun�ϝυ?Qa򟲈�c��kS�_<'��W1l��k������\<�����k�Zx�a���Ӱ¸Q���	�3O5���P���3�a��hj�������Ю���!��m���\}~��46{*x�뒮�`�!D�E�>{���O2 �lE�rs� /$M�%������M�D0��s��}�jN�Zш�0$@��Am7���ש5�@��߻�"t;��՜�¨�ߑ����d;6a+�*Y5�������}�ϜK�0�mgվ��Rԫ�����C-�^�Sx�>�2��J���Z ;;��҇��:&~�g�\�~i����P[[_���j�M��U���qǦ��]�w^�D=��?_u.0�(�x��ӓ#���� &
�fSp�n@w��������LvLIP^|�P}(��D�f1;�	$��ٸ��+~�c�Up�K�ս
��ll�И��v��H�т�YJ���w��)�8��76�U�� ��#+ۃ_V\���8�C�=�"O�j������1q��K�O�c�����ۏ�K�}.qp";����z���N��O��������^�����>\΁�������@�����)�^Ze�I�J*~��ү�w�He��0�&���©�a������\�h�5:�P\���[h"�i�v�aT�[�mUTQ�n�Ǻ�,�3i��ۏ��X����ɒQ��S�L��yTB�����ߏS����������M$ʹ�8����
���Oz��A\tt��|W5� ��6�~�<x�\Ļ^��ȷ�Ѓ��M[��h�A䝕��* 0���w�BY��λ,��Bח�`��:^��栢�Єu������W|k�v��#�.m�W�
N�P�X.y���q\�� �u��yx��j�&R��q���Y�J!��5�^E�<���yV��t4�EMO�Ӹ�`6N��*�b��+���צ�6�r��'$�Υ0�4�4��#!"�Ƒ���`-�4l����|��(��i�d!W��7��k��MSK+��V��ˡJ �xc�����űj��\b���^�bh	a��h��?��E�(>es�N��k=鋳�ǿ��1K�������KA1���h���,�2�ta�1�(	�sq�8 �0�L@�_
��Z}M;=��K��uz�=��g��"9<H��sy�f�]e$�_ �P�zuu)"2��5/�}o��Br�]X*�ˡW*D�X�mJ�o�t�E�V � �һ������ b�T�Zo%�ʐ��'�e���ra�/IN�\��J3I�N���B������ȣ��b����Z�:��������%G��=/ǭ���K1��?��iCvJ��Qf���`�#%t]"����٧/^�Ϻ��ۺJ8�#��;���3#L=�4�7td�
�_v܅	Mw�i4�i�C�S-�O�&�����i ;>��"�ӂ�|��}��S��\;+3s��F`�)qT����W������ ��T<F�kLD����R�MON�>��?=�kj���S�u��8u�ڶ����6v`��E��{� ���8��S\�(鴯����>��]s�Iή��b��8O)�b�W��wi�؀�D��(�z����
C
I���|$݅խ���:��`݋�a�v��ǜ�/ eIÚ�@�5�M�dj��I
Lh�ot��P�^o���������O<f�A02T��k][>[��%Vځ�g�	�_�i�kh���T�_����
���'Ó��v�����<Qt�fK�hA�^f�C���S#^k��5��o�d�))��]P#���yoߚ/n��E顶����� C����֔h�4F�袷�ϑ$�������[�d��������C X~nn������;��(�	C
����eeQ�I����ʔ�&"e���I̗���#���w�v;v
�t
���8^1xG����Q�+k����G?���ī���V�����S��ӌ$����� p����V0��7BZ�32�@I"�ra�y��,S�x+�w�tX�%��}�B��
�̫	�s���1C���W����&.|%HJ?�����	
`ì�6�g�G�k��W�a��-�Ta�%����~��R?���0�Q�'�m�S�PP'R�L�୐EKp< �ݾ�����$�� ����Z&��@��zu��^���W�LP6�)D9�Hc��<R��v��U64�Ӛ0Q�v���H�������@�x�����mZ^�kwHRAE����J�F.��6��ֱ�����$��j吔1�I�E|ʧ�R9�
u�/^���M�0�Mp38�A:X����GQ�����,����HydR���l��ٔ�8��_.5�����6��x��r�8{�X�S=�%R�*x�!=��DG�"�5:�?��!z+�N�Y�5�f�}tQ�F����� !}����v�u�۷xYp�=NN�lk��"�Z`$�2*"
��]==�[4=z	Q���h3����[�v���)�?������y���ܚ���rV�ŹE�]���ʦF�z(tŔ��L�J���ظ��3�.����.*���׼�:ѩ�q��5�-0`Xl`d�y���C�}'DluO�[&�';��@�8�{y�̔	�"&[��ծ]L���nK��)Ϲ�a��ys:g�ГE�����#�'ge���F�.����T���H$o���e����<��hH��Ma����#d�h��������ގ�����w	i�}��U3�q�ajj������I����c_h�SHH��X���C��l���'��v�����.H�?��-����U��pQ"���w��[t�7^X��R�/Yn��{�
���<�B�/�O��E�{�ncKI	��
U�e�K����]����**)��.��/��V�._�s���$XoӺ�_P�cn�t6��x��xg�_xo�ug���\c=J��̽���������uu}�C�O����226����~>�RPVQ����w*4n+=q[�|�
��D}�Gq��6����N3?c��#��QKf�b*j�e�MG��D���b���1����^?�,/�B�P�Ha�6t���UH<�à:7;{��m�r'K����I�'��3�,J��ZlKn5ͱ,�7�\$����_�ۣ
�F#Lu�$b�O4JRS�"�|�L{��H�ӫ .�8((����pp�I�{�z>8T7����䐆�v�L(&�+4ŗ�!���(���&��q��a4��P8��P��ku����M܆ˎ���.5�T��t-�6��Y7���ӗG���B�I��T��΋�L�&�(F~̡���s����?���"��$V���� q�j�EYA =����J�� a��^���ɑ�QCj��Ű�b����07�&*���t��IX�-C��o1٪����$�ۅ�UJ '��ٖ2��W1#��UpV�ǑJ�^&������O�������9ԯ�=��0��U^v��uھ����1����qn�}2��Y*�0�.,gF�7��yr�1�
�ֻEe������)i�%pnadRaJ]8���N5M��D��������!���j���2�2���[�)2�W�����S�R�ڼ?�O��716ͽx��0�ͯ^��Ŗ�Ӭ����������z{��T�bʘ�o(��9�<���klԣ���}n5�'�u���9��������D��n�qk�b'K���Ҹ���zR���$��ť��m��6|����'�o�ii��L��(ڎY�ײ��W+=�PhA�B�������Nퟟ���>�(����"���6<���}bA�/�)���B���EÊ[y9�@	u4Z*Lx�G�U���F��h�")�2�uK�;��_^����O{����l��=ז�..Ǵ+y�~�<a�bQ�=��GF�=�;�훊zex'�Mo��vH��?Z�c	;�����(�@K5�8Z̈�"�O:I�7_޺z�F|��v�J�g��FP�<�;�K�r(�"|&Yx����r��La�:E[��~�N>AK6�$�޶�f�l�}ǀ��q��A/;|E\M���o)���]{T�㔚�?b�,D�P�s�meEh2��6�{f�#���I��G��W� �/��p�i�;���T<�;��6���_�#�N=��/&{�������N�D�Y��������@:�sF1r3ٮc��XM�2e���3Apa�}�l[� o�%Ỏ��#iܽ+m���h#�`���:��k�%I�F��F���z�Yt���L���t�j�e�����|D�ej^y9�P���h��;J�!��Y8��wr�E�H�b���u�/��i���N&!G7�)�Hs��P��ѝ�YL��V�gҥ����!����]V�/�mYy��p�K�k4.1co�$�רy<| *�:��J��/�~;dO��]��Mڒ�T�wq���E�n�o����|�k��SΆ�$b]�aD�w�4��
�����=���E~�ۗ&.ܼo�ZI��d��dZ�+��~�8�^�_O*��9|��0�5�2�w2H���^��,���;9Ơ�10���Ϣ�*�ōxݭ^up������3Y)�h����u�T;|����o�h���D�R,c=����w�S��?~�������C22е���?���.^n�8k��\���b��Z��Y�qk:�d	J����JEOb1Z�(Ɔ�WT3��$$L���.,ws031�%r{����#V4�dR��[-���ͺ���0��?_����ap ��%$X���X�c�����x� �22�(bTkj��6�	��ocX�)�v����T��������㇈u����u�$ڂn3p���S����rf�4��W�|���./ݔ� ���yn,f^dw��Kr�����b�W⻆�W����t��`��_���͒��/�`nĻ��b�T����K͋*��cv�'%�R�����X(F���P����W� B���{œtPω���cݷE^	���w��nٌ�eҙ){]�/	؛���n��v0T���d]'X�!ѷv�z�K��F�� ��,}ZƸ�Ǉ��W�c�)+^�J�AIOo�w��̀I'�����������IO��-+#��=
R%##�:�x�W�j�U�K͉ ���T\ܟ���g/��2j��#����ri�K��|�C:6��"|�7�D�����ZZO'�.Ra�	�l֤ml���)���cz=YŲ���͛zs=y�@�����j���9~2P�ʶN|@�ٿs�ɀ���kh������}�v���111���ŉ��U���|�9��â�{��B�1��̴��X��̵��hi)�xrH&t3�M���%���"�ߙ��ܔ��w/)).���\Yi�#�ļ�VH�oNp.O|5����Ȱ�=H��4ei?)�����e���Z6}�ٻ�µ��b7��M	��QH�|��`�����W	ľ_p]�e��]sm-��f-M��	�=���:ʹtV�w��x=�@�����xfpN�*��Ő�I��]���p俰9p3}R�'��G[����`U̹�s�ǎ���/QS���]|#p�<��/���"Wm`�X9�-��{*��ڙ����M�×Q;��籍zz��$�G37����#jM��Cu��1���#�� �t�=��4@���ZZ��� �Op���We2�.�Ԕ/�ц�?x�29�}u::��Օ/����2��5��E*������|U��Y���8R�mo�A����a�;'��>˅U�o��
ħ֗�G��_�8����A�
�2��,���Mu [YCM-�m��W�S������[�8ַ�w��e���s����&��i����i/r߳a�׻��1[DS��[}��Щ,Ř)/y���y�D챗�2c�sm�!�2��4� ���OYo\T�ӆn�TQ=��>\J�g���;y�Mb�&����y����v�7d�Ug�W�
/eF�#�,S��l��/�Y��{�eD5��>u0A׊n���OzH�N�C$�U�Y�)���$��.��,�n����uL����i��^������~��f����qN���g���1����~{f�si�g�G����Xz:�-��.����l+�D�s���8�Y����?�	P"	��2��Oˁ���``xI��/��o�6g�;\�[���:�@�<T��?ƽ� }eP�i�źhm�n�������[���+��#������ڼ�W����Tc��p���9�bV4~zdS��S}6�Ow�R��d�i�}�E�K_�0sD�v���8���>�ЇGZƪ��SP�Ҋ�l�V/�>9\���|A�l3�Fi�u����6l���~4� Up�,g%����i�)�϶�.��.;�
�٬��rUS�ɡ"��	����	�/�AuLb���+��_����
W��Df)Q"�ǰ��7�]VR���dZd�)	��Ī��.�gg�G[[w���3�Lo~�3�|�=r m�`�M���2ƴ�U��/GP8�|���D̸&�'���h�o�}��1��f±����q���W��6�g�p&��V )MtS��+P[R	�;0dJL��f���>�^G�]Ċ�cDϣkC�W�)�U��x�k|S�_8����0��ŵo��;�����Ҿ�y��|<���Q�8�乏������#�B;E�@.'���S�-�=�ä��=����ߞ�{ʺ��b"ǲz�S=����_9�B�n�\��i�\Zc9�� �T����7o"SŴY�c��܂�\��(9�Ŵ+�mgk�����L�,��*I{߅��l��COO�P
���G���V�{�vqny�&��J~��A�UخL���rT��}f�^G��m������C�����!��E����R�a��F=*A�P�VI������WWb2���[�>ۆ�K߃�*i�ʮھQɁJLW�-�!%t�CKK5�qt;Z���U������(�E�T���L��FWg���u�Ԙ�n����s�T�
~}y���	Z󥍆���e^1�ow:���EF�k�Ւ�Vj���``O�]#>p�c?٢�^(���`����/�Q~O��R�޽����,���<��p���C0�0XA��{;�4w�>E���D_�R�PS�cmϲy]�8��QKv~~m�$essec7j�}��xvtA�OuC�d�����_2xW���z��g�GO�jPK�.P[O�
��չ�U~P����D�6pT+!�rC��VD�� �u45�EG(+`��ߘDO�9���G�E��n8����͟���k��/�-�MK��'����Z�w;9(��J�GӸc�	^�V�qX~����cy�阝ɏ������f�Sm��1���V�c��TS����O]���I���[�5c�Q��3�o FtOM.K�g1g��s�׷)e�R���Ob��P��[G�S���L�[W!_]�0-��-�;U(�!PF�O��$��ЩR�t���F%�/��|���e�]g���~�u�Z�*1C{f[w�:���r͵=��+?�?�����!!�c����D����0$[IXC�Q���͔��W�+7A*���3Z��гIli5	������	N�d4�Zy��\��a��Ixͩ��0��l�+��~�+E�Jm����fiL�6,~7�R	s�aB!�{�f�����f�3"x�-�g<,��e����Ih3�Y��ʤ��Vn~~��o[��E�*u�À~�l�?�dca�������>�>r���n/R�Bv,{3s�F��(�z� ��`����Σ'�1$��
�h�5�S	S��a6̛��O(�#o�r���҉x��6 �gW�["L5*�f�C����:��N(��J����������%T��|��c�Gy�cG�&=>���X��sn�7���*�-�-��&�2>.^]�]/R���_^���7�k��G"u��:�����g6��ϸ'��4&�,E��['�#s������V�o�l���:�-�_��I�Hk:Ū�&�K��WZ�_[��*n���ܛ��ZJ��w��$qou��񧁌��Q�"��˾1�M���/��y�?��*ʠ�XJ@@��n�K�DDX@����\�N%u)钖�D���Z�����}��w��9�y�Ν������33f�z�[���o6'�6�h`���J�{t>��l�y˱'���v�>YY�P�f�p6���F"����{Q��e?2���;��z�E=h�^Y�1c�'�j*�o��.(�����N�+�PО����\ jgh8��f�s!�^���E��[r��v�� ���A�%�u+�.��SW�גx�[�4��ݿ#�����Km�Q��6������u3��?�2�V����<OX����^��Gc�-�P͉o`��T�@�6������@����G3o~v[W�: KA쬦��^h��.��Ͷ��T�G�R���m!�	6����|�޷��>��|ڵ�ax~JD���-����K%�è#m@;�[�9��!ӗ�jȶ^]��1�}�q%�uR>�	cڼA|�����{�U��Bj����ğ�{��KO==���lN��:r�4�CI��`�S�=m\�g��/ybq`愔���J��>��btV��Y����A�@�u�;��O�H|��ŗ|EW���^���Mo?�a ���p7�k���Ȼ�7X_?�٠���c��_lg��g�n
�fK�)H�]��:4�2H|�Ń��1�9�j?ШH�:�F��R�C�!��<r��z�f}n�9��4�!3v��Oe�H��:�<�{����%��С�&y��~��S����fp-���V']NGA�rHd���-�\/�M�j^vܫJ����I�2���l�p �� ]:��,���Q��� �=Eo�,���8�s��ܪw�~�÷	������Y��?������W�+[�������?��7C�CO-�nK��8���3&�{R��{��6Ŷ?K`y�vl���$�u
��o��!��8y궔sy�1�7�2�t���1wۖ����}�#C��Z��,��T��Ϊ��̈́�Ә���!�B�����9�{��]�!AX�q����5������(4Ί��m��zP�<.�=���Y�2���qm�)^,j4Ҙsm���C�l��$�l�%ׯW[}�������ǀ
�s�k�[�e��Z��[���ޣK�,x�$��y������'$L�;�����8��A��EL��S�J@0��J�X ��4�>�����*�""f�%�.��V������GpXH��]I7�}��	&����A4�&�UЃ~�g# ,��-<A�me@Xi�1ss�'U#(	3e����T[��N�c	rKE3�q�l߆e��93C]fޡ�Xc��E��tL!jՏ��Cn|PMJ�$��?�&0.�0�~�=9$�e��D��KO?�ݐD�� ��Y�rא4v�A��{'�J�ND�U�)��g��>����k� ��uO���"���8������#ȝ(��_z�$	C���Lz|�\����g�����j�3��m�z�/4b^j�
HC�0Y�z<�9�kF!y¨Α �!n�����P[\n�8t�dG��h���ss�;�<�I���g�Cƶ�z��º��p�o����O�Ž��O+u�����Z�H�� !���ή�%��2��If�v���gZ��O0�Y�+
�q���PAO�~���69<�~�9�&7�:Xyc��׳�-���¬���N�V���=�8���@P�#������p�������I5g©�"{I���8�>
?���|7�H噙��8&.�Y̠l��^��r�9�drB���ͤMF��i����k�w� ��28���̦E�iu9U�<��~ǏұK(�%�>�`k��ηJx\�H�S��b#ix-L���䇺�1g�����&\� �y�(���_���}�ݦ� ���*��>H�NH����c|�ݝ�ͩ;�+x����E��.���C��w}����F]Ț�H��Y��(CeΪI)�6Nd��"�����KmC��T���t�T弛(�,A$��Hľ�.-�z�_K����Ѕ �7>��{(�T�_���;\�s�B��	�����83[�>���y�����j�;�`Z����E=,��ϰV
�����~x*������0��D�?&�\��f����u�7��B�KLs�����4�]�F� �
�w������`/����+E�u�>^�>'��|���=�����w�=W=��(��{�wK�7�o�?��{���f|jl�FU��\R����~R��k�����D�wJq�8���/��]��mt ���3�jM����U}�Zʟ�J:Cs��>��aLz��� ��hܝ0���E��ga:zT/���I,�/�)���8��t�ꉩI�3�H"�����H�ҭ���nռJy�nV����1aHz4CA�6n��][ *��lr]�%��\�pKF���l�3=��b}qFrX3K/Ģ*eA�	��C��!N�<�o~�k�s_����*���qTe�s�6#�����c3p���Ƿ�̣�^��x�w�]?���M��L��Œ� �=:�e;��G=���|�M=t5����7ǜI|�I'�~{-�n�I�Z��3�n3�䖻v'JfX��Dm�3�1 ģB��p��w���G���Ee�o�mh�捨�̓���^�|X���6���2�['���f�#��d��o���H�+�W6����d-i�6���|���l�����Ƨ���9Y�-�$��~c\œ���]�|݉�f=�M�U+���&'�W�����"�!6~�>+��}F�%y�WQ<���:�إ%�mHV�@w�7�g.����~e{�����1�\h$Z~T����ӓ�wҘG�<VB<~�����_�ٖ��Z��{ZOW٠��IJJ*��.�S�Y Ǌ��j�/���гL�|Q�HO��*)b���dE$x�$\��=�r>���?/TT�q��|F�d�^�O[��R~��U��WT�q=�/Ρ�!bs�@� �a�D>���''�E���h]$���Z�:#�RJ*[C�#���Y=�)Ұ{N��3\;�,�>W�Xf^�s�#6����H.��s�������q�¢��c��G~��Z^&=��Hՠ��Ŷ6-�V��e%��|4X�W�E��Ie��`�jM�� VJ�ek�J�pB)jxk<��T,�ߎmp�S��ئ:�G1��G�<y��F/�\�*�g�~=H����.���(�\�t��i)?����6e�D�x�>���don.m ƞS�� {��A�s*�k�y�I���B�S�DΡ�A�Y�v�J�F�߽5�h<��ly������]?����}bz������۫�wkH�$����!�c���4�@5?����p%�]�r��w�KLbi�P[f�U�X��5�M�R�yD����o9���-�߶P��n}��CS��叜�"t�"��A�J��2��Hl��=� �D`�4�A3�FS��M�*�Ɔ��-�_�1��ݵT��P��;��B����#�Xo޷�������
a+��a� <���4}�d�EAm���G���Y��W��R�L�;�����E��4�����np��o��>���*�,ǜ�ĉ�Z`��8��:|_�f�"t�Ͽ���J['���� ��Q��m�m��f�zY� ��٥uzk�Q��5�j�_E�UN��{����72u���sP���P�nZ��)ˇ�W5���@�V���^̵�sa��xT2���ڭu��k�\LQ�����B+J��g���v���R���RnҼ
Tal6"�8gr���wg_��6�[�a�!��;���z� ����Y����x����g5Q���S�TZ�E���]�9���<%t� LW)���f�vr�6�0��:�p�H���q�܁0�^��$�Z�e����x&���LP
%1�/�$�����7g��R�u��&tq�S���U����r�ݠ+��)��K��Ž�9�ׅ��RsO�*����GJ���x��e�~��*SG��W��陛���! ����B��M(��W�}C�����Ǳ�9�P�`���奦�0�~����̌�R��j��b]"�C�pSi�d��Wzy�_6����נ"�+��m�&YȻB�J'�t�M��j]~tl�`�j�)����QT�qw���;+�Q���O�s�D+�kN���T�5����������b����&��J2'cک&Ÿ�c�7����v�j�^U;M{�s�}|�ki� �~� ~炵8Ueˠ�xSP��O�<OcAon�L���-��8�/Es��;���}|u��������Wylԁ�S�+��m��mDS�]YZ��a@,}��j���ߌ���km�`B!���e4X>3QFVa+,/���'Cҽ�������/r�׋#�e�O'�B�^�|��,+#���Y���x9�-q��Y�q�2�p6�,���\,��DKvW�W��<�'�m����0S��>[|��}Z���	���*������o-_��y�:9֌�Qj1��"�F=��4r���
-+����;\+�>��K8jPf���n�VΩ��ܴ�{��M-������Z�}��Π�#���s*jme�W9�o�_���HÉ�>Y �(��\ p�m^d�'������n�m�FW%�t�NO��`��I:y�\���	�6���7�NQ���q � ��#&J{�e0�A���K�<�F����_L��\��ag�k���p�'��>���*���TY���t���:��pz�̼��$`���5��&�����'��Cg�3�Mlਙ;�V�`mt�%'�A�P�,�ڃp�A,��s2ifM�ۼ�M�,��}��Շ<�92vk����3ǄO-���̍�|��01u����JCW���ru���Y��cH�����~�ټu�l���K}K �J��w)���y�̻nv��yJ�Qp��(�����W���eSFْ�����V0��V�m������&{޸��>�7QG��:�"d�b�Btty��x�d�g��Y~�D�Ц1}q���8(!��?�ī����oW�|k17�H��^��䇏��HK��1fnC���y��i���UU���Y��k������H��sy��X��TO��<n-4�%ⓘ�_��?�,,�n�]YB�;�P���Wo�����óu�=����7#�E�N��<����!x��]N��!�
L�LH�s�l2S������QG���o�t��v/�)#����t�&�
?�
�������F���"�(�e%����L����1Q:5n�nB�E�Qp���q���Ñ�聹2c�	ӫ�F�b�g���T�X
�Tt� �;�cw���L�b�gi��J��W	sO:�nM'j�A�\�4�bQ.n��������;�-��3ꈺ���+���������� �� I���2y�|�����ʋ���j%P��K.����ԵX�?0*�?-�4�N�U8���>�y��慝�&Y���U�ڎ�B�"����XϾM��x6�����7�ŋ:���ղ�b�?F�^(��j�Χm�n��I�������ad�5oɉ�)�W�h�ss��.����W���}�d��*��s�^�7B#��Jlv��vf���P�����b�2�Ph��zg��%�W�1ʔ��֯�\n3iv���^��diA������q����qn����O�52涀	I�>�n/��&f֕$ܕuoB�Y.�����>�J	�!�V�����^�71{7�;�����y��@�R ����{q�ݶ-ʗh�%]�@H���	w1`�8�#��@�B��9�?a:�4!�  ��}h�f��_�����B)�+c�z�A�c̹4� �:��oŁ�pJ��Qcc���@����/h���£!p�-!ݰ[539`A�*A01@����"q�(�����[��*u�d��U�)6s��2PBѧ�	1))����便�:�J�����F�ƛ�W_�u�t��1�$�������i�������2#,|��$B/}����ƒ?�����"?��ɉ�3:��O�]�Hk|�sǚ ?L~����-mm��))�]~�p><�g��\��\Ĵ�{Y�S}/�[n�@����6��L~���^��+�W��j<�?9�0@X�>##�	����>0�"��|V3�'h��~׳��O���L*(9�7<�G��Б������/�~!ׅU���Xx
��VDI��σ���g�9�CFC8s�Y�4�m'�%wac�B:U��i�%��`�bn���������/��a��@I
�G�g7���n��7w��h�T��`i���%5�RP���F������E�i4�{�:G�I�bߒ�`z� �9��W��SYf�06��8��&1"�4��e9��;%k��G���p��o�T����J(�(CXvT�?3nC��}!j���L;�$�C�`y̠Ǻ��q(�0��9���n�,}��ۃ'+�s^���φ>H�P2�)�u~��z�T'�G/X	��Q�.u,+��L�����G���T�x����3;�#M^�K���\�-���P���S�m}�C(d��|"Z�[:�Rذ�[9̍@�ă�T���~���ǆ���7u��Ъ2�[Ĥ�P�8�Vu�R�^.�k�KS��G-c�y� ��.[ш�������~e5����f���?�U����g�O}=���5@�QAG���{�U���րm��-u�Yo��r�.^*4�O?n`�M�IB��b$5?)OSE4r���/ť	�!�����]O�����턝y�
&�@���:�s�9�����.jD���x��kK�)�)�)�g�Y^��x?�Ϟ�P�"Z0�"���N#�>�ܧt����n�1\�ШPP�����x��c��h�}�i�%�r�3��L8?ni��;��ޒw0���@��Q��*��75�/{�@Z��:&4��9�a��#7�A�v��Z ��,����U���fb��4fj�����v[5��Oz��b�b^QU��k!�,<�֌����YpgxP��6�a)����΁�� O������y!qLcq�iy5��d8�i�����_����L�[ԃ��9!`�.�����]����fr+8nbቡ6I⇷�tx��_����?	I�e(�=��?�!I��3�?�R���{�s����f��[������_/fAa��fAF��}3���t#~��F�Xm��OX�YLe,Ύ݂��&
a3|�`�Iy�{������S/M��9n��u����F���|�ڐT��Y����X�wܵxK.�5��<���4���c�EB���}��O|��|ſ"�&GQ
>�F
�����%ٳ���d�`�`5]�^Q�|%��߃ǐ�PwZi�
���q_�h�]<���A}�|��3:؋I%Q>��srbɳοjy��{�$�~�F������]K�)	,��4�'k�/y��A�5��ҥL�Qh�aY~�-;ʋ�֮�b[����BK�&��S����py'5�����H���w��g|�����
�t*��7�`��ȓ��r�O��mTPau�(���	'p��{ҏ��~w:���Ǆ�TP�dŶTC�Ӎy�E�)��%�o��+;��A�A��z���x�O�yq�1��,�N�j�F;��
.D7����M+iJ�b�ZA����&�%�V<��c7�:��ؓ��`F�d���*��`Mz㪁�����oZݟƆ��[#�d�Mz֧
t�����t[�-2���O�[�I�>�V �xQ3}j����lr�Tl_�5n"��0��7��뙔"�`M���Krt�Mz���L�����u@1')FBOO��M4�֥��t��2�2�L}Hg�.TΤ� ���.��V`%�ħ��r�o��=��i9(Hr��S�pVqSً�)��Q���L#���Pα+9oV������F=cFf��>V�s�̔���j�%�����5������OGC��+� kQ��[3����Y�������=���ex�W�8��Z�W��I�A�{�E��5��n��H|��P.!��1¿H�ŬB;���+IudbA��N_�c��]�V��2���������N��וa�2���x�< +!��R�'~��%X���}7F5���2�k��L�#��jݺx��W���hk�� L�|6&ԋ>�*���:-�x�pSLX��q�L:8�Nu,zo��늂�4M�ϒnSLD�����2���y[�D���ڒ<�Of0���Û���/�Z�"���Ő�Ch��m�b@	*�s���ƪ��(�0���)�,�7a�W��U�&��(�dK�� ���֤�^Jz��& �<��#��R/_~{��37�>T��U��R4f�eƚ�t<�O�E�
d�Ȉ#s����e�g�
�"�:�z���$4���z�s1}�)6��U62"��]X��:`���#�$>��D�nAN+�fra��[�;&(�;�\���İ���Tǈ-���q{�k����Pt����/L^����#���5&�S����ƭ���sX��}A!$��j�4�� �ùNY�ٺ�K�D[���K�v��G�߭L9���
�㌏���ڡ�Sgfz�;�Gi�=϶��^�+P�iӰE|����������򙛛ȤyP��6�{?�P���ӑ��Yp�����!݅EV���!x!� ����F<��w��`������B�B,�WI:ܝ�P�Vڎ ���-&�z�TD����4(��=�Y(��,}�ow���Glkc�/2��� �|\���t�����O�� 7{?Z�E�M�! �qB�s��l�S�����L�`7Ð�ȡxm�J$���Xy�E��nk�K_��B�>HEq'�e��P�8��0#Im��F�a>�Pщ�\Ls�5�Y���y�#t��@�2��w�Wy�}b���kH�=!�z�x�q���Ѩ�0<���	����q����0�$��X�Dy^^�j_��EQ��<ӥmb���.VF���5�3o�w�چ��׭�����S�����wJq\<�\	��Z�n�<]˘h&�x�6����N��'���߾}��R,S���mUIݗ,�|�i��i�3:��ed
��y���{B��g Iʹ����˷�q�&��5Z~�	Ę)8B�I�����
�Y������",�OLI��(��k��a�JԾ-��ƽ*g{��-TT�Pc����+(	9��i�[W�0\�/��89��H��ގ���qQ��ϕ��_`C�G��S>ǡ�{#f�;e$�(X�9
�$`(�!��yP+��BV�q` e�Z,ͩv1ﻤ�Q]����\�"L���p��ޅ�]���S+��,vm��37�{ʯ𝻚q�6�����|,o��'	�5�>�l����XY�)��{7�f$�
^y�x��%~����ؙ�vv-t}.�Nk����$���kԅ�%�J��׻��¿���~�����D��J�"1Ɨ���\�8��݂��e�my,�L`���+sʿ�Q42/rP�Pq��`�O�)�e''	�{}�a�W,��/mS�)�QR�=���#^�i��!��y}r��tGx��R�����4�Eq<�U���FR�<�&:�X���o�4��P��]u1�"����q՟��4o�BD�b~�z�SL�z]�D���欐U'!G, ��`p��Y����{oގ�]eS�]�*�h��j�I�gDK)�N˽7����qM<�'B����Qp�~�˃GM�V"�W7�׳jD���rho>!_����=������oR����0���k�\9�;M��NFߩ'�s�1�D��_Vr�u�� �E��i5�D�#�
T*�f�XGo�=#S�����H�m�q������m��Xς��so,�
�ur>���UlO'�ܫ�ᶘ��K|Xz�K��~#�NR�K#�y);�.-�+������:ahG�m_�x�n�g=�񊓱9)..	[����2��E���}4����XM�`���IyP�IsYYYL7�����4R�0D+j/��:^J�W�N�i�/%m�i�jvv�F�3Qux!�:�-q;����~�p�.}��Q���|WQ3���ބ��b��'�93;΃�����j�����wa��`Ȓzdnnn�~,=}�܋����x��R�����%	y�/R�`f����#k�Ɏ>�	6�IO�E��;��4���+3&��٥g��>$�5���h]�P�qX�v����~K)"�aJ�j�����Tc#>Q,����c��r4������kS��ٹU7���$���m��eŐ�y��Y�(���=��K��y���_MUE^�b����a&����'��n�뻕�B�c�#HW���jI�Y��^@��p�z�g������� 9n;�{]/�^T8P)V��ts��f�D��y��&ϙ��f�I���=h���y$R��԰U��5��$��8�D4ص��h��*D�1�B��\�'��!�����������W���9��o&ܬ+�񀵉~�M�����g�9��涷�o��e���~$gK���y�_�?Ir\��p�1<��"s}<*I1�wx��"b�S3)콏`���F�0+f����#1�%�`�QQ���/K�CDNuv���ď����k5��'ϐ~2IQ�Y97paNH�����k���S�|.�'4 �MN����!���< �K;�q�sPz�!�+H����#��Բ��c�<�]ٚO�Ƹ��1 >j)!Oe�Ɍ���KI}o]ߒ?8okʈ�
e�z�a��Q�\�s���������z��ͦ�8�8��h<#���Ǜ���S�NB����f%�"�&�7j׽�M�"C�ӳg���F��:���&�!����#�ߡ�n�t�6�3���х �r��8�;�2�gN�9M�N�/��p��v�U���D<��yX�N�U��_�=)3�oY�w���>i3���Q�C�h�d+ss!��t���1�'��q�G�3�8�7K1�K���v�/C���������2@�H	w����7�vwžFz���H�Xu��_]�_O��R�<|�0�M��j�/������ut�ΰ#�k�g�.:���aI���2s��
c���t�M�"�엠�䠥(���}�yU�6o���t5"�a1��1�G_6����׿r��ym7���M�0�,VJAt�^����%���Ч�H����Kg�4�#��N3���͂L�	I�Qp����U���U��T�ԧ�
��j�ۍ�)Z��7�W4������+K�S]Z{~�����@xď���J³:�-�LՋ9�w�ׯ�a�Q���en`�9����	壜;v4�w�fF��'�DwUe<G� �״x�l��=8ȶ~}��+e`�^�!�*O������PZ�|�d�.ΙW��M��j��~��nݿ��U�o�2ZeS�ױ�=j=8�����r�^}�?Qf֏L$�3�r��6�
���u�K�F�Ãb���� �֛}f>��IT�����$Ŧ�Lp�z�f�2�3D���{V4�6P�U��jf.��̬t��jp$Hf�] (B��<�b`�z?�7�sME�}����X�\8�@"��W ������L`��1L��B/��C���]f��6����u~�f�r�xiWMb9�����;���;��̬�-��	��j�fʟ=�JO2�0��v�k���Y�/2羐xɓr�£{��D��	\�x;V������;�#��2�R���8^�=�>�	D�,wE?���>%�ٻ����V��<. �o�C_lISa����9���<��D�՗"��/{j�Q�[���_�o�zGs �6v�$| �Q���s�����]��B�l��h}h}@|��XKj�=���-��| �J�]��Tr}IIt��I9��f�}eO7�M�QZ��
���d,o�Qw�z� �T�u9Y�Eg�w�2c��-�� �jہ^��{e�HnZ���ͼ���d�������t`X�in�'�kk�4�w�P�}9�z�]�9�0��X-�Bbc��F��L,W��!v2�f��Oc���Z�^�f�.b����Z/�˓�>�|=[��_"|����Z�_?k�8�n�,��q��햿y7!���k�\ܶ�*@VN���Rl�-��ɳ�%�v��,�*�VZ�%���.��p���P��$�+T�Rt��zBx��b�������v{38��u��;?�gehk�&V�I/���:5�Բ2į�ߐk�|������6Bs8�M�N ��9S ��/>�i*�]�"&��I_/��l��`}��AW�p'r��%B��jȝ��O-(��_4�;#�Z%0UV\\|�}��c�*���w��]V�����O�9
~��W$Ft��o,@p.yib�f>$>�ע]֗����Tٷ��鞫�#�Z����<�#���t���fS�i�u�d>c�JS�R��z)`�kۛO5y�q)1V�h��-}�x��� s՛���y�����!^�=	 �[gg�}D�dz���]�"�w�y�?��p�B ��@"�)!$SbJ!?L��\���u�z��5�V�A���2�w��.�m�!B�g~�����sn�����m���/w�Pֿ�5@�Q��gN�
��,���|�DY��$�D�>?ʢa��ү���L���K�W&���˝��	��s�}a��y��.���U�����-Q�J�o7�Ԋ��%��# ���/�u�Ş����j�-�	9�<I0D�HޠV$�+:�I)�^����g�!<>���Q�j��"���
����Dd��JfN'{��}\�@/N
=A�_��9)��]t�Փ3 �}ᄄ4��V�Z�u��$@�xj��GN{.v<�&�ЫXo"oa$)�w��X+����&>�����m�����p�a�+ӳМ%,ȋ���b�@�_������DsV����榧j����v��Z����/�A �8��>-�i�ѝ�'\|�P ��&�%���a@�b+�?3�ҡS�n2bb���ⱉ����C�Q3I:���>��j3Nj���Ax��^����ۢ�I�y�@Qf�j�i��5K��˃��4��]�C@���J��Cz�E��8�x��-�[+�bG�M�OGѺ���C�q8�H�♿���F\����#�m��BWѱ!7��n�@�`���&�Z��3�v`Cڼ�1�����5���i �&N���M$۔��֯�-�
���E��?zɽ��7�:?���҅a��(��M~ZA}Y����p����`���9�1'#�:jU ��<�z6�LQ_p<fu61�&:$�[vQ�?A
n:�o��#D����-x���et)s����Ԥ��V�'i8;���	��\9L�5���u��}���Ka�_���G�"����Y� H������ �!�<P�Ҡ��0:C��x�!>U|@�Wo75a%���h������^lY�VN���G�x�$S������O�y�H/;�\�r��ƀ��2�Bh!�0�=�e<!��Q�#�Ŏ=:�#Xi�M5�f�q����^�[�czx�\%��s��K�����!�OY�⁦�9���{$��Jfw#��#B	����"�X9+V��̙r�+�ڥ�I[Y�n/WP��~��C^8���A��`��ߛѤ�d���_3�V<|�������s�V�L��[��K��B�����:��ʊ�����$��H�y�&���Y1ؽ=`�/_w|�/�i��_d�
���g��.�
�OЊz��%�]T���.�DO'Zݑ������������ۯ��D`�*R��K)~Y�Z�6/_>���+�Z>hLT;�����Jb}���ɘ�����U3^ʕ�˽��J��s���H��3�i��%�-)\������+P;#���a��3�a�T1Gj��w/Ƅ�a�T`:��M��vږV�GSئ���x�!4���VK��VB�8�h0��G��nSb���m[�{�6)vǛ�sy�>���P���o~��Ź"���nyz�.���������5{6)�j�4m/��K����S���'J*��(�d�)LG&>�"`�J&���=5�5�a�u
ǹ�c��n.�?�#2U��U�q�.6����^H^^�.�QZ�E�w�5�%���%؂sԴ#C�5��E?�0�
��?�������jjf�z5��>��ޚ����r(��T3�\���4���=����q�xpx/�<\yWL�Q�!KN���ǟ�'���l{�͇錥��wÌ{@'u˚�l7t�T���,M�o���O���˻�����DC�\����*��Aۘ��a[*�Q��X/�I�Y^tW�Y1�����/���K���S�Z�X���'��A5I�ް����ϲ�9�+�� �M�Z9(dU�`-�o�G�b�q^c0�w
�f�bT�d��g���γ��-!kn�����|L|�<��A���bf�8}e��4�g�x��q�y�p��.�+��s��l~��S��!���#�Yj�G�C�ٷ���T��U� ܉QR�VO�����ޘ�_e�����Ucozcobv��8u�a@�I͓��������g��@/r��6u�tAC�o�Ct�)�5Io���6[#�����3�fp�j��%o���P?s>�3��K�1��|�y����B��ѣ{�B�4P�!)�'���� ^�UH~D{�%i���8���7�u�0�"<�0�����5�}�F/���"���޼~�'x;�Me	l��]��Oq�P/�/�������wUX��
�����W�"��6�ݪ��kRE(�w��ϤtC�ͯԮ�j�� �0�� �@��T��^������K���mN�A;�O���^RNl-��ů�I M����Ո��;6��ְ.*�l��p�G`�_D�����!:���TC�V�8ƛP�������h��{�Y�-"��,ڛ$�R����{�\	�&F��v~�?�� :�PGW�[�������$��Z�(��n63���њ ׬��Ơ_&��ǚ��ڳmR�w�2>O�C�r����uR=)zH"{
1\�Q^����GW�|��`ݔ��ĴV�;j���ޝdkq�E.���&�/����Oj5���T3Alr�����7�bL0��߃/��c���!��#�xs����ohM�ѣ�����4����)�D��� z��������o!��(���F�*��������R������A��7��Yk���EIJAE��zt.�{���.�&U��~��8�V��}V?|Y�3��h�*�UO����sz(���)��}+��b�ݮ�b����܆}n��6�˗�����Y�����&�c��I���Z�+ɒ��X���b;Z4|ʝ8SO�%K�8S�~.��yOg�ĊV�,��h����+SOOmgf�d��&Ī���
�U�X���qo�P���\Ȇ���U���1H���	�N���#8|-(H0��x�:�7ka�o��1����M��J���Z���[��iϭ���L.}V��d��`�.�;^�� Qbf�.���*lb~�
�i{<裻T�Ȱ**�4�n���ħ��e���u�Nd!R\>X0.̇L���Zy���(l6���l|z�M-�喙%��|k�O���^�{xz:���ý����U��<b1JկčkF��N7��ܮd���z������"/���1�<��y�k��V<a�za���P�&���(|��(w��,N���׶�7BC�Rd��8�&�����j���kM�f}�:�y�,[l%�~s��8�p�m��3�vM�wƆff�?#� #'����]��k��k�+�p�-���]Ō,����!����Ww'G��y��p�����jRy�^����^m�fXR�6�P5q�^�a � �����5vl�	;�/�����ޞ��w٘y?��Y/`kj��#�O�fY��i#a�	�9Q;|���.*��k�����M?_<V��x8���$���{�sxt ���ꮿ�U���ߪH�M\p���?vn�kih#2>�T���W+[tJ�ռ����w�do��*��[�����r�w�ӈ�����&����f<Y>y��ec�����:���fewnۭ��������?VJB/�=f)��hd��{�>��^����f\�����;|�'.7��hD���Q��}�Rgj{�MC0������~�%����n�L禗��a������xx-���jS7��M��s(M&1�K��ʃ(S������9���������=|�T�!˦(��V���(�RD�`�߇�T�����U�y�7.o�㲋l;:K5�u^��#�ЗE�o*�8~�.塊��B��Ґ��$�����}�1�t� #�2��րҸp����r�	OLGde�Ǭ�-��83��~��<�7}2�q��+������P0�{�e�8�;�F��Y�ǯ���a۳	}�^륆b$�/�]϶ɦ�)I���-~���=��o��h-�����+�Q,C`�r��G�Iǀ �$�T�l�F�/S�<�t
���?�hE�/��b$#�6��=���B�%��Y���9Iih����}�D0�{�7M�ܾ��hD�/���~3I,�y)"y���.��)FD��~<v��a�=���sr�"���i�}{"�6&���?����ǆ�!�YX����7����'[�������>Gk����_�Թe���?)�I��L�(��+�(U��`���7E *�Kr��KF�?���C�{�޽|:���Nœ���m�����3�7Xշt兏M0k���P��4/BoWD�ߍ	�w�=�,a��Al�>5�;�M���J���و��aŋs���������¸�
�Q���� ��!����]ĳ�4M}��7E�����r�p6_�������j�����GG���,��D��$��-׮O�O)��֨5����N�o7!E���q|���>q�,���.�b�y��:�2�:3k���"����[�E��që�����"ҡJ�Hw7�K.H#J(
Jw�ҵ���(]K�H쒒�����<�����s�\s�7ff�
�HJ�R����ac��| e��HQ:�B]^8�?��D��]��Y��W��}����#[7��M�[j�1��Y�Ɓi�����W�+�y�X���&]X�	�t�h��&�����&��
4�c���,��?{5���4*�A��_]'�����'���܉z8V�߭��JnN�2�Ɂ�u'Jc��ذk,=g��5���=.�|���V���2;�d�ݥ�˥�*;pwfZ���x�?����O�K0�ِ�K@�a^�5�EUu�,������)3"ǉ{vv��H~:v8�=��*S�gʋ�|�����u7m���[��J�j����G���?ʅ�iC�X$>�@k��o�&>~��|���/�;z�m�>�ʎ�c����.����a�'\��!�_���^H僨�L�����qȍg'��y�$(M���g�B���'Î|�|y1Vr��X��2��ݹ���4d�vN}�"4vEJGGG��5w6���R�-&��,tQ�d������؃���%a��二A�]�j�vS�dVk�5ޅ��0<#:Ss�" � �Ϻ���޸��JW%����p�y��Xl/�L�z���[��y�D��I)_߅��t�'�{�ˋ)���e���Nzt��>{��Z~[��*���0��mD�/��O�0�\�:�>N�
5J��N�W��ٲ}}�Uv�P1¬��D�N^b�lTI>��5�΃.ʂ�l����_�޸��>_���?=l<�hڙi~��_VVV��2X_^^lKʊ�����§��$7�zo���G��*Ɇ��W��\���֧�g�(I�t�n�:��$�N�f:e�����t���b�7�֎�,K!��,�R2rj��������_�z^CҌ�����{n�;ST�X[Z:P�ظ���<*?�!\�<Ou؎Qt�˞&��p%��:�ZȅQR��v�&
3z����
m�m3�p0-��h�'v?y���N��(��Q��B�:?�moo�`TI�����i������W��4�6� evJ;�-��/}J�ӟ�TL�},y��Bor�_j��1�pE�l,,��sڅӨ�e�}V�N�S��|nݜȿ>����խix�o�Ki��0ɗ/_�y	g|{���˷�)ӻ���U>&VV���w�؟�@�Lps['������ͬ�owx�0�r��keƫ�##�[��=�M�}�v횅�*�V� `j	���n�ф�@B��9𽙹y����y'�;�:Zj����|Y�'1�T윜�X� �����*'_�~]�{b�)��8|K\e�V`Զ��]ˋ���U�Ni��� ���6��E�h{�	�x�
[P�T��fW�s���֎�G���8��ׅ����vhw��j,ߜ��w(��0�����a�c?�ҫ\l\# �'wv~�'´��ύ������K',i��|����͔�롁�p8"8���Ǔ��IwZ�T��{ߩ�e&=J����8�����l�ul���<�n����Qz˹��zѿ�~69E���F��is�!A:1fN��+��z�_i��ȝCZ~!J��]�k
�!���_A��0[6NΊ#<���� ��h��V����r�����%��o�Y�z1�:[H|������߹Ϲ�N����_�S
�1�m���Z'���DAo��__՟���֊���R���~AcR��/!�Ro�z����vG49%�b�������6��..�^��w���!��_Yjv��q>0X�b/��z��;�/�9�V[sz����S�o�_=$ӑe�`���F�ȩ��͛P!�`|�֟/?"X��iK��i�X -fZ����i�i�d��oxSX��/�,R�PO�e�l��_�ҧÃy�u枪�+��ӵ��z����<Q�d[�-7}����M���xЙ�/��?���3K�����X�oPR栧<\댜:K����E��(��҈�_�tM���w����&���4?�'~���#{�m'q6l�ȷ�9�p1L�y���X��V|�3��N+���+m�s�iB�s��W��9�S�e�'�^�^;;I�C)��wI�ƍ7�k�]�)��]Sl2��8��G��-�n�H?
ɾ;����q��i�M1a'@N��,�w��-{����A��M�;�`]�K%���F��.o�~�&*[)�)G�e��B���ڎ���1s%�)��3\�8����q��9���GR�*��=�^�R
�p�aE������,�ɔ�롆=}Glo;��a�`Z����L${>J!�;�2ž�B�@��sإ� ���ޅ��&���ďh����J�[v���^�=n���=�6YW:�� `�~��M�J�a��������͡��$��˒`L��e9��q�� ��52�k��c��H�l��b�c�ձJ�:��}|�H8fP�TT�\z:��y~��m��@i
��c��|YA���~WMc��89shK|����G���E9I(KEl�+�
��X������S׺$�|v���D��[��oi�e`~�y�I����V��S�CN9��#��=֎܆I��KͥjM��.��U���Z�r�=nB.+�Y+�Y��ae@a�A�VI��&9Nhe�[z�*��@�g�`�����c���.��'�1f����u˄��A�7��;�5^�p�\�rz�~<�q�Ҥ����z�%R��C�u�Na(,�6p��3��ڻ`�8��J�[��
�u;Wpo�Y.��fu��y�_p~K��4=�}+�X��t�e�����(�~�1�*ׯ�סr]H����4�H���NE�H4���`����\5&@��tLW�$YT�wW�+�5�Oq/;� t#�����%�>��+�#@��pq�S�=�2�[��n`�u�9u�;�`?�$�,>;Ƿ�k����j�~96a=:|-@��fff�		X�k��n
��}�P�IE�6�SW7�����A����5*;�وw�{_�]�_e��:m��γJ��Y<X"���FW���+�@������� �E&%�Ol���bw��Z��`��9�	�a��wt���Hb�����x���[���g&�(&���v�շn�ǃ�h�x9�a����cC�M虚��ߩ��
/5���	o�5�&!!���:hQ?�G���S��IН�bN!'ĝ�-x�v"ъN��lF������	����>QDbm*8��l���)O��o��:������qE��}��}��4�v�eRR���7��/��Z��<�Ȳ�߮��^���q��A�/K���wD��^Szɗ��2��m�}٥�
ޡ�O�c�my�k؁���-�Pa�r
�	|9T�Tw:r*-,zz�5Oo��&��� <!w�u�V��ŝ����.\�5��K���`Dw��:��0�ȍi����z?��=S�鉺Lז*��NDB�c���y�U�t_�����9,��>+�����$#'#ceb����k�m��=�6�=�y��z�ć0Y��3��\��U�-��?zjVn�!Ӥ�+�����j�*fx.��d���F"��U�}�t�jtzr�3n߈E7���lR�#&�ؚ���i���:m��v�eR-A���`��壶4�s�P4��_��r�t�CWS����n,�"�B���L3}��U/cD8�1��V�TE�y[(�P�c��=W����`�Z��tm_�J;��n�
;j�A�����o��+]��K�!~.H��9�T!3��~ ���,Յ��,[%emh[=�S�ɧ�"L7_��>\+?$�#�Qp� ڃԯ�nﶊ\JB;U��h����>̜"�H\�����a�j�+}EӾ<U����p�;��{�7��>�x������{M �ا����>��)��,�~�`5ڐw�6�T<)`�P�Y�x��h����~����R�7]��N����V\gܕ���C���D�6���^t�H���������ͳyM����"�>�/����Z�$e�ty|�<�p���x�[Z�"�.7*����/�$혭�}�v���L'z�R�]�������̧dM
S�w�u$-�ߪ�Q���}&�����6�y�&�U��"��zV��oZ6wT�Im�_Z�_>.9��jפֿ 0�2Ġmk[�fp�l�Z�ܽ5-�L�;v�N�yHD�R��[�BQ���4>+�=&/e'��>T���y
^�O�ɓ'|�V�b^���^����?؞V��ho����ɳ�k����mg8�z>^�R�:h!iղ�7���� qx劍�5�-�4���6��S��S�m�	�cč}�\��<i����Z7 �(�d�@A�Ѵ��=����0U�iƗv��c���w�w�r2�'�R����m��r�n�D|�����ʮ��0��XΥ��.���g�����|3[ޗ�Zâ��Ƣn���cp����{��Yw'+F�?d
�byU�]����W�s��0T�!���!Zr_�{s���M��)g~g���m����7ˁ���;r��ξ�����rn����� h2Հ0B¼�Rkk뵯�8����0�M�7�g㝤ާ|��+��k�j�#�E�we�Kb�'_h_��o.�w�%�X���(W���B��9{��3���B��>�9?�N�w�)��ju���ˁ��5��J�T��I)����K\��O��6%���&��{Iyv�a�R��}BYI�fu�.�=����b�"U���[n)�2֟6`����^��6k���Raφ�r���Q�Z�2����fr���^�U֔õ�SH���Y�F��/i$� Ú5��*ge����!�������f62_[[�]�ނ�q���C]4Zq��vK��o���j�d�ѭ[��4�e��K��z�A�nW�Z�3��`�D��W�y>�s���s�q	���,���8�y�]�U�v���]׶Mɱ׵|тuiǺ�7[��o[�-x�܊�0+�D� P�)��.vAD"�"TI�j��A.a���]ړ�ʉV�����-�'����O�yŤ�_� ��Oh��m�uIP� �L�S�dLmwЮc"7�M���o���@�,%}C�&	��KB�5Cz�A����K����dya��[�ϊ���:'ѹ�W3# ��v8�B��g�;
�I6@N���U���e�.�<ul�U%/�Dfn�w��Jn�t�iO�5�ԏ��=�3���C�fb*�[H�"^Գ
�p*���U����b��_�j�����e��|��>��]..%��6������Ք��_�㺃��4RO̤"'�U�k?�I��Դ�ٵ)�Z��+�o����-W�n��lF%�Uq�s*+��tq����`�Be@���y��ط7X�=ɢq/�E�~-7խ7\d�6ӆ���Ց�yp�q���on��&5�m2���P�~V/����^i��W��{M1E"�_��)g=)��t#--�c�r����ëf*��O���g���n����p�`�ݸS�h��0z�	h�ML��˅6�7[R����pg�n=_�]6�
숆�e�e"��� �O���]4]��$}�~a���1���r� M�E�`��L�V�����?��?�M�/{�R2��(21�I|!/�D����^����� ��a�rQ�������s���Wp4�A6>��V����,�ہc��`p�g�u_q�r�\�$axQ�Ky��Ԋ�6v�-=m��}v�Oz��=���5T�,E�dk�'���[�$X�S���ö��i�ߩ��"[T��tdq,X'�Jۓ�a���܊�)y���ElI|��4g��|.O��5]*� �8��Y��Ϊ}ї��˭љ����G��G��'��Hq�|˳b�ϳ��WV���\1~���=J�@�S�����~�][����8�K��6��N��\k��k[�����o�=W(����X�ӧO��U��/d�����n<r�[4thӾT3].qPK���\�B���(()sIn���Ȁ��0������%�s��Zyyy�Ua���o9���g����	����W����_�Z�!k5����q�n�ڨ� �����[���u���W�����n�ˬ��j�lؐMt�:�� ���Kk�H�>�BPz.2�������z�����,��U�\?�q�8�m���%x���F�ӡ���w�?kf������.�ĿD'Dd���1�Z�t�~+���xg��h[`n�� �����v[�}��%�4m�ᡏ��`PlB�Ofg�x2���t�XZV]NR�q�Ϟ���d�3���S4�.p����'G�W�^:-���s! ���t��W%�SE.��}��=./25?2�Q���K��N�n]DG������G���If�/��-P�$${��^2�cF�#��W�zg�߇>U>���R�yS>���7�<���])��yt��N�!w�r�H�ф}%ԷMPA�;�̸��BL���VJ{vk�5�)(��G�椔������#��'�@�N�#�E;=܌t�-f��>$ANfOCn�~��	f��+�^�����漠�@���Β1z���@����5(AR9�.(-�{��0v���_����u�8j�fȍ*<{ny���ݛ����g"����z�蓠�iX�Y��f�%R)�����O���tl�d#�ә6��UI-�{��I���|nk�a4����ZC���ށ@5�1IC��fD�����2Z��|�ea��8b#W��c��t��ւ���kQbn�Uv�����{���@�-33O��>�g�1�jQ<Z��$;��˿~�*8�.)b�sȨ�Y"�S�wu�:F��e���"��}7|-.�LT;B���ˬ.�����h���1g����i3��HM㽣�m�tR�w��<ep�:���,�x��?�����_��g�^ �`�t�����e ���\���k&�Ӑs�/�-�P��Yk�h��1;�~KX�1�|>QR�Q;�:?1�k�"��g�r!$.�T�H�[�Q�{�eA��i�x�D�@���z�A��_ouP�.�5�\�{S�';��B����>l<���-�	�[_���+6�;u�^R�@�@��O��`�|��|����@�˰Z��x7��@��Gw�y����*�9yQ�Z���?�,�U���ҺˋW����
]f�]JKҖyL���⋫YL.?+h����?,��ǫuAU���B�5��_�~�i�L8�\{��S^r�J2�p�t�{3�?,nb�]��^�6t΋P.���6F���;R��7X&onU�5Mg1(`vL~�C�r��Pd�c\�G��l�Z!����-.�����K_*�n����,G�I
n�>G�CNm���Z�i�xɧ�EJ�����?��	]ٱ�T�E���$&����k�G�ܝ_|�6�G��O��\�r���@�)�ǩ <sGW&]Z��Fm�e���mN�GuzDN���/���sj�5tɏ�G窮߬�m>��[�DSj�?~�:�^��L���^��I]�b\z��IM����"��Aq���ܿ�������Y�䭉�ܛʕ �0&�1�@]V��"���{j Y����ɢ���/����v'	W��mVhX��{v�K� �.p�MfK踔
�]�i�UՋ����(TTn{�E
���NJ�܅Bn��<�U�]���H���E�a��$P��v����<+J��Հ�v	0�T�����*l�!�*��eK��c��Ա-��K� �(��o4ʻ�~)�Q����_�\���)uxE�B��5'~o�����w�yY+q����i��kö���ㅡ��ޚ�ǲ��f��0�<��m^#^�kH��B�H�9b�n޴ MX����&���$$Wi�K�l��j@���e����I�%c����� 5��S� �gU5�Ѽ:`�.����3���[_����K�q��g;Ӵ[����l�hv���v�ɛ���j�>����>W)��6/�_�/S^�.����]��	¸�棉�W����l�{)g�a ��S������V*��U�+�h�@���Vڀ��j���\�x��8,��T����7g�@�A��=���PCq�w�S�a�����]�
�u�W�HX�"!!a�^y6м=JGGS3�7��[����LJz�h������ �o\\���J�3燴�b���V]I8_���X3�تD�ճR��o)P5����ܴ�^U�` �%�ɮ]��3���˓Cn�����Ȩ(������3!$Z7��.D��×�C����0�r7�)ĕ��Ă^���1��\u��������r��*���U���s�|Rj:�l�В>g +�������cg|�H�n��>u�����-4����0�y0�C�O����\yV��l�y)6�0QS.互��:���)IÔ�G���)%Xo-t�UXG &rIn
䦦6᬴�
�Qm������X�&���?c0N�y[(t�1�}1tW𭼬l����+����ܷ,�FJ$ �G�:���ˎuBIƾ�>�G�?U��)6ƍ����EvHΰ��W��*�5��i<J�R�����k��;���\��A~�zl�Q��Q)r�e4�X%������Ƕ��T=��Fg; �--�����Cհjjj���=���י���?��C�ޘi��ݾ��/�@S+�k�V�(��3�|�|{_��N�9=��掛�N� �_��K�����
W�{�񌄆O6Iy��N���j*����z۱�8���������ҍ*�Ǡ'0�V\PLz�_?"~�1쬢��'G��W~J]�5�8J;�6{R�Qc��=�;v>H]�4�k[�0@4�}�����g?���_��;K*�����'�:��氧@6q�(+챻���I���o4��Q� v�w��r6ڗ!SJ�ϗ�ѨT��v`M�U����|*���-=#����.$����#��G �4FFDd0+D/M�McbL|򎎼PLi���[sma��ט"cc��� �TS[C(��ܦ���t_b�� �vZ<��2��%����e`)`aH�B3=��Rml�s=x�AD��k`_�5�c@G ���i��-�D���� q�?p%n��S�6���Օ h@��:�҈agy�Ge���AὁU��qG�NNe��Sg�E��)��FxY�mmzz�'����R��:������x����)))=:+.�C`މ�< ������Qg�Z�
G #���@��ԁ�ȳK~%�P�W�b�[�I�O٨a�"����W�١_j�q�O�/����F�c>�v2:�A�C��4ɠ��b��θ���
!��e�v4p��9/�Qd[�8;����_N5�gY����hfFt�W>Y[	�9�s��;ڐ�(z��/��9��WGO8����W�1�YN5� `u<<jCċ>��j��¡E8��mm
�_ZZ�
����6����i����������6�5�����_z��V�z)u�F�$a>���7f��ox����lGF���>0l��;wt�r4���_,sc�XvNNMe���V��2���Ӂv��
��~��4��۷/�@]q�H��f�=x�N|���G��r���5���u1o��l��!��3���̷�&/'���F�����(aY�ޕ�^�
HLC[�Ѳ,�Θ蘘�acO����ٖ�B�^�h�!�oWT+��S��P�C	_��r�g�v�Zn�$�ф�g��Q��ޣrm�t�8n666y��R�6� �Ɓ���j�~%�zk�����P���>vc�%^̻ZOr��.9�[�����j�/$@���sߢ������U�T:�ICSg	���px>�^7%C�:�\��]\o��Z��|�-+�࢞����-��"�sT�sH��ѱ��QAL���	�� �5�Ճ�r!$��`�Y�){y}�f��:ĥ��b��X8�!}�����>�T�ٹ�w��&���eeDͨ�U`����s�픜:�$$^1S����G%��a@db��889v����Ǜ<;�&ȥ�[);��pL~���4y
��q�P�/@/ �{�O?C��A��gjw-����b*�uG�?.pi��]j<���s��Ą\��ý"�W�@��5��ȁ�X���� �]�o1f�4����G�W����/8����t��BjA�s@� �<ɣ� (MD~!�ɵ�nî/�e@Qp�-cQNܐkl��p�*�M��d)P�tR'GGg�$�|b߰7�A[}9��m*m&U]��s�tdq��b�oV8:�A���\w0:B��*�T��_�؜���.���*.=�Ĵb���:ĤФs�(�@*D��|�1`��_*�!��I��� ����x��QX�}�`��1=Xh����OL�b�b�+e dg�+���sH(�7��5���\PZf�,p��0wk�ew¤e�;��S=��ꔁ(X��3�Zr��6A.G���}	 B�D)�]�)�c�h��D���}b����z��[YY���������$b��m"�E��4{���O�8��`I���2^f�HR�I�}/p��h{�b�%^bI��}�'����Ya�(ihҿ�ؠ���q�Ei�9`���]��+��iy{+�
Ï�4&j�I7̀ 合�����7Q���n������L|����1�J�;hl{(,B�4 ��W�*��Ł�����W���ͤ�	̺��Y�oެ���}k�[8�����.~��_7�"|�	�=�)h��F�2�����ݭ�.K��NGG��_��@ݘ�e|\ �}���Wn-��;� ����ii��a����Џ��I�VY�	��u�LMMㅐ��I=};u����פb�����՘��솄�f�2����ޕ���MN}��W��KK�4SPP;ߝ��j���%)�/R���殬�$��'uk���H��u�DH�`�e���8'K ����l�H��p�#����:����+Ρ �C�Nq`�����R��Id����?rΖ�����T�`��� ��S����
ѶU���U�{����=!W��S����7Y�x�ʒ޼��A�)ݘ��)��D���(���\�>�v��uЈIE��Y�%�1*�Y�A�I���0M�U�H� `�zv@�h�4n߈'�ر�`J4�����Ú��0��5��>d��5_�%S���a�|�ü��BɎ�Aa��ci.�*�E+���vc�Pm�7�7�n�0���q������*m��,b����� ��Pe4_�B?�K@�Φ��\�.��f�@o*�[��#��N�K��O�����{��Z��9>��ޗ �������Iկs-�9����J�6��o��(�P:�|���G���Icզ�������R�P���G�<��c&���КX�k�q4��ePUй��[ z�l�0��n�i8¤�U��/K��MLlM�=!J���S�L��f��j���l��b̮JHH@�M{�@[�\WFL���Bߩ{��/�ɭ�#�W��z���}`I�Pbu����x%�n�����uc
? ءeh� YŔ�@a�b��AǍ!>���#��`؂&e�H��VSSˮLHI)ޛ�T�Z�m4�5�ʳT���E��-�����Vn���>��bn�|��u�Qfd�L�i

m�6,��~D�����U��V��r>�I.��{��i@��%Ǳ�C~~�rˮ~������m�3ߺ�Oy7��IQe���i��X�[^II��E��5g�$8�hw}���ƞ �c�4B����ǃ���:��x�KB^�I�0���g��"����^轱>=�V�+#�0EFu��0�>h���W�H �� z���t®P���]лZ ]�-�,~�%�� 帠��/"�l�7=�Dm�[����W¡�~��;��� U�CA�.� P�c�|��(^@Yݩ�)�W�57B{@'m�/��_�<��x��(ӛ �c�)nL ���j..֫ddK}2���c��q��{L:���H��	C�-��m�m���@�eWX�ˑ����H0�Re�|E߃۽y��;��_�Ǝ����T�����$r����Bƈ���Q�h�pwu ���	Cw�~��o��x�{o҂b�'&>>� Q�5q�B�3D�c�fk"%FU�� 4m;,�d`���;�GN���R�sP (����{-s�o^ 2�ɱS�n�x��6�(�ōSs �xa�l��s`�����+�n�[)!`�}��Z����eO~� 
-�-��
�i�����Uߣ��5�>07^�����M�u��h��"�l©�g&�7�\��-�b,הPw��e��8>�ڏ�hY����%�
��o�$ǿ���1Ar��q�H��X��_��XC��G�P���Q�XE�"��(���n��%5��K��$7�?=~�e��Pql%�����S7�����e���P� ��1��ș��:�^T�{�c_3M��t�F뷮D���չ\�F)v�Ф�3�+A�n�$����7�5����4�V���M�Ƈ�iz�0C��Q�������3�o\&"z���٩�J}�$��P�8�`��@��P��kee��7AyZ!�+�
L%=���v�*U����	3�������� ;�0x��;�XZ����V��~����s����@��؟�d�M��)�j���]t������n�X<7D�_g���k#<�Q�K�C��!��R��"�o�p ��O�}�u^(>���uE���]�,$�awn>�>{���
��ZY�eff�SI��N��\�jI��k���o/�"���a߿�fee��Á�S��d�"e�v���$���6!�0��^fe�М����U;f �+NL�b��۷|�u����$/ {�V�x`����g��A��^J��Q��:
%��9�-Sh�h,J�@���&�XЁ4|V/����Ԩ	Y%xNμ_�RF�&���N�z,*e�$=��n692R�UF�4:��;;;�?���OƟ'z����*��T���:C��r�������|�͠��Jgg���4��e%�U�&KM�W��<#c}~��q��,�5��»�=��\�Fo�d��O�䍌���Ԟ,+Yۃl�ݲ�%8�rP9�r��@����g{���N9�6L�#�w���~�zY>�I���q�@r�1I[M�"����H`�zR�� ��
�aCxX'_:^?=)�ձ=��l��|��}��X��I7��=H��
�9�&� >?���R������7rsY��7"�)�Y%�ť-&���_�l���0#��(h�#$$�}�	<r� 1i���?�v���dٝ�gS\���vr���Z~���Ĺ=��n��l��R�עw��6����S�G@�����Y(t%� � ��5�Ҧ=���0�ݫ	�n=Up�m=Wϒ���Y��u���±�-?����>I�#��1�f�U)>r �2B�E�����3g�����ٍU@JlU)��M"c�k�n�CV�&ǜnv{�\7�F�Ɔ#
�J��k�Ҥ�=h|��#��:"{�ǋHi�B8~��� h-�`����0 �0GUϼ���(Ƴ�[s�A�!؂_�e�Oy,�~�}�~�ڵ(E�ڭ��{�s��E`�T�>G������d������x�J�?� 9����`K�=Pd$�=%�8 ���C�ϯoɓ5������3K$F%h3�BT��;������da�X�?�������@���[w3�~Ӹ�ً~}9)�Hȥ:�NFA��H2X���� �gN��D���
����=v��Г��_*��h�g��zNP��1:���,��E\(�XF7@ˀ�9���6r5��Cz�ͥ��m���ύ�6n�b��M�U�+$�~�:��5�anXeM�x��� ��l�.t�_1T��}��b�*�x��w��3�I+��ҝz�5���ɞ�T]>`0Eyt(-�Y��d`�3�V��SK�~�j����VJ6�v����g�I���,L$�!	��hC�߭��B���q[���1�wo߲U�n̶�F�s�tհ��}V#�������
F��mʽ��{�w_*�{7��ϟ"�Y+�3�B�!B�Y5�V�{��K���9�,��)���=��&������|�dӭ�Ɛ�~!(�(��]%���h�"���o�3&�����a����Z�ZI�NQ�-VR	76q��T��}|઩Ke��-m� ��Y�j��E%�6���B��@9��4)<p�|�}���H���d�
�3�322���R���u�b$��DA��a�(�ЬT���;�����{T�]����GTQm��3 P�q�����C>�����UH��*[��z���O��*������y���Z����9�y� �F�_�,�������������=��Ȥ$l�G�]��ͽv�j��.�+�La�NM��7�ݩ�ײ���_����'X]�Yդ��g8�����&�i-��s���� �@���ERRRN�
ٕr]λBu��Z����r\����(��x�j�n�i��|����Ōʌ�%�iVNΧ��T;��7o.��T��j��ȹ�����\� �E<��ݵI��O�>9��D.�R�4�L�0D�l�{��m��R&Ӯ�{K�啯�ff�vWC�4�e��DYY/ݻw�w�n٥'����;���żهh�}���(t%�}�~�wt�TB�6��R�t�R
1ښ�O�\d�OEC�DM�T;�oǸ�Ì��`z���n5]b�G/�ŊT���B}��}����JNa���	��!���-y<s�N�0�L�� (O~��rg��rw%Nל���P�5��V,o-O��N滬,s^��+��ȫ=$�
7mJ�}����J-:(���u9m�*�wo���%��զD��%���0��0"��cE��+'������`����:�<J��U���z�Le{�C?�{��T)]��
� ذ�� R��77�bb(צ�2���DH%*�;8:B�}Uv�_�%H���ƵB4s�O�8%W��X�
�***###�pa�?%������767��hAZ:���;222F��qEEb��v������>�@T Y�ZVV64J
�哶��q�T/m=��&j������?��l��������o<9P��u�ɮ�� 1��cߞ�/��C�,���t#�O���隙�Y/�����Mf�4�%�
d_����o�#����@�<��A�M��HΧ)ua�n�ȶ�(S⇾'"�|�ZY�:�:/t���:��n7���o<od���w��9����i_�jGY����0!}8��"�:��J2tA��h��t���e�v��z� n��g�_u�l�u9kw��.-�i@�����f��)6�����dT�BDD���~�Eш��(�֗���s�����ۼ/�i������RS��i���tk��Ci=ٟ�-Q񴦦ffk��]���]BB���=ZZ������ڷ�����YYY�
Y�?o"�����EK 	��/I�n�C\����?�\}z�i�7�u��]���v�q::: ���(���$�-�P�N�e/J���6�~P3�N��
J�Te_����^��m�{^����?����NIk�j7Y��YO����^��@??�ׯ_����Կ�#���f��x�m����ϯ[�� �vYRF.��$ic��ޝQe<I<��X����$�o?]�w�`0�����Y`ַ8�GLTߊ�!����ݭ<��tSlx�g��g��m F������6j��\[���B��Ô���_Xc2�JK��_8�O����˓�HT\ ���˫P@CC�ӨVW�c��>A��'��������LS_�\�1�fD�N�5xK�Ҿ"rnk��U%YpAR��BW��ͼ����Gf�w���[[[���A%%��� !�Y覒_�sp�m+�o��Q��%�#�lc�9VԳJ3��cw���b��7/�i�������o�h���u~>����k��=.�l��g����4��AFvǀY�{`��G�<T��$��re���+m�{�$	&�=u~�ܼysȉ�6��/�zke�Tr�c?��k0m���5jj=ԇχj.G�K����w�R�g�;}�{W#�h��p����"���j%�f������P���8�޾blAYY�W@��mq��5bW��v��^׷3��8�BE$##F(������k7o����lR�o�,��[�-�$F�X����TA&#!���)��H�7 ��?x��А�������fSV�-½��JJ$1<&�@�2'ρ�X�M��6iPt�Ȟ��ݒYz���v�w%�Yi�v�ܵ�J��(T\\����7%憪�*n�ϗ@��.2^JG���v�=���ަ2E�-t3f��p/���V�@V6��o/��b`<�Ч~����'���9Go��MVv�'��x���K%pc,���A�����%�^4��_&"���GE�& `��C�����_�eHz�$V��~��0����G�	���"���,�^�ƃ�]|����J�$� b�#�m���,�;,,��cT��m0���j��y��S����$��nkM]]$h���?ctB.M�N
������S==j���Z��ߴ�{�A ��<��M��\>��u(o��]�_�6S	�jj>L'��8�@���@�SJkhܠ�6|H��F���Smmi0�K�������z�=�J����٩���Q�a����ݫ
��d�BB�W���5[>Qr7MM��g2n�9FzZ��?�(��W�ۏ� �S����������� Oc:�%Ց?��������{�~�������g��(�u9U�('9"��}cc�� ��h�$���[���k���������[?\����'�6#�S��gڰ���t
|�u�wu|zy��"��j���P:<y"��Ռw�F�X?�>is#0���+��A�s}��D�6���S,e��w׍b�D�/�v��s^yU�?���k4�����t�o������l�1@�'��Pm�W@�]�E�l���f��c�v-��5��ǫ����B����+x���k�H�a	��R_����M�����@�k+6Ȃ+&>T���J <�9xr�������JX%��E�NO�5����xa�����K��$7f FV��ZS?1����ݜ�8?ߟ�������W�"}�Q�ٍ][��ȏ����^��{P��X%�?6?�]1E���EO�bAAA������?��rկ�lv��5�3��s��|�p3(8��'�U�Y��k��4%��Er�2���Z.�>�c���� �[�64TT3�Y
%UU�V" yK��_���Y��1�3c��mEFN�V���y�cT��0�Y!ũ��1�DG0�����i�B iL�m�{B3���}�RdLw��_ ��V2��@� 0� F|��hy�G0��Ȳ�۫E�>��g|3���%)kk�BW��?sa|RRWO'����~ƯB`$h�΋�q��,�Օ'�o� �ձ@*V�?��+w���p�����[@Um�ߠHHw���R� ݍt)� ���%����]"���:���?�1p8���s���߳�Z�8��;���~�����E�Wj�����_�' �@�(	������D+z�y��yP���E�G;��a�⣫{Ti6ƂG`�@ �L��5bTR���T��=�\��h��	�ۣ"��q5�_�̀k&��RMkl�q��2o	
��jY���JBD��Sr��A�EAMd�����~cQ���w�C��x���=���|-��JAM�?����x�'����x�1���DW:��{JJ���WG�2���Θ���S��Jw��T�ˬ�����]�C�ؑ!��\�J¢�HQQ�gwc-��oҭ!���I��I7z�{�pA��T�\[Dw��vT˵iUG׼�ih|��P�����#�n�#}�+�l"!�f��r�e᭵+�C�6z�r	��ZZZ?��Q��������ZZ"��ۻ=�h�4'!�u�w>^A�>TVS�|�ĴYoc�����]�UF���TfJ�����h�4�y���/�:��t�@>Ae��*����`��o�����J�3* �������P��|��xc�B�i�^�-�b��*YtƘ?^E�
FrZ/I|x�tZ�Ӧ��i��+9zc;+��bw���f&I�w�t�>=���d9��6m�FC���˩�$Cp����O��0�JCCcw���䣛h�w�\�z�>w)�{>,�h=)"1��kqo5� 7 �:|�=�kE�흝����Ud��ѽ���l�?�Q_���1ˇ=��0C���﨨`����+�II�+�*(�*�s!�
��.�M̙�V�	��<�
h�f�Ml�d� )��Y`79����y�� ����1q�Y�V}��r�d��^�S#�ό>�>�� %Ė(`Ԣ��DsX��ƛ�W�A:㸪N
ο�xp���'�U.'@�F`|��#kګ��(��՘�d�ɫ���S��>�(���BB<��/>P���˞�$fګ����������R����D44.9���`��6{B01tl����ۤ�!�P�9Q>�B��!��c�/ͫ��o,�˱x�I2���:׎�/�~�l�e<33�����?G-�z�>55���'��hr��ܾ�����; �/ԘFu��*�u.6>/�.�0{�n��%088>>��C�F̀�S�ȍW��QIf� k���k���6��3�\�;����ks �!�^�̌��������e)j(�q�}`rT�;nè���{�T1�)2T�?ܟO"|Z6�a��pԹ��E+"��7��|����i�����6�~�]D�;���)l_����ҎcbcSڽ#+.��2j៘VLߙ��"�����̫`���Aq }�
�����!�iv���g@�-(�<|�A��\E#11�-*�,x� x�~ȃ>�<i��y�a��s?Gt%�S�ot��<YoK�]�����r�m�X��):ݥ�XS��P+���@���x��쳇G�¼![
�-�ut(�>��`2�hw�O�W�2����~8�It߰X7��O��4"�r��X�:sx��%�=�8:r@8��P#�������.��-��B����>��y�gZlG ��^^^ss�5��dQ'�����Y����e����}�j�D2����]�Bi��v/Ϟ���Q�%���?>�����l��Ϲ���>�-����et�?��g&&��:�$�0ԓ�F?�t�O�Z���b���l�4��z�֝-..�6s�����Ee����ޞ$��'�.�H<$�ϟs-�PG��E�����>=�����k6�Z*`Q�C�ն�7�F�!��� �{�3�'''K`P	��\XK�A�Ε�)���!�,k��_���1-��uxn��RjD@/h������}y�J(�)��!�H��ˢ����|sn�1�r�1�0�H���F{S���666@��!��ᙞ��+R*��ɡ�^�(���3==�����	����H,K�IG�<��ay�˓O�?�B\(���
#s�\����x@A�1�)H*$$dE�h/4�S�
�-)�,T��Z�(���턟�>�2%���C���>��@�;d�MY4�N��o�4�,(� `q/綩��'ƅ����5Mܵ�D�@L�j�YX���=�8*�6�	ҍ��ڪT�'&&fb~>ip%Sлo�����G~���̄��?"bbo����Bvց��v�-������z�	����k p)zad�}��ۼ�Ç��I�f����ntz'����g �KIII��˧�?����&L�.�L鲮�Ή,�_[S����3&.�ݵ#���UI���K�֡ȩ�7F6444dr�-V3Y��-����uZo����l��1�ME$����b>����ޞx��K�A��ҢKpJ+�1��UύgddTV�j���^���i�R��%��i.��UPPn�&*����C$����J�Ņ���F{ӔQ��>d_��5nz����>��y@�	HO�Y���C�o@�Q]����}ߨF�T�݈h�]����q_���ה^&��G��&���̗ޕ=}��Cimm"Xd�����U��YB��xwI����]N��o=��3��G�ZZ���LÊ��<2*�"G��H����k�)���(HU����_�aʎ�럪n���8��n�<$b��N�ׁ8�>�&{4t���*<M�t�V���4��l,6�̕2+-�I�^^`�u��V��������m��4637�TYUuw?�Tgy�w��/�ʥ�T���������eiϐ�	:b7I�4����I����S�����i��#�?�$-0D��}{HHH lg�4W3�K5���;(�%��wߕ��
B0��֦x����5�
�]J��AV(V�OhM���Q����1�V0ݣP ~��l����א��܏T�ǯ�j�*l���7��Ks|���*�g��Uξ�{x�z�Tf��ZB���nV.�X�����j|��R���ڰú�����0��,cR3����~�_�r+���k�-���!�u>��|��4\í��H��'�QNGK
��1fܠ��9��!U��iֽ}�9�]���h_��v!�Xn��P�a�����u�)��/������k�ڵ��Fi�D�N�֤�z�S5-�.f8��h��B�Q`nDU��?�c.q��࿆C�T�[�Z�~cSk9�B*�O��������X����������]�KYK�O���N�e`�۩V�?�܀:P�2�֨� t�n�����r����4zI�4Q{�����}�A�M;+�)����ϴ4-�u ��^Y_��dbe��I�0W����	�����HAA�-@��npjsū���#9baf��fC����5w�A�1���åxp2�/֠Z���ʪl��U�0���i�lmn��x\}�_��w�)T�Jz����$��UNiYd�N��Tlʑ^�v�g�=|Wᇌ��8�8{@7�>�nw������T;�h����I�(?8ԿA�^h��j��8�s^��::�ٕ���bK�T!;11��M�������f�x��_���epy�g���
2�MY�𸪹V,�C<�kO@Kb�zt!�s�)UZ���B��GL���֝����&�����~�r�"@��e��ii�щ��{k�iiޞ�;Jt���.,(Wfgg!s�!���x��YGۣi��"h�
VV���Y�7/˱�iu,,@������>u��	dFez?�7;϶������- ���oY2_�zh��(7"���'AŤ���e�*.��[.��<V��e�
>ъ�uuu�3�_��.cd5�n7��ڹ�my��u���)qm1�t2
S#�1�������]ԫo(��b���6��b���f��(;K�飦��?6�y{w�40���vQ��%R�Z�b����|co/4�٥A��/r�<<<!Oyoow��d������Q#U�����w�K�i�11k�F����v"
W�N�	'���4k/���w�l��l��E�H�G3ۥ��4�dee�F߳� �,�2��R<|���^7��c�d�?�4BG''�� Oec6]�~Q��0��!��,7F���v^A��SJ����D6Ye�S_��Dֳ�;����m�e�dWT0G�133*G�i���6x�gy'2q�q{&�~T���������˷Z^SS384�GSS���n���ګ��
ب�8�d��1p��i&֚-	r�S�&&� '���^Ů�+ٻ��:q�Z���66D��@�+z�2Vj�o
�^i�zz�{�,�4�|Xd��Wa���Y�wԨ4���h�{y����>�<�@����H
'�[���şO�t��:'�7����S+��x$c��������SJ뗵.�*����z�o�?��0����z���7gz����U����%c����������5ɗ����U,A(u�.aO���Oη���MQVUT٬�M1�����l��b\0�c�+ �Ev�����u���Y��z��5�!}<x$���6��U�mNG�FF�uWG˸�G�Yf�A�~ ��h�f�^OWj�'~nnn���zӝ�@�KHA������Mm
@@p��������~��_V@dhM����@U�>A����j�A����J'4����"��ycT��d��G��@T׀ς�3otL��~oK��\��������k�mG�J}>��Uz������c�4�,2�����Ye���D��s��$R�+N��P!;��޿�8���eK��K6�G4�+>�����B�y�=#���FH��usRE,u��
����¸V��XT<��ot���] ��3K�{��3�s�����
���o��:2�]GAA�;�HQE�X�zZZr66��{W����6 �z�b���_���Y��os?=��^���;��i�7;��U���j�|EOFs�u��ok�����}}�֝����P^L��X��ShȬ�'g�hW���\�j���:.�n������%06�{��1�?�I����N���3�#++Y��*��RR�srs�U�Ճ��Ѫ���Ry�������?�Le�p}dxR;46��],�(�,?�ś�V>Bդ����e޺�g��P��e�!?��ђ`�^�������r��A�]��U���8e�qk��!�0��V�)(��@Q�,,h			��'��l'IcR�gS�:jvHBA;�����~Y��5T�7�k[چ������C�񉚩>431�;u-<��gl)M��4vj���,����Ic���/�\'�se����|t 3|��O~tosx��psڮ1�Ð߀�P����{��`2Gl`�������1t�V�\�_����Zf�鴸�����V֔��e���	����Aqqq�A7,�uoo�+#""���$�'���T%��}�1۷��;�qW�gI��Vw�$f�> ������V�jj�P �v��A�@�+���K��ӽ��@�_��%t�Jnn�(����m.֘�a�������7�D��>���#w�$�����nt\��,�fCTr?i*��A� ��j����Y�9���2�*�4Nd��VE7W)�Aa'�@EGG���$&���E�{@�yw��)��lE,��"�(�<j@�p�b.�g�'&س׼͙u�/}$�����'W�}�gt����IU�u"y�~��`����n�䥦����ٙ��Y��#�G�4�X;[cP"�wo����`�Q���d]�)�������:��n��E����@ر���(L���[�w�w�K�g��!WZr"3q�wB��@A��԰xܒ�'7~ۮCJ��:4��v��x�Gss�ں��*#q���A[��
�o���gר]d�G�"$�7-�k� ����l��� ����P�������b\�l,�3�щ�#<�<�ţH:q�F����q;�+�J�x�f�ǁ��C�x��;22�s�"d�O�;c�g:�`�2�v���a�|���yI�^�ߐ����G�]k�mkkSߤ��������L���~�^�|Q�;-j(ec�q�+<yGAQ�Y�Z�ŭ�^�`����BI�K��nw����.o���𡆣����6���|@��������|�jrN����?� �o�읎�誨���}#pa����Л+�^��sl��2.?CF��q���hN���-91v��|eο�c��QЯa%0I�>�0j��Iq(ܟ��GD�������-��3���ᨏn��鼎�^���@9��)��@6� /�"g3I���ǻ�N���~p���!�< �DEE�c)�B��`�##��Q��D�#8����O���o��r�36E����d.��G���G7�զJv}�˓e��S1ss1��sN��'~�(����a�<O�w�[�����Tn�j�����j#������o/"!a�(�(ȶhPݎ����6ւ�;�K���Փ���#y�"��o��Qy̙3��*�ݚ�e��.�j[gg;I��N�MR`lKuБsp���ɕ�{��l�y��Y�%�������ׇt������xZ%��_���q11��qT#ɬlҿ_���v���^�n�r��>P���q\K+���VZ-��ZQÿm�f�a��V��H
��,���!���IT�Q��
W#��I�Aaa��mQ>k���\���m*��t��mJJ�7��Ly|H9!�����5�ø�U����:���]����k����a�f��c
��9��k��F2�ZrP����܏N���}d�w��O����];��z�B���L�K�����;�>ͺD����Ot8!���7�8c(�).Z�JB
�b�A?͗�2ץ��ͮk�����0�"��E�h�p<�l����B�g��~�+T�����v<�3$�F����fa5�wqq���ni!��Yvp�p}�� 6�wpPR�0)��qV#)����J&
���ۜ뚈��v���=���rh�,bvv,nׇ����-'��l�h���6��c���	���J��Lҥz[ԏ���k ����� ��L�����$������%$$�*�~ش�]a48GDF�ż��\n�fT��������p�t��`���'O�������a^��t�,[�,'��)L.d$i��A��LO�%��<\o�3#}�ښ�N ^J�Y�I��泂d����8.���s2�w�����3K�K�8�b't�� :E]��2��u�~�<7�Ԏ��������u��C���	�Cb���OMq�d:zoS&��u0�1��r=�-+�U-.�Sx3�qͬ�o�m;����|�8�6�Ѹܜ�W�����::Į���[� Ƅ�r\(A���� ���`�����6�A}=51��		)++
%�����!!!4̸^�n" d?��h?|��UPyYP��́��42�d�AAF ���v?�~�}� "�W��coK���������5G'�ժ�fٍ��y����NT"w'ϻ毜�p�L"@�mq�U-�T� �ZꛂI�h�f��e��|餉z[��>$BN$j�����^X%�P5�����奄�
�la�V}��1��+�\�/c@:���p&m�m{�p=9=� "�\�At�ã���Mqs����z��gmm������
�CCC����SS#qQT¹]��p��Ƥ&��h)����	m22�2��_�����Q�g��I6}���Y�n���P�aB���?^���*]�ģ@�-�~d���[	�_�IM,��ܥ�5C����O��f6��"S2���6�xA����F�7�$rv��^�
��$8�ds-�5&��a�����y�I����Z�+g�j���G�咒�;���Cͧ�o��V���G���	�m��Q��W>m��/O\($�4s�݆����X����὆�%jvy�۠O��6�M�"��	,�ZkjQȤ��o�G��'�����pL�-�6E�|�?W�;�w��z<Q��;�L����Byҡ�s���ȍ�j�8����4Pw4\\8 9CFǫ�A���^IyA86��'�6�����7���O#[q姉��Y�s���k����,�Ki�@D��b��xvv�����'׵����Û<n�B�������	Vp>	�j��:{�ee+�ˈaR��2��N�����~�ˋ/�q�?��"
'\$�rb<��,(-岣�	��{��K�plzUp�3xTT\U#��$ph���|�<l���C�U{���zҦ�m�ؒ8����*f����-ꥮ�,�����%C���1��t�S�����58�+~03/6���'�y{^S�x�|��r���v�������頡�r��&�v�hK;O7ޙ��xx�@��1	��G0����!:F Q]���LX��MT��~/�8��^��}̡J�A�9�p�{�kO/3-�`�x�y�s�����r=j�G˵�ÉB���]����]k�-�̀1Ê�8~~s��&�:aLGKI�;N[uk}����?�͊��v����"i�����B �S�)�.�����RF\���l��T�����P-T�j٫�т���<z�R�%qII�\?w)���S��6��z�唱�N��i�A�Lm�3�V�{��c�6�<�%� h�� ����?����	�014���ڀ����

�##�h@���v�u�P�\��q��'S/-g���7|��).�6bS�t}}3���`��8k9fO/]�vj�UUsjk�^á��W �
i���H�����>�X/�vn��u�%F<���d#�K���ҩqNS����G��S�b�뮧��	1%m.9��呰oäb3�l3QI:����+JJ�[/S}߰}']�yLf�[jgKD:0������#��6cB�(�Տ@�$�)!�I�5^ҵ\~�<��wK�7;�}��߷���F^��3Վs�=J8dφ�ĠQ-�4���%��j�+@���𷢢b���ٞ#���K���`��(��n���sZ}d��x��j�@`���ѯ�8vB ��U�p>av69�l�{k3Qb3=rz#jh�	b��O����i�xv� jǣ��7��T�����#م�'ce���~yjERy��Ừ?���\yc Yڸ=ی��wqg���Z�Wt
rh0�HWu�fYoD^[���ѭ %� -E�޾c�BA��w�\ʮq��?��J�E��!&Q]�bˁ���O�a���MgfU�zn��rKK���	��� �	}�D�8;�L��(l��Eޞ��� ?�񫄶{�"�c��y��P���N����!�>�� ��sb�ο3�ѕD�i��P��Ϯ�s����k�:o���:���7���ط=���U+hh\��Xx0U���R~�.H�w�9��7v���-§S������CX[9,��/���ձ�*��:�]ypV�_Z���kkN��l������`p0�RY�w����4������M���ǳ���M~u�[�ޯcw;54|��		�k�j{Ys~�^��/���~s\v��:Y��7g_5���GS�n��憰cu��8�C;s���X��'i�v��d�=۬�)*f��+vrr�U^��ɯрґ�^�K�X�	�he����MEQ�����<8���$M�̡�j2F޺Z�� ���9�ןZ��Q�,���{ݾ%�_���:�6��rz��T�"���٬N����\��o
ǧ��E �%�c��M���yXLrl@��^���'!��WTf��l�6Ũ���)�Sڤ�t��Z:J~��-����-�S��Ee&BF;���"�L*��CH������>��Bc`��%E��ߤ���ז-O$�fa	�{r��w�t�����񭄁Gu�[��ViqE����r*b׿��@ͧG �#�u�H�q�����5B��C�WQ�_4\ר �����V�����:�]9�y^B�°��߱�g�ټ|y���~�~~r���A�ep�7��4z��/R��!�V����9A�=���2ջH��ޏ'��#�QUU�����h�=���N����s��0���'��m��n�}GW�U��3��Z���J+'�����lu�kZ{�n�",�<>>�h1Տ��Bp���T_T\\)�@����!q�ԗ~c��Cc�'�j.��@�\m.�̵>�?�3	�g	�Tx��u�@e$���˂0�&��y����M>r߮�q.&��Y���i�c�/O�ԅ?/o��VxV�㏿��T�K��3�$GK�E���j���ş���QnN�9����44�1f�b6���]�f8k��,���t�����7�h��".<Yu�<�H��[���[�����.WT	��Vd����Ҙ+-��⛧�Wm��P���r˘��(�6�����?�M�+������i ��E�3_h8
� ��(ը���=3jhn�&LeІ�l�\�<>Z�����̈́���"!)YT� �8���_T�X��}�82c�$�Du��H�����`���y|$Xx.����������
�A�m�˱�73�h�� x#��r{Kl����s�Bӈ����S��Y�a_��RLs�.Y��=�ݍQh��+�+��?���LǑ���G�� ��<�@FH�0�4���҉&���Jd({7��3�#�����s�k�^��z��������S��NS�p�MOYE��"�ۉ�n�䛨�\f�9� �Ojr��Q��SHR��[�����L: ����ѝs�BO��p퟿��~�xp��㭦�O����l����HȾ�u������=�!{����3N�'�JHI�}{�����o_a5�<������k�@߬�A��P��}�m�!����:�Fs~(26����/a������7^�[������84D�pw%%������IM3����loo����,i��kj	٘W�O�����W�V����{*�<��8Q��95i����gC_��D�onl��h7<�� ��n�a��-C�wm�zF�`JX�[iz Hz�
̑��4����>�v�zw����l_QS՗~����bv�up_vEaȳ'o�=5\����v���+��g(�ZNSj�aAZ~#��}c6��ϋwd�����{��0��k�]�,���>3K������<DoJuXq�-f��>�s}3W��N�#v�4V�9���"H��W�+��P[lqe/�ϔs���7\�4�
�*����e���,rJJ��¶���Y��P-B#�dl������E�l<����G��f��h��#>INe2K�ݽ%���GV��L�R������0$}}}����,��!�.�ju��'n�:�>�E7�c1�RNK�u�T�Y�Dy�j�U(��M,O�G\h+jLl��37cdl,�����L]��bQ����?g�7��g�
"���/�IZ�&�|CC���׼��2�*��~�^�	w��\��ױ6���
Р�J&�01�7�׭��7��K��x�qc7��6�l!󻄥T�cx�_vn'�ތ�����q4�ܿ��6Uf1tũ+J�Nɷ�WR����|Y%�([:3}鸧c~��~z.k�Z�������!�8f���R� ��3*�;-*�t�7���Ѽz]D�Ϭ��Y)}���3���������*�ϻ��~��̯;yk�
j��6n���w���L�"&�u�~��C��C���f��j��������m��Ĕ����j���r�G��?�k��c��"�VgQ�os���x�c����f��49���b��yBn4h����;rkC���,U��چ]����,���� �"!4�S�'~�\��#3up�pJ���̶"�ӋU����U^��������;k��E�w���"e����H._N�'y̸�{��&��NP_T6:�#8Vt��ӵ�WZ��f�Av�h.X��/,������[��f�&������H��"K�DbU��f�U�1!���#���4�e���lN�uw��111�F\��iGA����kv>����5ӎ��`NA*?���Y�P�n�Y@@ �ݡ�b�{��t��Bӏ��w�P��4L���h�،��	�Zn�����AX>JSV�$
���0�`��2�ֻ�X
������+�0�~f��n�ZZ4��
�%�[*���e"S\��68$.�Gr�x4i���07�	b���F
����G�!�ImB���&�����:��;j��������`'GхD�E���)�Y1��VȂ<��8�֎��@�	(h<�=�"
i��х�$b������DPS]ͦ��I!���.ޤV����qA����a�C�o2�*O�1窴�#MޓF��������A���I���|||����pLIfZ���ts���k-�-�����o�u��H�2�Ȱ]:�=z����M��̪�bqD��T���������k+=\IqqVY�����h�X����Wl�ծ�����T��eȭp��o�}���W��ӕ�jW��PM��z��3�j����H���WF�TW'$��B��\D�H,������%G:1{�7��}��|��-�#7�J�A��Z|k�I(�M֙-���oߒ�����GV�������k�ec�����\�q��/i���S�G^�$s8��h��D�+ !��Y��׶�P���C?�<�tu����Ŵ��&�UO4�!����O���8P�1����6_�W�?���v;g�p�R�6��ξ�����ނ|w�`�Ci!v�9�c�j���3!�_8,��<?=\��dU�t�M���>U���������"��0,���Lvo�o��'gZ������3z������eeeU��k,���R|�C��9�8P�)��#&�*�ZiF:��\dfYD�q�������[o~v��_EE�A�C>U1(&�0��a&gd'ZnM�k�<����%>�v������m8��A�H��&9Ar6(r��h�`���:ƒ^�v2۲� Ò[V��w-?����52��� 1��r�I�_-+ND����\�H�RR��׸���(���7�D����ې�M�2�I�^�Upd
;	�!�<�����ش�x��%�V�UVl���`vfF �<~�4���D1�X	!v���f+��*�z5U��R��zS���#~Գ���������Ծh�_��7�������<i)��x��6�J,���!S���p%_��s�S2�=�Cm����6�Ml��s��;�"{):�黄�Ұ;����o#�A�V��$l:C_�_=�WĠ�!�dvk��EJ;�̊to�\^٬3�
s�������C3U_\˪��g�ײ����x�%�AYe$��Y�Ә�D��Ξ!w尽PR��ds@��Y�ͳ�ǝ��e)2���슬��M�_)l���@;d �,Kߞ�V�QVum�	���X��l�v~�lkk+�)���Ũ?rc"[X����IO�e����ѣ����߄M2�%�k�?�pq���w~��"`�Kva�T򆞞K�uljJ���g������@�үIs���̜�H�\��S�_ˣaS�9�~e&���ִ�DO���?�A �hs���� ��6�zp��Ժ3`�"���#L���1OY�;��+�
Q�yҔ!��S�OJIF�, }�<*=��&��c��_"~�B�)��EU�'��kނ:����Lxڍߺ����(8C�mI��w��D�.�V���\�5Z+�ͭC>.S|���i0[nCL2G�)dƈ+-�%�7����N�z��;��۹��<0!{ee�f������Y���|�R;���w~r>Z���;F��	H���=�Y��3��#�Q������fxA^^��DذR���z5�p�EB+���0n)J��K-jW�@�?ITr��6��&=�l��`���d��
�K�����<X�>��^�<H楱b��E	�)g�L���Hl0�/�k�,��;�y���
 �ե-�'',HϑN��}FS�A\*�wAW�P�8w�e����������2It�%c{0���x�p�^��~qUW�#g��Vg�jr�i�0��m�['P���K�H��I{#/'�7�օ�q}H�/��Fi<�Zɜz��)|���}����+�_G|8�O�Р��|��:t�OH��UoS_&i���!����mZ���a,hN�V:m�?;���q\�r�:��&�C���K-�ؖ!E2�Fl�N :�3���qQ"�$}�BeR��$L��H&>1#G�H�%@>ȃk4SG7�|�llZ ��ߥ�Y6vi��7I��f|hW��'X,_�o/�]^^^Y�۶�}{�	@$FY�n�!�U	I���	W�[E��CC�R����:N�B\�z�xg���жur�����CQ��lM�����(�����HF+}��L��*�m6�P<.��r��}�����}�#�ͽ�5���_Y��H��Z�&�C��Y|�d��v����`�,�)D�p4zW��0�|J}r�����6��*�>�Ƭ��'�H�|��l��z���*�͡�޹ wa�FX������iLR��	ZN痈�Qyz���A\�~�ncA^
�/�L}��ڍ��B�����\#�5*�U�Z3U@b&���FI?F,���7kb�Z'�%�+a���7���y���U_;���J�s�.�(�	���q"� �`����o�N4���H����|B���D;�e�eX�㣋���7�<>�F��q���Q���zE�1Z��W�����ZkN��H�� 7I�c��B������u�+�^���GّT��x����H^yҩC�줈t��ʯ�m�>���f�A�����t��X%d&��c/�Y�g������[7��~�6$^��Pd��+ڎ����߾i@%i��:+̲E�|���x�O������c��==��pN44�ٞ�����Ûc��[Ň{C`q��;��F3D��8fT���'I�9����Sjj�6���������,�UIٛ��VI�FL%ᇸ���S��tg%���+��jƛ��Y}�4C��}�w�yr��)����)�A���N&N�qRn2'h�"�����7k���W�1�I��Mv���[O��������c'�b���]�W����R����৿�CAI�#�]��)g���`���Eh�;O���������/�7�1^*�r<(^P��0b����*1T?tC##r���`��C�B���bZI�	��������1�wc<�O�quuW:�)���'-�4��0������UJT���t<U�HJJF��{��U,�ᧄ�����#"�n����|>W�fq�5��y���T��t�X��Ą����g�^��%�+`��O\��䏖�������_�8-�Pg�mi�ɡ(t������`�J�{���G��
]y���M:���Z��1���9B�I��:�y��`��mW�dI�I�k�	��#�ɔ���^6[��i���L�B��'��~�+�ٻhK�I�=<"dm�:�Yg������-J��>ՑV�!����������%��M�]�	j�R�%��s��k�̝��>k��E����=��(9���q!T$5�T~_��/��'VW��[�T��4�>�7:�Nw�yM��fCi�N����&�tW�<�T�K�o���a�i���`L��>�9x�h#G�U� �
+	ꟻ�$���9`[g�����3>�����R�=�-z����e��wCNPD����,�CQ���d�|Mu���/����F�*ϱ�3�1:��ڛ���ׁKߣ�˧E�dW��O����<?�*������� �I쒐��hhH23�W89%E���/gn~ո�xOQc^Kk���K�TgKݛgg�Ϧ:��-x��»x��H1ߊ��b�ߟ�ۗ|�Iv�	�tc��s�	�O'�p����?�Q�
��	���So6��4����l:���b"i��oT��/���(�q?�jU��2M��Š?we���N�Lm�TA�0L��p�]���a�xKb\J"2����������2+�p�;�Z��|��h��s~��������zyM�����>�����!뙂^���q햋�d1�퓶f���}p��!|����kٙ���'
0���ˉ��G>	F�"�B��ZMn�r�^�UD`��,T��Z[uhI��HZ��0Ě0j�䧏�Qrw��]M*��p� ��4����w�Z,+�0�d{T2@��y^s����*�`=�y�l��S�v�S�q�0S:��w{{�2Շ'W=_�|u�G_�~����4�@�47)��0���`��wv�S�ś6�P~���>Ճ���21����qr�7�y���V:������(ͤ
;�;h�A�%��E�?vܟޟ��-����B}C�q7��#��ظ���kVJ�<�q�����M�}|��"EZ��_X9�h�Ob��O�Ჭc��E����*�W'���mǭ��oEDZ���Rػ�q��M��tE�h�*�XG��z|��[V�{�^vV��ş|S5�`
;Q��c|N�R�����t��/4ш����i���i��NAF=�oP�?���������ֽ�������:>1�<h଑Δ4z��#�M�!�K�� CH�$I	}f�>&�]ޏ�0?�p�����M3�KK�7�{?Z�D�1�to�6��I����NQf�����Ȋg��3�ߔި�D5`ߛ648r�D ��O��&UP�WG^N.��¾��p��mTF/F��rK��+����e�{AЏ�	���_C�x�>?�_]҆B��l�Df����y"$6+N���ٸ����$�y��G {�Wޫ�Z��h �6FR��m�:�Q%��|�3�W��gh+2����U4��͋2�;�tr[[?��~�͓O�B�ƺ1��c���:���l�)��w *W%�x�~�Ǝ�ȵQ��\)��H�!c��5[��fK.����%HѮ���l���_bT%�O���v��B��p�05�����L�C�
�iv"�,[(k���Ψ�|jjj��Z�;�E"�K�.>�:I�O\\B������o��k��ض��m;OlO4�m�6'�͙��Ķ�v��z��#�}�O�^�j���4%i<������uc۰`B8}�o~�ZbdzI��������i����ic�G�G�S�$�z�=ә���;;aD1�[�"���Nգ��4G�D(��73!��=|��D�HT
�Dů˝�������_��CZ�b�%,*F��dP�)��T5,��F|]�4R��Cvm��3�\,\&�f���+Y��D����[g�0o����ݴ�(Mĝ9��T���
����g'�.�@�F��K����ӴF@ �.PNN�w�G��]�%�Z��ηб~�o`��t�����qh��)���@ֻ�i��")�,3g�ݼ[ţ#����,�?.(o�9���E�d����E��V-L��*=��]^
7?�a�ƣ��Y �9��?���������։��髪b�=>*��Q������`{���Z��2������l���l���JS��|�ۑ� O==�01R;.|'�<�7��n��y���s3s�wj�ğ�����.��Ѐ\�g�J���c��ᑈk9iyHd�%�e��΄^�|�#�(�W�j�߳f�'.�BJ.V�?�M�;�V���d�a�+���8�ߐ8��f����`�	��|�LQV!��6��e�",��E���?�Μ���DLo#�X����6 ~[��D֚�L��>���:;ccҡ��B������⽨!����z�D@�~s�ʏ�S�|�U���yC��D�\8Q�J��	�jv�k��D
���g��`K�����F����5��ODȣ���܆���������F�Ay�nL:�+O���m���v��]>�k�� h4���
}�����{�=��}+�\ \����:Y�nN�����ZN�ǽ �H
�X}��?ge�8���Xp�3��[���`� �j�/�H$(���i>0�˄���$��ڗ=��feee~C���g}1@�&b:�5?�t(���ÞF���|	l���O�i�gx6f?�H�9yYAb|8ܝRk\MI���&2 �k �5&�TF3�9N�v��G�c��k��9�_���
� ^�c�����(=rߣc(p&���+Z��i����QpF�8��Wc"߽�x=� ��O���dv�^4 `���t��	u�,Sp��D�gܸd�C��ل�~����ea����y��4q�]��2��P�^V&���#��l��uer��t\#��@���G��T-�
��ʹ|�˳eqy�zR\�)��B �G6�zXfL�VcZ4b��@�,F
���7�dE:���0�'�^O�������x}�(X�Nx����\��
��?���A�"K���Ә���b)pƭ!�B���R�^
Q)�I�������%��g&C�>��'"��P�s�|�4���Q�a^Z.& `�UCIt��H��|럐�MX�?� ~͛�����|���W�ՍIeK�Ζ�.�,h�� �n�o뷷����~cC��@V�{zr���(����g?0K_l�MH(\_c	�!`�7�}���A#����%%%�T8p�Eq:::x�>]R�Z��;D66'�-Ϣt%�]P>��\�Ϋ���k߈E������x�v&�J��u��]��k�ӳ����i��-��5�����K+�?�ưm�͕S����ݍ�
xtB��`��AX�����v�0#��S��L����Vd셻�E�^�~PPuf
�DZiM��d�8�f6��x��N��q���}�_p9�����H��=�d�P=L��7���:�g$g��6$�}�����Ȇ��h$�9k��xy�ՕETm뽑��$>E����$�=HK��/Ò�B�,U�^x�	+��dU����sb��g����̘:��Eʂ;\�Ǣ�a1�����v:L<�T�<�#h�����㳗��w���7�w��-׿(���wDK�DdǬ��R�J���jj�*���g�%� 3^��3%��Ƃ��ݸ�]��Y5�Y�GB�?�����8���P@�~�(������p@�4�\�g4u�?�*6��}�O�:�j���_��6DMe����B�ڳq1�n�z�!>b
�h\�j�C[��=ޤ�f����Ï�[���-��v�?S�9�B�VX�򽄜͝�ŜK]�"�uޤ��œ�D9�{Ͽ��u���U�Y�p���j�T5mM�W{�x���F_��ʫ�~|\����nKw~F�����������Lخ;���0[�a\�����|?�R*���L�* ����J%�bh��.��'�!���_��)}�	�Gr{�,2�c��oD��A�bNP�DPss@����+(LM�9}ү)&�,���ynИk�5�Y��T�>����z�����/�VA�����6���Non
�Qӏ��ˋ��P��$�'@���C�sN���l�����Mv�G Z7'��hש����ߦ���/����E{����U������GiK�Nu.Mc�B�0���h9���;t�����R��"����K�!J���6�Z�%��F�T-g�e	_'Q�ڢm�_ӆ���J8��q��n����\Y�;�[^��F�.�'OiW��cæUgŮ��A���j?��r�b`�x�ML�c�)yP����̌b��t4�Ա������m2y��Է�Ŏg�}�I���,���OB6��PٽH$/Lk�R���ُ�������6Z�M�$���)L�%���~x�!��KaȁQ�����|�,a�f��*�����Q�4��ݤ*nio��~A��@&�u�.��G)�������z����ūg֟H���:�/|��G�9}�焣�0��o�үwM3�����dd`A���Q�i�����-57.��_�Mz]w��&��O�H0�e�˝�8������������m���PZ����m`=u>?��B�����u:A����@6F������v0��������C�xě�%�Y��>���$Е�v:�6Z�\�z�Ө����;��X��;���j���T6{��=r���t*�z�$�[�H]TK-��;d䘪[���0����CPq����H��[M3�0�{m���:"NB8��,�١�|�jg%:�:vX(�\�x��Sxe.(4ӿ�:T��2�,�]Q�t�dId���D��5�2���k�T�?B��|k���@Z��F9���1y��,��GAO�yJT]��$��%�o�}�0E��3L�P��joP��K������"}�m����Y�"x����CݯV���n˖�~{j�I�K��Y�f�\�&
9_�V�)�J>,)d���e�Q�ykg�x$���z�)�һD*��DH��H@�Mӥ���! p�"����8�5��~w6V$u皀ː�W`8o���s<��̖���/Q���O������f'�t0���j����o�w�c�N������?�;���^~���g/j/w�g ��5�baAiU-^N�!O��>���v��&>O#�k��ߨ��#ý��`�fW���-�,BCC�㻹s��������U�,�X�8�.���!ʌ��5.���$����C@q��Ο��F���&���߿�/^<��|�]t1����+y�W�N+c���P�&��,l�{j��r���YY�y�v�����A;:1&��m�O�w3�t	)�w�N�����q� QE�z%ASX)ϳ�+��K_��]�Q�	�w!��$�W}"�T���������җ�4/�����.�^��YCײ)����>d.M���GQ��J4����X�����vw�X�jI�;@RJ
�@���K���B��Į6v��J������!"��n�Z+����:~D�%�����$�\}蘗U����¢�:��F>���&geE{����ޤ���&_)�&�D�#�;_�E���~H|���o۶hX�����w �Q#�3�u���ᐇ�(�����;W;�u�l��	����_pS��|�ϻ6�����<�\�D���� ��޸��x������ʦ9���di���M�W�e���˷���5P���,)�x��{-��H���k@�����\סo�A����K�X����]|2
�L1�k�0Ij��+W��O���F(����m�����y�Z���������� ��^��d�M�dΌT|Mi��0X^׀��.c��V��%�˧�����..���{�j��
t!�r�����96�E�4�fB~Qf��8��m��I��\�K�?|�mZs��M����oe������zC���_���m}5YE��Qb^2��n��ݪ���`O�v��
�L�^�é���Q+�BR�++���}����
�C�Z��썡���wl���"�?./,GokyL&��:����6�͖#�襷~������V�S��s�aK�Y����H��t�^��Je˷�@��Vx�u�[��k|p:tqA�6\Y*�`��0c7�S��|�"N�O��F�z�����͔��x\��[2�W�M�=�q�����})>Ht�OP� !R��������o��C��'	�N��g.�������PNE�{�m>þ�AU��)!6[geVXM!;;�Ϛ�������[2�]�1�Oɘ��x���F���\vԞ��C6���ڜ�:;��v�Z���ƛ�����knλ�}v3��Ü�1��w�ty&�/u���42�ޡSA�3��)`껹�����4D�H � \Iu�I�-T6(�FvD,D��[G{+Yt���A+M�� ���X�2_�f�R�צ)_�n��˒�����hm9r�M�������$���+,�0�1b��`����=��H�w,�x��<s�Y4FF\Qb��/ׯ?�1�W᤹��IU0��j�
�>8�`���}��X�<��Z����-��/�h�1�;����X�q!���� �@�����<�1m$/���!Z{���}�?},�XN�<��9��d<�E�,�aĥ��}�L�l
��� �������}���U���aB
Prg ��ٴ���Z�v8R���El_���55�[%�[OD��M�(��
��ǒQ�n&�z��^o|䡭JS��J.?kz��c��{asN_��9b�0�=�[�jS��i��ʊ3zZZ�T��h�z//�k�<{�g�V����׸U��
����_����� E����I\ {��)��q㷚�}�_i��880mY!J́"��nYm��
?~>J��~��弓��#�\=�.���>""��{a�p��}���*��0]�d*�ݚ�;d��@
��x-���r�hB�Yt�,ӗe:t_8_���ץ�[how��G{m:�2ˤޥ{;�U���*V�J��OJ�|t.{C�~�Z9qy�
�*Ǔ��D�9�<����x_���X?D\����2��g'������9������lnM���]��0�Ғ�Y�VWW;�����N'Q�5�&��ÇDCd~�����F7Λ�	W�ȯ�E���/��E �`�ՙXyn���j� ���b���J�ǥ����� 5���z��Y��FB$�?�ƨ�afV箱SF��s�bT,��<�yC[
��Ĭ�z]J�J[F�0'�c�,h�v���ֱ1U�M%djZ\�_�Z��P��C��Q'z������-��v7{�1�M��g�fm�h���b��+h`��9e���,�32��Hٱ���V�v���J�t�>g�m"���b��S������I�R�ߟ+�ώ��>���_�$��ǯ 7(����:-d0�����}�#�[S�i�S� �|l*)o��\�1P��6N����le~r��mgHa/��e����}�
��2�8]��]2'3��c������cw�
Z����M�Cҍ�E9s���C���/�C^�6� ������ݘa�s�����=H�^{��2�B(�O������'
�D�gm!ø�;,Èa?!�F��|�xCͳBS��X��+Q�] /Ğw�,��y��ܗ�����,ʯ"���(�uv��?R�xxyߛ���m�d�4
l�t��$�:KWj�M%q3==��ΑIѡ�����vt� �Rt_�����@�2H>ڥnk��
} 蘀�۠�W��n38#�K�}�tbL�q�&���U��6U�����LH��>PC\�Z�/����X����l��R��U�[���������~Fϴ�T�b7�i�	;b};���'aJ��}ߣ�O���\
�dp�=a6����~A�S����������^��A[�R�?��̽�,�:����Uh���`���M�;�`^����j^n?3E͕�%L����ddov0��P6T Z�T"kfL\�	^�6��e��m�/�Gf����8v03�6`��K`�OW����I���Q��ZZ��+:�֤���D��'��G@���m�;�g���w����},�����o5S���y:B5V����Ǧ���ϔ/�q$e;���3n:a��}�M�s����\�. �&���Ta���%�7[2���RO]HH�w	|<�P�7�z[p��2ݮZ���(��ՍD?�H������&�2�����ﾵ{�(P��4VH�V{�;H�>(���3Aa����Uk^x�����<5C��Q+��H!�h��|Wغ��)�2ަ�(����1�AEBR�г�79�p�?�M��V.Bٸ�/ǽo�s�#{"�u�.n
Ff�ݚ��L�~���b}�I<Ƽ�}��jY�g�'/���kT�����a]� ��@r�)n�b���-@j��^���*b�X�'H�/�*����oc��	f�I�˃UVL}$B$�2�+���=cU��5���H6y8ֹ����x6=�/~˪y�P���]��a�{�� �>�+A��(������R�y/�����y   *Gd�l:�I�S
����'�����2�����e��F�|��W΄E��_K�i	�r�`Ҿ$����g����
�c����*`C�"�X���០&��(�9-Ĺ$��PLTF ��Y��Q�2�4!Ro�:��0��g ��(��l,�Z⟓�xG�2�:�3���!��8C����b�@�8�R��Ax�O��h1M���74$
����T�4_H�c�%��Qֈ	���iv��{����|Y%�(Mx�X-)���Tg#���6nQ������mȲ��eگ��	��r��L�H"$��g�����^3W )���˫sJ�vs�`z7e|����u�t�Y�d!�&b��R;���; �|+\�Yr�����Y}�X���jڋ����f�y��8[�@	-�ˊ�p��o!�"}!l6�96��9QqJ�V1�<� �Mè��@ GA����Qњy���X[�|g��+h΢m�m����4܅|)oY=#�ш�ct�݈��W��ɼ�M�]�'�� ��ʇ�S�K^mۻ��*ȁu[�Ԧ�P��"G�ŗ�Z�z�&��t*Kxp��ee����kт�+���'�-2P�HSV�piTǥ`�l:�D�Oz���Fv.km�n�T�R����d��1J3�M�m�u��ǅ�0S��5oZ�Q�g��3/�eW�J��3-
=J�=�� �J�����*��r�k��y�%fq~��fF�kn�T�P���C@�<(�A��>�Z^�~�!`.�7��ŬZ_e$���v�H�"s�J8*r���;#�fT:��~#��"n-cO��.�o����uԓg8�Շ[j����2��q���0��EgI_��>d隧C^[�"��u���T�9�JE��M&!�Q}�6�p'!�F���߆�6yO4��7�����	�ۗ��#���0�&!�)M4�N�q�]�eC���\:y0�K�s�ơ8��ϭj��=yj�7�t�L~��]�@�Р	7kX�Ʃ���:�gO{�i�Ek�6¶��m�T�0�3Hا��zn�`N`eٷg#'tLT֎e<�e��^T<�bU,�Eb����*�cnw)�o]���k��R�ނЪ%s[���G�i�#��`6�8*tgO6������� %N}�p�L�; .u@�i�>�Wf0|�]��7k�i�$�ן<�'[� �Sʨ����z4�Ҿ_~���vV�t�"O�~���Ҹۍ LBm�܎O������h�LTJY����,Fo<��1��x�U: �	H�1��hª�O�'��>0 �I�<���ezZ�Mm�z_���3��>�q�)li��$�xh��c'� 5;W��t�X��Z�6~����׻��[=�o�c�?;7yВ�~y]J�����PII�%�c��vp��X0ئL�O��Y´��R�ڋXA���tNZ-�L~��eW�$4���w�eMΓ8���<'@ή�������D�-�[?I�j6I����pB�.����ܩ��(�Z�e����3ھ��Z��z	L�B"��#"�{���@�C�6� C�=T�����u+�֚x�{�͠��`&E�|ݦ���%�v�r�g�L�XH��y���gcO��s�]q�W�p�e��P��W�9}^�`��0��=���Ң���R{�+��
� �C;�5��Sǻy��I����\�}!ѠG}b�Q`�`�i�:��m\�s��%�0� �?5~^hVѥ3�=�n�*�CP���8ig=�sb�Fj��;_�q:� �a���D\�m0n�!��W߯����޴{���J��_H�c��8���Yu�ğ�q>���S�X�C�/<�%�a,�*�]����!�7��p�1dRT�?5��L�n�L)q�h� 6 ���J�Y���<SX�X`� ��_!Dz�{	*��D���Q����!�����u�}�y�y(�����L�	�"��!���g�����4���~���)G�!��c�{g�Kl_�~��أb�� ��:��@�u0���Gz��\F�ׯF��-�b����b) ��\.�.̈0C��al��c-fd0��M��9�H��M`�k���!���� 5� �0�U�_'�SÕx �����B]PPP���$N*�M�#C15�=��|r�H�`�;��؋íE������b�r�Go�f��"����ðk��HA�΃�	#�4��H���`Q�2��Z}�JAӿ���pZ����-V�ْ��=h�c�c�yG�Fc7IZ�Q،T��BS���o��t����3��.B�AߊS#���ǹ��ɲ0h? c�_�
��(����Ho5�5�svD���7�4k��(4*I�Ɂ㔒D��e���2���n�r��悷"�l�d>i7�O]�x���Q>��ͦM�-�j!��힔X�tё���/�����c�W!���C+.�d:��3�JV�P��Qo��Ȟ0d�y�+Ds�O
�X} �PQ��:�{�څ��,ZA�7�u�X�D�����\�%	�7:�����ܙJd���t]��@��_��x�0ek/]ȴ��I��Wd� �,c��Ch��m���Hq�P�J���⫐?��/:��1�&,@3��ok���Ж���޿ ��m"7�!�>/=`tL�U���L}�uG����W�\��؄����K�h��� K�泇�h������$��hRjWݴ��0ӱ�h��Y�2��)��fq���ʽ��o��>I �ARcR�X���%�M�2��8����@��=mFt(ߎ�,�3�/LdĬٷ��q���M��
�Y�H�([/�����v��Pp�F�|+�z`��#��OI�n����&�{�c�i��nD�����q81��Z��2���+!�i�!�����Au!����n���I�eZ��WL�&Y0'8şW�h%��7=�p-t��ZD2���j0e`\Xl;<��,ѴN��������� 7G�
%q�qb��;��WTx����Z��U�k�:�������0�����ف��;Q!��G�Ч�p��;v\h� ��D��d���Z�r��"A}<"}���ZU�� �#�������ق�+c�h�@'X8���u�V�ƅ汫-Z�Ԧy���&�߆8�;2h|z�l)B�U�Olݞқ��R4�h�[��X朠���� t:.��r�*u��I[%��� �֫^�¢=�i�E�s!4�F@��)v��.�і����2��q�z� ���%4M�u >�{���#S���\���ޞ�J&f[�2Q,���jW��?�� 4�8%	�|��R�'�r���*��)9̦C-� ^�ɜ�������1�x���MJ�S��T��<=�|����78 O��k�R���`�)y�'b���hp�#p�NAE�=;�"�J���d�s����!b�O�
*�}�� � ��Lut�"�4f��n٠�Т&�`\�y�S�r����.0�:�$��]Gp�z֌��� Wa�wn�F�F����/��Ųj#�qfx&�q���L		}�w������1������2D+�o�w�:�VR�htE�[���S�iچ�LZ��� Ö�.�:�*�]�08���j@���������[f��Z��Ɲ(N
��&��!.���?r������ƚ�gg7C�8I8������m��1�����N4o�pd=�NwF���4&����!iV��1M�J�Vi���8/N��$�BzfvHOzx����������o�r���
l�J=؅3Ј�����T�Ὶ5���ou�{o�����p�4_�")�����������Y�0��T�,���e��H(�5-)���l�ќLf$O;��5�`�/��!G�n-� (�x��PAU!���)� 4�V�e~���('�̔3R�է����S��w�#��d�M��DH�熎�8"��0�K��G-Z�i�!Qàa�ա�|�RÓ%��u���.*&���o s��V��_���aӂ7��d@bT�x^6>���7J4R�|7���𥸻C�C7��-�o�p ���H;$E�l������CCC� �%�3�-@��ݐ�R����Kq�����yk^Xb�q"u�
U�U�\�c�r�K��l�Vz�(�Ms�E`�]D..�n��
�eBb���Ȁ>!�0*��GK��Ix�L����������hTnč��vhBBv���+(
V���R�{k=%��x��Y���&$k�O0P��B;]�����̲q�x��%�T�f��V� Dw������qT-�Q@tF� l��..lzi���ln�$xB�8�;Y�DȆËG����G�����]�'9w�<�}6�����䬬*�r�iZ����e4�I��!ūH��ź���Ӎ�Ԕ��P|G���ґ�z�!�$>�Ś���t�H��y3G!Ze>ʴ[
n���(4�Ӑ��9�B�gg$T�Vq(�P1�����G�(����#W%z3�_�TU7 ����I
��?�ZQ�4HR�2���V��YH��Ƿ��Īo�5�z�Şp��0���0����I'��0����������j6�oli�1���ÖYe�_�@�"���<ڇ+"b�*�r[̫<�}�pV��Et@-� �e���md�>]��)��̦������:Mٱ�X�'̈́ ��``RV�A��1�����~I�G`,���]��x:��l΁s�h�i	����1F��@,�I��bϜ �tQ�����K�~2V�R���	sDd��n5T���U����,�?
5���!�������2"h�ȟi1�f�looo�Sx�"��>F��v��=������ܰ<�ꐕ�=�Ј�ծ��"g�����7��6g�mؔ��_��qq�5��}K��q�iˤ�H��z����m_@V�x
ͅXd���hM��&�,I���քU*ů$���(����8��9Rѳ�E�k�z��U`a�t�t ^cV4�_��^��>�\��ow��9�>^�wY��Jx ��騛1��{UG�R�����nA��=�����W�'N�&pW�RΛ�qmױ��䑅��^��_q���P�B�������~� =R�{���1�u���XN~����zy1�6���x?{ݥ�`L���Ks-��Cₒ�~��x7���7cL{n$�ܖ�l�A�v�_�fy��BN�8��|1N_�|t�ba�慤B�c�������SZ��c�+���ΩfJz���@H�'�5%�`<+n$!:�S��^g�D�v�k4�ͩs�X9g�Edx�p����US��?Wm����\{�S`� �}��i�PK��c�6(h�f߹Εr��K"lq�l� ��gT���!��b�~�hC�?�*��5l7,~�>� ޚ��<��?p_É��]�[��?K~+�����&�ͳ���L̂;�^#e7�V�h�c�M���_eV�6��D�iS>������s����p�gZᔧ˻�P�H��=�)�D��$�m�����&��J_�?�;)��u�
f8��Q����89��IJ*�tVx��E+$�4gTJ����ɐ�v=���f3|֛�!�l�q�e��CaAcē�;[���o-�q�d��u�Bq���5�4z������培Z0`�+W�w��D�C\3� �)�`m�~�(����������g���D���b��|����Њ� �:(�[���P��9��r;*/�l����hz�Vs��õ���߰��'~p���-�a�ؘ��ڥ���1T=	�~�f�4Y��d�AI���^�m�I��yΗ,�Z2�J�C�0�}h7�=�y����t��Р p-g5k(r�/��=e�R{ofڙ7����/��z|R�Ks�5Q�XYaw�͝
����]W��K��h%?+Ҝ�԰�^�#�_)���RR�0�'5�9�딕� Ϸ,��]��5J�|�C��$�+J�;;�0)H_S�9BB;��e���#��yL�/��:a)�BPV�{%���Q:�k��x*6C,
A�/����o��aC������j��B�"`�U���Ĝ�5iJ�ާ��&x�ۼ��j�~*4Y�d��!��������z����DK��Exgp]�������g�7����hV�n��+�WPR2|9%�Ɂ`R�G[��o�Pa�/��$���(�)��)�f�(�;��a5$j ���&�V���R�$$d^K����k��=)�2J~<��[fُ?	"���ܹ����Ғ� ���5=UU����
�#�%wn���xN�l>po�
F#�P�n^�6�C��ez�T�����m��u'����(�Y�"9���z���6~�#�m�j��`'����f���B(���g�۟%*�)@�Rw��S�<I���a	۷`��u�����훂�ڜX{f�p0�9���;ݩ�L�U�[rt�xғv&���Ǵ~'�zZ�u��M�9�xjJ���%��}|
*A����:N�ȏ��j�W�qY��1S���d�!b���q�\��(�!�Bc4��yI�[��7�"5��RƮ�T=n��Y�~�&**Л�#�!!ӝGU���	���"ԙ�0�}h)k����v9��l0�����D��a���z">B!a�a8F��<ҍ�Ȇ�-/��*n��d���j06�����E�V�6��$�0���g[���d ���YW�{�_�a�/)�q �̉��BԢԡL���)+��2Ę�S0����p`&_�w��Ծ��~��f���A���j�+��n�,O�,�?J��禂-�ݜz��	�b�Z�B���S�3�}���~�EX���ba��Pć����+I!47?v�2�U-xM�OO�������������}W%���9zX(�E]Q�2(K�0�����Ժ��HI��'�9,+w����L:кC����.��i�rsƅ��m�"�n߮m��혜 !q�\^����	~$^��Gdl��mG��3�Eh�@��c���d"G @5���IKt]m��i}� ���"J�N�� ����A����a����
Aߓ�ܼU`��1��4AG��2�Zh��.�7x��k��h�����cE���8��V3�3��})��kX�c���K�9��hX���%g�0C�Ň��~ ��|%���9mN�q$­�'��p��*�w�#
���]T⮗L�T$"��f�c��w`U`XSmdzU_6������"�NPt �R�����Y"��4���h;*�,�?y�W%�����^�^J�8�Q''_�w5�m-�$��R~2�,YDH��9��t����ٽ��Ҡmc��@��S��a������^�K�FF�Cߝ���H���h��fbl�d0�{3ݾɅSƎDz��
k��Ԙ̥��1��V�/j7�������@����ѲJa���RԎ�'�:�x��Ԕ <��X���akp��'�`���#� �=���CHHү
$�64B�1Wz��z�«H��{�_,pM�Ϻ��P	�-��g�5@� �7���Ip)X/�K�:����i�P���]<�7��S��|�?Y��u��ӫ�����o/�9�D�t��^�Y�^�PB'2�_.�����;�	��?.g7��'���b�n|vYBI� !�k���smL�찁�Z˅�t�:�.`'���֭����&P��@Gw�8ŏ�Mr���pAS@?F��nf����J��,E�:�级�	�o  X��B�
� Nd[�wC�r���j��TQ��<�;<wn���#}������? ��{{��K���H��>�N�֣=������ﯜ�_���WR�O
�X�%a�������4�4̗A��%+,�C���Gv\��Ae>��,�`-�#>xE+��p�������Y.����=��`���۵��ݑ�ă��<t\6g�@f��ki=7�=�|�&JF�틈 @j�<�x�g8��ճ����Cq�Or���Q�o��v�(��ʝ;cώ7S��q2s��;O�2w9�E��'�&�e�6�!ҷ>Jmm.�k)]	����-�3�����N��;;�C/���yٔ��]�
�7+��q���A��PVV&��\����N}(�P�3�>�� %G����>w95�ō&"BYC�4�*Y@>�)B��{�zp��[�0!���h|�x��F��A�����&_���Z�� � Y��ͤ��A�W�n��f4�`�����}4S�(Pc{�'F
��)*�x�p��R��b�pʡcw����{�O��`m���z�R#��@������r��)��́�V� *Z���ca�#�7�xI���l�Ϥ��b����Ҹ�;��{q��h��!4��"|���^���v5�9���	P(|�$�������1ش�	��sӸ��)�@ab��x����ݟY�,�Km���F������ﾝ��ա6K~Ш��{ 5���Z*	�O�2U�����
��	1���!z��O�����c)C�R�1seh���� R��O�!'4�Q�����xx�rXRgQ2$����mo����<ˇ���d�Ox<�c��ʖ�q�18"v�6!��]?�%gs�r�ԋ��nl�>.�I��;Y�ʡֻ�=���*
���C��T�6�٤���w�|Ehwww����W����Ef�4L���<ID.@�Oţ�g��o��5{w�z*��<�[�a����7�]����R���f
��ۧ��@��Q�6�ƨ�_e��~�]�(K@v�Y�믪����ҫ��D3
*�ީcH�E~{O�V�z<bAVa���E/���/�=d����Js�1y�z�ٟY�Iz�"uE8.�֫��ŋ.�@-4�OKO�V.OK�|
�>K���
��.��w�r�yT��#ަ4� �͈'ԦN��qMpyv��CJwP���#��� ���Aǝ����a�������҇�h�krrrcГ@��gxYY-�IѐYb>(`��)a)҄�U�&4�kg�����?��k���6����ϸ���5�����L3����|����b�����|�æ�H���P��wHQ��sK�2��D�u������8�Ɲo2��;T���Y|�Ai��U�ʛ>3�+^-��3U츲��s��ٝL�l�Z����-�������p�S�Kmُ�w2A�7Xz���0���,�&2-5s�'��D�E2�j�D�ȡ˼ʀ� iW���� ����h��ہ���q��m�2��_j�f�a@kU���Og�v ]��������'�&���l��P��E[[q�L�e�/���#��/�8��p
  ��@ժ ��m�y@�G��I��n�@�#�����Pe�@�Y�q��D�K���/!a��̕5%��؂������eט5{>�x\!�2��l@4��B,Ș3<#��w�`؀m��������n��i����ś�����d�i���2p��e#�����.6?~�)5E;}��Ⱥtx��ol~h�_�-b�,��o�wF	��O7�������,L������4|a8�-r��U��K��M�""Z�L�eX��6:@pw����wM������%@p��܂�;ww��9g��� �g�j�Z��b�`�}�U�M�j�7�EN*Kv�Z����C=���Ä굲����:�q��]��#�-��B�C#C��U%D���f�J�#��g桩	ZW]ޠ�Ұ�d�I�%:�mJ���i)�<��m��D�饤�rV��`�OUn�ڰ�<���TsU.)T�Ъ���
(�dT��
��G��ѭ�LD���m�wL�I�
�2��v8+i�*U���fh����QE�R��R��ʎ�B!��[�eSԓM�(.�r^����,���h�A ��Ÿ�g�z^x�RÍ��:����=��_¦BI-P'uA��`~���"&=C��X~�_uL�0r�λ���}`��j����e�_�unw*Ș_伬InMNmk���:����b��J�L����JYi8�^��"��ov�
����������izX����P��w�{��O��W=<<�+i�j�߼�z���+�W�7�q����?&�{��d��)G�5�W.	4#@���Ŧ�{V���-�i�t\�i�Įu����#x�wr�#c�?�bU�I2	F./����*�~�x�2uW��O�%��`7Ȑ�	��3�F�������%�Z;��|E*��uB��J��P���a��J��j` ,&Wp�����uaN�P�|%��"N�Bz�k?��	7+0 -�b�u���>>_�0H�tY56rk��4�|�*7�xx�z�0^�X�/�m�B��{�M�Up�k�:Թ.���
܆�	��=>aQX4�$�܊�9w�m*�������o�OƦ�ӫ� �ϛ�}��a"x��tN���i��B��U�ׯ8���d��@^��4$*�I(-��FF��.�H�QFE�D����[NH-:6����qؔ(0�5�2���A!f�({�Q�_O.�J?��r�蚙��È��t��ݻ[z���)Q�]_�}��xN�� 䈤�m����vݞݽ� ���"��~�q4*��+�ץ��C*������s�f��2 X��d��V)�Xb�1�!A�hΣ��|���4_�%�muD��	�����'�;`@ݚ�����hۤ�Y��Ӈ`樃r�@N ����Qo#l��=���S����l?�����0��&`iu�d*�U���B7_
W���G�r�d����1��3y	�ۜ����,��<=(1�授6�1Ƨ(�K�z�ۄ��e�{�F��Hؼ�58��Y������z��eZ*0�]�/�Ҍ(X��hd�|p�D/;(m���{ˮ{�5�S1�,��H�#��w�����%a���+D��s a������`��d�ʠ=���2*��׻�O�
�����v����v�Y�`����e���#sDt'2l<j���7�ۣ���֠��\��"��'�O�ho���~KVE��]A�嘫6W�*�CO��W/��-W~�?�:�[�Ԭ��0l���;?w&�B�E]/����8�����@UbTE�������d��	��{����2�F���EO.t?iۻo��ަ��;�]�c`�;"�|mb@�;�q����FE�hw�?�[�-v:q1Z�o��<�����}�0���n�)����˜��l҃ޓ�T��R���9`�O��+���/e���R�u��r!A�/��|O�.�}��B|�ONR
��k�좢u��=8f�p[�S����e0x�wR�t�^�ڪm�|fd$��r;�O�����2�؅X�]�������f�4�� ��?S09z0�V�_�\������^ɒC�T��s&�C����Y���%N=���8)I�vf�W����nS��>��P�oo�̙��;o�-� �s S���n�Y�-�Dp��n��ǁmL}:P�0Z9�1MZ]�Tzׂ<���T���gi���������!����vW��Y
�<<o�<.'8��W�JpD����ظy���U:Ƿ�sǈ�l?�)(���&5fX���K7�򠎳Z��C�������u�o\��`Yr{�QbkJ��Jo��B�w�?O��ak %���q#��:�sٕy�u�J���h��v:���&V�Dp��5��jc�A]�o<���u�Ů��4e��v�휜*�IZK�=i\�0����ru�[����&"�)-#s��P��w[t��r�������>BG���Y/��^]�.��$�G����r�;1�<a�����V�@�o�-�p7��z��+�ֺ9zmK}R���I��n_������^��K��f��a�����w��	�	�����p�PVF�l�?_3��>�Wn>`�l�6e��R��ՇGW�K��"�;��"���f0���0��:��y�|�t|�<ʿ��xM"���qZk�����8�����%5�ke;�w�:x��/���L�q�?�i�rE���+~:�LM�t�(p���a?W���y����3�Ȩ �C�����Mn�#���iZ.ɚǰ�վj�#�!�ilV	4����Q�ͽ�f���w���ޓ�8/'55�o?���`��1v�JN��!��]sKHK3��S�'̇��Ԥ; R%V]]=trRI��Bӏ�,;�ڽ�P��;n�T��~�
2� �N����;c��tZ�������Qӏ�̬<ʑ��v����^�����%^U��HII1��P����y��S>��*�-�9>������C��P�}�Wn�Dt��˭���C�.JC��G�q6Y��W�a���&������vG�d���L��@�X<�4h)��=�����"���{�N~��F2@K]�U-Y0a���c{{[I��n==!'/׿�L�ըF����Q�]x���E7N>��w_��b$��;G��N��x�����} 4h�_��w;��˅������g,IM��d4�b�t�\�Ǐ��R%�qѰ�[��)U�j~����WO��z��W����5��o����/U���:��k�/ݻ�̄��9at+z�&�ppt+5ǧW�^��:����4��+o��m��ٴ��0�+Q��l|.�Q�ɘHن��K����?��sfR�76�	G���e�Sewq�性��F�H������mm\��9L]����0�1:�)lol�T�T{�?YO�
z�V���G�!	EUUM���!~�h��u��j;`@��ѽ�~?glq;���ed�/�#=n��u���q$F�*k�[�z)t� �3��ul��0�6��l�
��(�q�z�z�M�4��=�Y�J2<��.|�H�?�3Q����W�u��x�����vb�\Q��R�ا�Ì	
	�|-�/k��~�0����w��i(�̡��r�;>So��O����-V�h=�x���ׅYB����k���&�H^z~�x;��ޚ�w�j��1�E
��Heq���h���>K�o	��L��0��:*����KL�������;����Ϲ��=K-���([ʣL�v���O�!)����VF��}��sR�q��[=��ӱT3�	�eU�mwz�7P�3ɢgZ�. �r��V\rl�y����.H�`�,��b��`+͍;*�!x�!�GOG��J
Y���b��T�k��훊~p^+���r!�^�VL��9��m���A�J�4eM�#( 0PYY���9[�)=S/��}tִ�7��~��@��Fƀ��.GUD)$j�8���T���M�V�-��{�:T��uڋ�9O�ǂ�S��[�����k�kĚ/OQX�=[Ja̘+A+��Ď��l�Zdnni����::Z����p�z��GK�������l���Yv�_��.cO��{?6�s�Th�曁=E�i�_��]��/ �֠��5�"�����m��qzc*&N�-tʫ�5Qp�2�+p����窊���5,�������SN�oV"X��mb\o=������+|���"�ҽD̮��M�'���8�@��1f?�)d�gU�̎�0@���{�k��`ڡg�
�z��8��5�k����r�ʾ������Z[�yY�e�������W�4�c3C����ݡ���$���LV�.2Yxtt�=��K���}���\��>�D�m���Tֵ~�}�,�赓�]�D�h�v�����۔"gSC���"�Q
�UUHm�~��Gj����`NW_%���|�-Gb����-�� �N5���,	-%�'�Y����^0<}��iy�i#�h�)��e��p��Xc���>�������vx�FB�vU�MDR�?o^�ի��OlI�.����XL��Ξ����4ґ2e�n��ZV����[�5��֝��6|kj���cKKgUU�dz�j#�N%��&�4�	�\LM����a>i4X$�"�V�Kd.���d���ʛ����͵��7�5B�%
��R�@(J� w�h�[��"7�+ď�|;�3���p��}�v:�n=�!�PQ��{t	M���2��L?P�S���+����"}���mL4�2��o��V�4,5O��s{8]t~x�^緦#�S�����@!���Պ7P�+^˔�R�޻B=��e�����}�����*S5BG����ds]��,��~�^�BCd����݋䂍X�㽊�j�'va�t�:�%VEee�w� ��Y�'� Jl>-��ڀ�(HᤞI���@A#� .Y]!!�һus=[�?��S0q}�M\�u%�|�62"[�y�.]�LK뚘�^����ZD��Q4~���rﰒ��ӧ��uv(tZ���Ԛ����ϞSgfX�Y-��y��T�=����f�&��YZT�����?'���o�
>��uQ��3m--mΑG����sT���0f��QD��׏��+�1x;���[�m��1[���6(V��j-��Zd��u��֛#d��Fu䪼Z�N�������iy�O"$�۬�#���?�����gV_XOx� �q,��S88/QQ�������,�o�r�G���=���'[�yx�������4����Y�Eұ���ק��Z��l�Z�'<p�ǃ�DֵM<m���2:B(���ko0�JWy�YmF�����@�o+�2PYy����=H'����������ݩ4`G���q%$fNԱ;))V���Պ$�F�Os_ez�5���Π�&=8><�2�v胑�(8�#�FCJNN�Z���h��">>~�z��xϯi/& ����!����j"x��S���1�˓�琍0F�_zdpHHTI[�߉�:&�H���hr����ܬ��s���h~�Ʌ~|�P�ѿ�uZ��H�JAq���n"�ʬ�91�!il�8�P�Ƽ�ff�[÷R������1[��M�����R��[2j�J�a�'�DF�'$&�;ML�&&�?��m�aw
 ���۔Y�b6D�~�UxT��U3��K�lmsE���28	r$A�5_\Z"���_^��v���
��d8:>N�4t�]D���I\x�����k4��آ�8d�� ��彸��m����A:�`�$��3s��u6s��jqgPS["�3k&sCQd;�Q�q��fچ��,�;��� B��k���x�c�|'6�7iMb�/�hݥ�F��6&��߶��8w���8�FJ��pB#�Tj���e�X��ϸ���LK��Z�i���w-�&[�iI�oph�5)7�V�\8/�p��0�a��J�����e?@ʉ�}��UU��$�A"P��Si0�忓�����P��55EXĬ�Ŧ�����Z�jy�<�
vT�D�1:� �l�����'̆FGG�'$���a����	FyT3����~Lu�T�5_�ns���h�[��0�VIUz#�����/�$��2�'sE�h�TA�Ob:�/j9� �� F����:~W���� �DDd�o�;�}w�x�e����4�)R{+�og���"JC�nN#�p �\a�@<[o��ʗ��[n���1A$.j�J� �l�-�@�Z7�=gc��e�Aj��p���\��Ӧa�T�mw~�hQ6�pl�@B�+\�Xanh��H�h�L'%�ێ�B�`�j�E�O����2�+b��E�?2X�-��2X���h����"��呦j=L��u&��.�#�y��H�6�_�zΘ-�������h~�VAAA�&ߛT(D<�Zq�M�>�I��$o����k\Āz)z��㉽B�E��13���|�K���	�����j��������{�ծ���|�V��C@��_��خ���粱�s�̄<���X���5������62]�֠�a�S�"����+��u�G���|�@(ZZ�#|||K���a��E��t����W�D^ި9�����ж{4T'�"��Y�ƬQ��������<79V���ako+�sO,�Tqj���,�:)57T|�Yn�z,@���P!-�E.�0����7��%1�P�*3 p�l7P/�~'��@N��i��Q�3kByxda$�$���W�k� 8���9|ej�JSޟj�zzĐ����>Y�'�5̀�������y��b񐒦�"�d���ob��d>Eei�{x:�L���UM��k#�O��U�����O�.;++ �ւY�[.�#��l�\B1�t�����^�h^�� ��'GRѐ���L��l��~�m��Wsf�x{넣�	L{k����[l_��v��G������=F�Ԁ� ��of�93��l)+��&�P�l����=	��aq�SL3����J����"gE��gOH����6x��
��7j[}�:8LvT�����0Xqgy�([T���-W�"L���p3`�&aM{M�:��J�/����	��pKW."�P)�rjjK����v  �9ɚ�+�P�J����,dK��\Nh�,����­׽-�%<d��U0?��?�{�i��Bg���\}��V\fu��N��s��EN���UW�����]�(�r�@!{�|�IG�'���UY�܌���&�~-�>@�22����o�9��#){\̚�X�^`'�I�y�b�, �t
��oN��+���٠�J���n$*��L�f+@sY/q�ގ��M5�ɡcn���R��+��w�a��U��45+b��w+�P�˃w���7�ӭ}@G��*�f�,�����u��}��3�\�ꪏt�W��VVv$���/���zH�������/..|;S� 8	 Z�+�U���J���m����7�Du�⦏�p^u�f�#gm�M�Id_Jz,PJ��-c|u�(���Ȣ�孢
u*vPS?9���X>>�YQ:�쵨������4�{�"����p�+ G���=�o{2?>
JD��c���u����7KsMN����Ab_z�����<<����?�1@�ߨ���7�p�N˲���o�C@���� JJJ~U��<���1��`�k`�,�?��X#�v�e��U�����	�����h+��P�~L�x�/T-כG�H�� ,d�ٝ�#���e�r~f�є���K+B�eٰh������Zo�d����� eXk#�2B�����Wbe���WBj{.w7�
�ls�
�_e�W�VQ��]U�259uI|�N�S�l�����.�b�C����PCM���W�i�I������A�vݤ6Zx��RLҬWA�.�@����wޒ\��`�^��F�x��_(��5����G���GJ̪��zx>�e��K;����n#9{&I�);'E������"#��2����{�����ޣQ0@j�߹w�ϫ�t�\�Z�4��N5��n�F}����5}J\��߿���O�I��닳"<G�)��]>Q�� ��#��N�I�dt�n�{{lJ��RQ�}Y2ŵ;Q���������U&�g^��EL��r]�ZMI���`�c&���=�ed|=����!�3�U1wtTj�n^��S�}��0�)
�+%��1edʕ�t{';CJ�B��t�Ԋ~?w""��T��蜪W�sq^M.޼p��jF&$�b���T���'�T媞X'�W3�g���r``c>�0���[@����o���\�[tf�:u��")I���H5�g[fvn
�S�D�W�8��o�����܌v'�.c5V��d��(rt4R���F�60v�W�.|S++����ma��T54pDա=Z������I�P�&���R׵>b��)�cT�m�t`B�NC�������irf*�����%Q���:1b4�]�-5c�Ȑ�%f�W�h��߉@Q��qqq�9 X_�nL�9E`&�D�lJ�B�0�z6:\���^#`<84g˞��ft!l&�{�=�a��LOe�!'WCca��˲��� ]A�̢s�V�����Y��������0iۂg3�R���Mrp�Ǯ��F���),w�5�[Z�b BAA�4��-�����]�a��5)"�|~�Tߖ���
EH_4�HX+�ښ!,Ȱ�X������g0�iRoo���@]ʐ�}�^]���a�ffF-C@����+��i�o��#���Ec�bN8џNՊ��ܻ���y0l�"�_���$o�SBB���hPrr����jz��]:���4��Q�:s�[�3h]�\ZZZ���ɩ�ʹ��ZGG�$��]mn<4�$�@��/�ط��Ez���>W�����.'��!ϑ�;��uu�\,ƼX��cL���g2�v�|.�>[��:M6�h��Q1%�P9LL�b��Sz�ح���»��K��#�^nE"�����'�|��v��� �/�����m�����.c���H�Z��Y�Cj�<M���"�zj%�Ez�#h]���g��J��Yk�[or�N�zsㄣg�Er�T����^��'��T�xI��H�-X}f4Y��T��,������4�tB����fM�Z���t2i.bh~?����>]Q)?���٫�꠳k����E�4]����k)�‿�s=K2_-( �) +�K�"C�~~4W���1>�ŗ[^�rrm�b�}Cͣ=;�'5ؿt��)[<n̛r�����yg��ݡBX�;�Z�'keeŨ7�5���_�{{�h�e���by�v�`��2s�70��77t�M�67��9W$��v�uqC<�i� ���G+�JL:�i%���z�/�f��հ.��8�[�������ײ>���{"�
��f���/������C_]]]���ˬ���"���� #�6���/U<��,@�P���+4db��Gfu��L,��p�S�sݖk����U8�#m|y���D`K�A�[��9�F������%������	��16N%<���@��^[:�e���,�I.�Q�X!y�Х���#j\�g�Fxh��ڧ&=N��S��E��M�Oxɰ��a�M�%��B>��1���K#�ҕ�'a�o!�ѹlV�4`n�9mVa ;nH��K銴���̲���v���!����2_��s����tu��T��l@p�z6�q����*�C�mz||���$;ʐR5��z�������p@zz��������YLQ������N�m���������L@�e�W�8+���E7���o�!߭o�/Zd�b�9�
����\������y)���1`cQ�w%��X=n�V�=Ջc-/9]��f�'����lA~'�戤o�:m��؀�~��&udU��VV�q��[[p�:���@kܲ�v{� y�?g�mvvv>��ė��IB5�%s+1"��&R���I�M��p�k�/\���o?��,>�k2�K�j�lQv��Q���"B�T>�����ƴ!Y5�֞�a�����C�7��y��ȸ�W&���M]������^��ʫ1�_�W7��ny��g*@�U����e��ned����6�MVT�F�j�S)(dhc������yN���RM~����z(�']I�&��j���H���	�w_��%�pݴS��^�,+�_[����CCҟYY�g@��n�}2V\��Jr9�S(�H銹�(�7j�qgj�9-SW��G|cM1�W_X��.� #�׎�@L\|(IH����BYYy&�nE47s�YZʮQ���{?�|���p��vXR���hp�R���VS�MMMêTM|.n�ئ��Ym+1ӿ+|�0�Bٰ{���섁����q ���|c3�����4h�Q �c�'��&�D-��K��q�P��{�
�$((��Y-�����k���Ԭ J)y�>?�g� 3Q~*76=����i�i�rJ���wfQaa���<���i'�%/:�e_轻'�oea�@��������+`{�X��J��22z�>ssk��ހ#��Y[���bJ/�ž:���\���zx��!o��f`�*6΁�[�S:��+�ptvn���� �6O�������O����	������g�R���C���b=��dc��l�z���#�r�HR����f ��x��h�g�Y��s��"����e��`~�����d�N^��쪘��7]">{t�;��4���RRByxLw�h3zܝ��>Y	�_�b�����kJ-����2�6���S4/�Z��R2N��r�P����j�	_���\���飝�������+dI��x��ZXm��9RӖ&,�<^�r{ܔ�	y=��!��*c�1��K�X�g��#A�i�b���.�=χ�f<F�X�v#�D�n�?�¤� m�3<=�������������:�']!WFM�ε��aW�Q��EsrIņN;>v"�&C�Ʃ����N�V�SڙE@��  |������(���1��2���X>Pc��nc�t��ࡽ!�M��0�?�>����@�m�v[��D��!/�<	V�46����G�����f(~��'}�&X2V���Eb3��������=�6�gf���M/Cn��Rΰ�zw�e7���x˲K U���Ūc�mǍ�b�����3
{�M]e�x�T��T�Hk�PksVf&����Po�rm
l�SG���G��{G�d�Ѵ㗶����W��X�_�l���������(d?'šg�_���K��!���W��^yoo&n��!������Y�].yjaa���9}iplk��,9.-&\��*�MM���$њu�@�7��+,͘hT5���_��Aυf;::�\�I���`�D�gfNA�I�[� �r#RQQQrr�)�"�6����F�?@H��/����kj��C���9���gpyD��fT�:Գ?���T�B�}x"�2�"���J����͆.lNKc6 ���4K�O𠮵5B  Y1� ���~�\펠���me"^ؘVH�Y� 7�[���b����e�s
�U?9GzV�b�D2��F'�򟼝�D��pY/�w<+Ռ��l`zu� .��/".�d��?�H�rgtm�R2��P��XPX���w�6@�EO�2��D��=B��cέ�=#�F��d�s\_>��XX�I���u(�����i���Q	?C�Ɔ���Jr������-.B���uk�W8���Yoi��B�����)�o��B����!�U=���1H����r�;]��Q�v����-�n��=e=���Ք�1}�o���3��z=[o���"	r;�l���B��;���5�WN)�sn��j7\\_��G�jj�wB������z�.񧥻(��5Е���}�꾸>뱓�c�#��g�[P[�ZZ�(��uY��*��jxߢ��6zE�Q�R��-m�\:�̃����\96��0a�Cm0����;;S힮�O���F �]�@��"�y]��Շd3���|q��vZG��������hw��;]k%��wy*�:�
z>������y��q!e]e����"��/���#_g�a]@���ǚ����B���4���)( ?����� U"
�`@"�Ԋ/}'����W�72�}�ct��(0\��v��3��֠m��#���]Xs̗��b���?yQۄ4-���-�dǛ���iv������&a���Y����y�҄L�� �0A¨�j�}j��s��8��z��^�}��ށp'��4j�����w�������Iu��o�qc!��E--| ]z�Ɠ�������!���G�D� ������%4�������wT�Zl�a�`?�uû��E ��bȓ-�r�h��M�ꂆ�6.�Ϻ���̥����QFH5�(�虱��R�Bݻ��バY����Tơ��݇��V�ҟS��y.�k��{�����S��Q���cH1A�9T5Meuy�-+�b��`:{�Q���`�D�6Se��`F��>/�;l0)��4C���>0M�����
���Y�JWq%�(�1�o���P$�o��g���ě]���;{��XF�0�%h�����b��j¥����<����,-vB�=-,����bϔ�ko���-��ֵ��h"E�����3++��@-f���H��k�ncxŗ��9{Zv6Q^^�d��m���Q_��˃}���ϭ�Rt�a�<	��ݔ�1���vh����{�96܉X!FN��*���j���2#�$�J2��O��8����%���:�f�///��;������Ͽ5T��'�PV��u�k���n�;{_�d�d���'�`��l|000�F��j>5�t�6������Es\"�N�67�vH�/�L�ei#++�3�|*s�ƶ�8X8��YYl�1�.`��4�[\*��!{z{Mƃ� �l1KJ�F�n�������_���|���/..�h)�%VK:�BJ�DP�i-h--�����]�n!������J;�����p�f��
�{q�M��VgKl� Y�#�O�}|�Ͱf��;��G�	�������͵޽B�����RZ�2iN��@[�'@@!��q;9�4��:�8�����oX�w��BO�����.M����X���T��QS7��#�Ӷ�Y�խs���}-�ˤ�|�դ�4�5�HnJ�T�)��8%�fp�m4)4��lp�)��c��['�'�1^<�M����Nq������hҺV��ZM��4��- �!m����!A�Og9h6�~�S�΂rbA����6���L�V�A��͵W�MU���G��qIkh4�ʊ�3O��������P���C�&����	�<l������h�jN���f��]���O'�l��-N�����Nu����p_ku��v�Qr4�� �f���?�d~���䐕��gZ�QnP�,�V"���D�����^��@BB����;������O��I�ʋ)� E�"̓96���q�3}���]���J<|d� r��3)7~���
����5z�MOr�(�T.�i��~Ç����X+Ù�@���7O��5׫��0MPU������g���H{�� ���,Z��x���s��~�Z�99e��4��W�p���6�!rF�}?��]���z�Wk2b�����J�����������ݽ{v�k��Z�khV��뫖U�9�>�@��0>���)KLNk�s<C#п��[g��E�JJ(j��)�b�֠.���&a��x���?k�C��⒐����ذ�G��uH'|�<��!�TS��i�7H�$g~@e|�MU���{�[�5���7�O��y���6�PL�V����6������y���(_vZ/���:��<��}q)�Giܴ�&)	�ʨ�3[�j��8S��n�2<2���+z#/q���Sh檆�C�C=ʈ�!���dzJ��  !H����n��yX��<++�O���TցR����.��_O�^oT_vb�n�$�� C�pK�,'�|���I�s��x 0�֫�m�����%%�y��U�u4#_�7��C��^
v�ھ���|�a:�Aq���j���L����<�*<���Y^CYٿ��}4G��w����7�����zBHk4Qg�Z�fǩ��whx�I[k������$
�r�J�^�)�����1*���{�S�?{V%2""��������1xp�D�eZ�GC<�%�,��&׫�`6|�9\�|�*/,��WբV��!�����A{��h�ʃtzp�a0d�M��?��`ljKu]���q(��n��5�%i�܋Z��=b�v�t*���y��̐�K��u���|7ԀO��	����?����7������3+����ō��C��@WW92���`f��*H�{zT���-myN�bJ���rh���v�^���s9�+���31��H�V
D�DdI�P����рjYm�1����@>�#�LKUS)���W�|ӎ�`oց���RLB��3*aڢt���{�űX;�4===�ߝ�����L��yϐ"�I�Sgv>�����w� �ɅI;;�H�	��ǳ��XN�5���qA�_̬����s ��e��8>l"��c���t�)������@s<4�k�(���ߟ�ύ�nKJK�˼;c4�Honi�=�П>��#����<R4ڬ�.h����pZ�L�����r���BEE���ly:��$&�}a#U��^��*R$��M�InL6c�S��c��,����j��
X���?[��G�Z,��b� ���Rys��6l@v���������UO.�urb/R̉��V)]v�e���U50��]��c�|x���M��35�!�hs�Ծ�K@�����r�� K����<�(М��|o����=3�y�yrѻ{��Y�R��bѹ��¯���Q�#*�Lr�C�Ã�_@��0��/d%�]Px��w��1H�m��
]PHHP!���7�3�		��<�����o��ϒ�0=3�"Ȩl��D$�w�g�}����	���K2����\@nn���- �7_Z� إ�W���-{d[�VP
?;�B(K�8�>�+�svN�� �"�A[ZZr�UWb���f�5��~]J���!@���B�Ύ����p[]V������L����ũ�V]������ \C;*v$_]���p����ڭN�dQq�
�Ja���@5�����7� uv
99���d���Კ~��R���n;�����]Sy����Fd�T�RY� Pn �zU�����9��Yh��
8?>?~JJ[k�nt�O�q�	@ϣ��Ѫ� ��,,z��������_��NaՓo��J�z�
���s��@�p��~~ n�!�b�� �o(�'�� J���j��;7A�����5�������`M9G
#A���Ø�,rgNGt�Lլ��hz rW�p�herr2�=`:w��?]_�Ѡ���b���):+j&P�������By����>�*�엤*:�2ˡ[�^њun��c?{<0լI7�X1�t'c��׆����j&7�⃋���l��_����_�>8E�@��Ȉ^��MRRRqe���==�];�[��l�V9��*%�f= �q{� �"�>�^��Z���|w�ei�͈�H�(!'�����◓��#��j
�1z���<�������#<|��㵲�6�3�(����IUҊN࿽ԭ{զB�q0@}B��ic�5T���u��Mگ�U�v["B>�g�g ��I����������5^y��2�P�}��UЃ�L]��L���\G�i�굚���]l��QSCt�@���T��U .�2�&=m���}PVV֪�����(�Ŧ�OcC[#��R���&Ϸ��'"��������;���Kc�r�,B�V��������4Y�?�H�+����u3���5t�d���������8ŷ��K�L����L����O@��8���{p�HR�Ԑ(̭�+�����t��G��P��J@u��6""��Y����H��
�fo�����:���~����eC���꺸�<, ;��s���;, ��TO��e�b�O�vt��3��6�{x~�U�ځ�~�/��<"?'�Ċ�V�f p�þ%������On���p���O� �.����:�/k��<�G����Ev����/��Uԧ}����������V+>�}�8�FKI�揬�B��������nB�Y.W�1�˖�J����CxMLO����0��TU1��/(mk�+�����L`b"zEeen����R�jjj�/_�����Ҁt��� dG�Y����Wff'� J��5�K��YM�j+� z�Id�ng�(�gyq�ka�/ԨC**�?���Ԅ���%��D�D���� "K��E�f��:����+nmų�����Yyqy ���QЗ��*cC�����t�&�3o��to;�7�z��2��,����(�����N�t���{������S��;��B^�5��g����G�z^`����FR�ߢp�~�]n������#�������B����O�2�9qw�պi<���
?a\]�S}�*����`���L��k�Ө�?^�2	�����A�>��_,90�����!l,��E����.f.�Ts"�3���;�����ݮ��fzӪ��S ���<���(NsKG�ߙ�ŰPdbR@��G�ãU۱��:��Y��8𽬼<>;;&*
���2�T��M�������I�n��d�A֚E�k�^���� 7����h*Oܡ���k 	��'{����*��p4r����ǉБ��h��.@蛛�* �}�A%$�(+�A���_@�m����d��i�R�F��!�n;�(�� ��hq��T�zd�r8+�F!����U=5�?H�qX��a|�D�B{�q�uz�(  ��uu�aUu]�ߤ��4*�����4��4H���tJJ�����t��-)- �"%�g����y��<!��^k�q߿{�9�c���gc����ſ��[ޒ�9�0�~�����t<`����5�Rߢka'�����ohh��s�Z�`���gig�+���]�7[�`o��뵁������!�F��<�������xM���m5��Ĝmg��`���%��6�a�mXetR������V�������K��z��wc#�W���� t�u�:�A.���|����,�55]Cbll8�B��LLҕ·������Z �(�P����H�5�>
��]~�aCP|��[b�"+�\C�n�s�NV�A��1hD���`��{	�������y�	����_�>t	�x-�UC
��pN��^��@��_�GN�b�}�@��k��8�N�eF��P��&����eyP��Yq��o)~4�|����c�MJJZ켡�Pt[$Ϫ%�ǳ����|3��T!Us<���1���l��ͫ�؝e��>>R22F��x��b�ۨ/_�l��У"DN:��jw{�dM�� ـ�x��@��@�y�L@�P�,�a�D�UJZz���w�r��'����6�5�|�����x).NpT[�����t��'����aC�������zs_�wpl	�W�&�m����ݸq�;I�RBB��z/5�����_�����^��ɚ^�����f��G-�m���ѿ.�����m���"�*C�����������CK5�m3Տ��[ᚊ�*�������N��/"w]6u3)'�]��]�������E5j�`��n�}3�Zg:g%##���Gv�K��� :�d�/�$�Ua��Wb�?���C�C3iȪ)Y�;�WQ�݈vvuQ0�	�l�A.�wϷ)���Xц�r'L^7�{���>���d�w�'��&�����J�^^���F%Tjjj�8��<G�n)dv������ş1��өYY�����}�b����ej^^X�F�ȏuT��$�v��svx3���#�����&�fLKC�,i�����b�R��q���ܹ��Qs�5U��h��}�/°=�ug%�-�; ��Re.~���
��3c�p&��k�L:�A�n��0Q�C}���S�����i��E���ztq����ODm�lQ�hO�HM���������S�X��~�6,���BZ���R��P�(#�m6A�L������3L_Y6�GIc����4O��B擁׷�`~�iު�O���VWWWx���-v���ɸ������2�z����B�5�&���44���Ώ|)ֈ�%cA|�2�=�ۀ">y}�[�q�.�F��p`����5�e�hi�����3�nҫy3]�/���m�����\�O�188�J�}
Y�W3��;�a�����J�e����']���]�����}��0K������<�^� �}����N
L,,&���V��z>�7���W�޺�.�hn^��@��f
��BCF����f9��`Pj*���x�o9����Q#T;�)w�g!���6���w��54F|�]\ڋ����2z�q?�2zlo��=x���!�ըQ5d�H��Uko�������%1�L�������T��	]9�-,t�J�xsr�"�n6���!^��E�,��ژ���K�&��:��*Gٹ��8��	W���i�����e�T�b��U$���@��5$K<d`um/.[̾��[K`$"+�	���q��ӗ�b��h�j�]T��X�8=ς ���V'x��C�GÁACM-�y���Cy�7oݪ���q�?�:�2]��IL�:�{��0ġ��k|Q�	�N��ے}�\ ��"~vv�s���nf\��=+����~ݫ�� Ҟ�?3]��[kK.)�y���v���,Dɣ#WZA��\I���R�KeV��37ϣ�`�W�"����l��>�n�$���Ur��P�s�?2Z픧��ѷ�bo�c0�I;k��qU7����}A��X���ɜ��"{9L�>֕�zϷ�V�5�J�͜��!Ѳ�֖����7��}��^��nk��y��ݲ�'Oj��� )1eYK� ��'Q�+m&3&�b�6�KK�"=�x�2C��|�Q.B��-��������P<d����Jp|�j
 ~�җ1��S��!-r�=�[Y����ڋWR�6�o�Ugnx�-�`��u��ʺ��9��+��z��
2]Q�uZ>pm���ݬ�������MH���ݿ�?�Tz6N����â������%�$���ͳ-�K���o�x�i��O��6Pv��L�.�v�V@�g�3��Jŀ��=#J�D�$bl�F�=��
[�ګ�괂֮K�뢢�jkk����|��H'�yO��s}��V#������[������GKq����'	���{�d�%�����箢��t��e�K>z���zki	?p�F��/���Լ����Qۇ��vvw��,1d���\U=s?�=��H.ꃉ�x�8��Z'9W�ܳ'z'B�7�b=J��� A5*�}g�=�|�<�H���	2�Z,mk���v2([�Amg�S�0���,�))������GƯֵd�o�����[̉V��ޏe�,��h*|x׉�bI�����Av�!�N�������ϡK#.����HP��
���p1ё��l�����i�qg��	���=M''.�ʔ;�����%~1U�}����g�h�./.6�n��yXl�. s���/�T��g�9+:i뽿u�fcs3F���R4��h�!���[���U���c�"Ꚛo��.4	ߺu��$��CJ��R㕥e�y�WP��>g����Nyr)��� ��!1�n�_͗/�VD�Ē�AH@NN�>�x%Ge@x����A`���Y��9��b����~�\L�����,*���H��~�[���>Z��� ���V�;H<e��@ .1E��J���;����9Mm�R�T�F~��ҕ�aHTQ�WS���Q����O�c�h|̄��(	eeЀG��4�͙�&v���t���f���.��*� �jW��Qɲ�!R�{�nDߣ��m9�dhm�d�������O�s��W��=�dNkni)�t�?!!�	��?6��s�o	����`�%b1����}||�S������N��L���H\�-��A�BH����Vu�a��O�[D�{$S�e���p��D�=u����~�YK}��8�n&"���٘r�U]�������+�?oޡ�&�mf%��`t-�K=�fr��<|�d��h���ؾ�Qd��R(Qm�Z�;�髁���	���s��}W��7Խ����}�X���+]�;	+��������8<�VVd���2�=ל(X�I �X�P�,F��K�"/p�U��X����FާB��@���8�_O��C���'0&�,h��8�ݻ�߽����A�@q*�������K���e��k̍�1��u���N��'��Oٸ�&CzMM���뢌X�{�^�qy֭�&�s�8����sܮ���o�����l���9�]"���$�kɺ�.��R�-�W3sN�(}���J�J#����l���H����h������l��R��v&b�p�L��_���ٽ1Z��J����鈵��'N=+sB�;�T#}�n���Y�Gc0Y��P���m7��2Ey����MRC�fd��-�:m�"���٭���+y9?{zZ��d!�3��Eh�������������f���<@����D�SSN��)���333���]ԍ�q���H%ѳ޸�F�4��9�qb����ܢ�Y��!�DGY�z�kׂ ��:����mm���è�g=a,�ŵx9^f�n���g�c�wt�=�Ӄ�ݕ����?Ї�����},��+l�,<�;[�a?�d�R��[�Ц�"��[�Lo����Y�NH{�=.�L�I@�H�Yȶl�z܈����{�a̻\��֗���nX�L_+�j.L����?�����U�c�Ƹ� ���`�4o��ఋ��{c��<�m�5̪�%���f� #26�#,s�_f|��.��y��+�;���C��NJB���1�lE%h�{�dg�X�NLN ���r_�iX��D��݀#_�w�cO���1R��]˙/�'	z8�_�/����wTO3#����;�$������iҷS�{5G5h�4�O�
�����E�Uǁl����L "l��\�X�MZ�k0�z�;��#T�Ԥ2o��y�y������ܔ��R�*��"�"���w
�[[s�<�ӱ���33���W�gz<������;�C�%MMM�06�K�ϓn�* �I���D�edQ���A�:���{l�r�:2m��ؓ�i)��<����(���.\���L��Mx����I��;,���3��|R˻�w~vvχ�Ν��E�ˋs�*�[+�C�	|�I�,�,��D d��Ǐ�^5��[�u�����_M�B-1��雟߉U0�=H�ԭ:h�}'�L�]V�Aa]P�+��QS3>�����h6��R*�M&ZN5�09���*<5��`i	�\Q�Glj�f��;ޗk7``�q��OΫ���Cv�bbb�.��"��é���?JDX�I�8�𲦿��I����K#����oZUU��_�W�yv~� ��m�}���K��p�n��m-))����g.6?I�Z9�����&�3���_5���Q����?~x���x���g9�2�Dl�������X8ϯ��wڜ�ʛY���H��|��Q6��rQ��%���va��
[��Y"���I�����'�n+�ؾ6�!�߿~e.���8f͊v��]ه�#�.y������F�/#>ff,d!R~fl�3]��kG\TTH��Z�6k ��C��m0����	�;0�9V���؃�E�:ߡF��d#��l())��2K������ê��CAҿ�Z�ݍ��i�{�o�{6DI3===^^۾�ۦ �J�+.N���f[��?����l�q���w���~���?����3M_�>l#gee-7� ����?�r�֭@B����3%&K����sM�e�[gǻ���aa	���2�������f[��c��AGX��m<C-O=��6q������f����<TUh�իW��bb>��>���5`�w����Mp���?
��!���6[Wǭ��U���H���u�ۢE�N�1�=��~h[�6��[���3���l����Aڷ{q�?|��V4�P�p�x{f$��4d�W\���D/�?>�j��s��Y��'r7���҉/"�²�XkW"��<�9؞{t������I�h�>%��F�����M͟~~~�@ֳ.�
�W�]g� �թ{9���*(��l�����[ޒ�~�2�ɧ���$u�98X�[����,Z_��t՗��7��oZBbH[��x'���G�p��8�O٪�V�MPs<x�iXc�Ov�!�q�v$�Un�,YQ���f��������*�倯=����z1޸qC��³L����Z�Q0U-�d�˺�P�ˉbC���̓m�9��C�*ؾ��4�L�/GBt�222�33ɀ��&-T�O�<4������)��Z�$�u��7�����
�S��q|�Y%^8�?�C�����Ez=�� �p���\�BrX�y��۝��ȟ�=�N��oDw��j����0����0
FE;�18�je��9���+y(���m>�[���Ύ58owk�t�F�p��x�З�ҵ4�ˋZ��ϷlgD���=J}��ixx�z0�qm��RQÅ��9t׃�p���b����`�R���#{{(>��v5�O��\(��g�Ol�+^� ���
�3"u��)�t�4���d��8�K���m���G}�0F���暃��={V'�c&U]Y�sq��@��Ä�Q �}&�Mw�YQ>�^��	Ī�8䲭2{�v�1I�������plj�%/�p����"��85��":Go�KU�k?/!z*�}�1Ӑ||r�M9��Zi�	�]��M%��;��VVy����^���������=+�O/;y趽���~��d��J·֖��>��pB�l	}B[��P�K
Λ�U���<C^��u������C�+σr!h�Cm75��)����c�cd-JO�y �Wb1�Y�}~B�أq�w}���3��N�3���2�ַ��w��?!Xc�(}R��p��qy���C&|V$
Iq�N�V '����O/���#�S�\�k�33�M[���Am�u@m	B�+[��r\v%xDo��oA��ܔ�vv?����i�'�}%����}_D�!�8�S��"��0 b]�o�J�����zr�����W�OWw���4�۟�x���i����w�z�U��;A4�?��NOg._Ew�%���{�~�y���S��:`h�f?�BƷ�8�<S<&�cU�!_��ޟ�0iYّ.����%�Xii�Pd111A�#���ٔ���R��í>�'_�A�F_ԌB�Ĥ����!�}��L�g����l�-F�ޱ����WS�y4{�A�lƾV����G\ʥ��Rf׼y���?�TG���$Z�m�qPE��ȶTAf7��:��2�0}���_d��}�;Y�X;R�B�������8�l�{Bk�q���N?�'�ݨ1��Gs�SfIa۰�>������9�ZQI)�f��h277g���u�v���7���ԙc�#酿�>
���׿FG�}��A˻��ם���Om'{k7�֥�M0\1���p�^�h����(�� �Ƣ��2�|2r[�&�|�S�ܯ�����|U���Z?t�C�wc������gǎ=2H���ظ��QT���MM�(S�@��mm؂���eeg��''k�|4#1����mh��Jyu"��H�xa�����+p�
������C �o���f	�=}J,A���Z�\KS� tٻ�HEV�@��HQQQO��"g�|���q[x�=�r"2�aU���48H��5���,pu����4 t� �m&��W3���A���R���!}�$�(��G4ӣbiȽ(d���ܲ̕���ܵS7(�D��%$�lV�l�q�0�d���#��Vb\�n�:�Y�g?�y��s����8�*���%`��y~i)����JDP�W�Ɨ]E�������[����o��K��H��y(iiiKm&��Ѐ
��w)QɑRR"�?���[冀��C�H&���DlD́�ܞ� ���-�dQ���أ< $�G��R(Z��!p�lqeŪ��4Dn�>���ya��jܜ|o�R#v��"��lSvꯢ2�vP�C����Q��� ���^k���q����&����j��ʇ�n�[l}}��A@�v��!�ɾ���V[%��v������z?�vr�V����&fffL�9�;L8����W�m���v�0����IJ���h��j���`�o�SS��#��߾}���7���5D��0Zb��}T< 0��b2W�N�n��������d�
��=����;��z�}�s�ea��ۅ��Z�j��j��%=r� !S�(��d5�KQ�	��W'G��	���:�������������g���I�$!�Am�Y�L�
l����'�^EA��0jL�����l=��p'%#�[_cq7@|���F��bY�^��s@Q7@ ��s�p짻�/��^6N���шqR$t͓�����H���������q]�\y����|�Cn���K�I���6�}���n/w*�YU����ѝ��LHnN�uY M��z���d= �Z�bѯ�� �:�ʹ+�yA��T��4S���ش�JTƕ���G}���i���w�� rn���'$����ޑ�,wS��� a��M�i���3O:ag�c(�]�.�� ��Sg\�!�f�����������v�*i_Uo��҆!SȐ��ø�ấv�c��2����H�L��|�F����Z;��mLT��Zή�\�c�*ZE���SS�$	�~h�T��$)%+�<2R񭧫�-�"wA�t����z�A���/��psȣ�陊�2kN�8>59y����z�t�������*Gse�F��&���;wIH�������/�*���$�6TVU1ݽK�L��8������M�?&�����D��\7�F����j}7�)�U��[�r�g������'��%4W&g�lF'&v�BB����ז'��/D��2J����@�!3����V@��$*qK�����`c����ݠ��l��$�r��L�Lk�����kc�Y2�������f��U�������eZ@��.�	a�����(�I���ǟ]O2T�ˬ4z�K����@:o� �s}?~w�o��y�UeC"!���';��T�ӂ�y�U%��o]���q/�S��l�����\�i�2��ݑ�=j����&���! P�v�|��Ѕh�S�D����>�l�]å�777�}R�]�mcfe��������r-���O4?�N�@��*��ℬ��CyfUa;#cgw��y#���\���j�����Ȋ��ty��@�`���/ʱWa�+W�f䚚NNN���pQ��[o���F98����/�(��&M!=G�NT�?�ocff�L"�/פ:89-�ݺy�).S�V���ޞ��ޖ�B{e���g�z�@�e����FGKNn�~��Q�KV�I��ۈ�@��r�0���9���d����[�"����D��6�,��j���a�N0R�	�#©D�U��b����P=�D���[\Ą|���y��m<�9�8�"�-RRt H�͐5���䶄v۵�7��xggg'6���ż��˯�O��ԖI}j7~����2�*����_35.��WI����3��vZ�ll�;�]�ֵ����]>%�?����d�����(<D��1J�K�5u��-�� �E��} ����E�P�c�@��u���<������vo}��
d��}��].Y8kdU����~�!Z�4�ׅS>�1�p�.gcG���sFU���*�����u:�www#�P����C�蛑���֟ �X����F�(>��Y��8齛����R��$5��؁���3���7���t�9�4g�'��AW@p������[B�j���?A����L����gMqq�q�����ְ��϶�c����Ez0 ����ȣS�8����%�V�����;�C�p:0 �o�򗻙km5Q^�|RH���S��� y����g���充��l���������斗e�$o���@���Aq��)��9:6�H�����������NJJ��N֭�CC��~�7��~��5S ��:���Q�׽��dQ������`FcCyZ��!��<��R����_����ȭ�;95���܃��}���H;=J�W��g��w3T:tNu'~�lR�	�[XX�zCԉ����d��m���P��[�j03B/R#٪R�������'U�;���nbWՄ���_@����M��"ms���⁈��!S�e@@��!8J%���Rg����a�����`�_w���T�m�l.^��k�W�z�k{?rh5�z�����r�$}&�Pb1�<������uۍ�˻c5��0��e�E��f�;TJ.YV�ġ��U�){�RT6��7I_�`���"[��l��{𠩷7��Jf/:!!$<�����1<Q�u*ȉ���ڵ d�>��uP��,��}����ik��1-�uu�̃�g��l�ݹ�>��uY�r�OBR`�����e1�TL�	�9���J�Ќ'�}cs�������e%c�%�BV�m ���P�z�Ҷ�F����z�����h�H;8�FMr��@U��H��V[���{6�3�b>����bL��ዚ�&� W�=��+M�螰p�l������t��66/��M��oܸ���� 2�lOD�gdd,�+�q`˯J�u~�X7�nG�(�z�U(��<�ӧ��l��>%%%�=����j�n�����"���F��!..�����c�����'���Fg=�H�P)#cU�.,L���kX�z��n��U$��c������
��h��r_r��~�3�m���\rk,�>bpsa�?O����_5����<r'e�-B�Ҏ)�k(W�LI �Ĭ�F��Ě�� [��oAfff��V�Ӑ�����O������P��/\*]Y\4��8W�473İ_t����ʧH���I]��,,,H�I����@.���9����@nX�:ZLUh�[㢊��}KJx��I�f��@�D{J�/.6V"GաM�6��"��0h�	�z>.�)|�|��a��D���qۧ>eC!��+�*�+yQ֠��~~�f�^�,���+I+=~<�hU���C�S�0M3\\���h�T�d��*�H&Ґѿc�To/���(v�"�p��u�u��R����p�^C������_2���[;r�x_������C7�C��N���t��g5���cab��EE�&Ø��-!"$\ڿ\I��-��8Z������6�F����߼V�R1�C]���o�c� �r�8�_��7�*�]�&�^gN+r�����@~�|��$*�����j��!��sXġ����j ��M��o��94��:�伉,vONfA��P�������b7Xm�U�s���$_�������Įqz�ˠ7�1d_�p�e4��b���}�zu����j��Lr?�Lո�'&&���%��{OL�B�+���H�U��(~d����%	�����f�/�\��0@C��*�&E��&֧9�ԗq17d�M�P((*��jBa&���p߹sgy}��K�^w�t�Yx�v��ow��M�X����!Y��CF+��א�Q4��GN�r��ꔧ{1Vê��Q!!��Q#/��22n�@����[��=;v�z�lyX�Np�^�]���oQ>S��Ѕ���V>r��`iu��DCq�SV�z:'���>�І@�"7<��F��$�*�D��z�q��f��2���:�>�t��?B�Z���+�o���p��y�N͇���\�&p0�	� �����b�F�
F�=ѓ�&��H"�SP�tvLWa�^/���2@f�휜KJ��څ��Rʫo	�C�u�[M�~���}ں΁R �Ĳ��]�w�>�X"1z�������Q{~0Q����L����k��_��a�?��$?��*|!L@+H�q�j@L�ɝY��3G�����׸t�R�;kjkC�F�w���{���a|����:i�=d�_o��d�����m�����Չ0<tM4&���ÈǘM�H,�?��(�s��>p`��̬�07�syk��1u'��o�Ќ�C��Ɩ0�x�
;{N������x�Ӵ�x��Q�3bw��5t�m�+�CUrL�}�9J{<||�<<<�n��%�i4�{�F2&*l�XY�h։�Z���מOMM9]TVX�����a;�������?]��C�*ө��zX��j����6��+�W�v(�R�9�R+�z�����[��=B�qri�Ü�����۷� �C)���N>;���j(���	�G��p�	�: ����j�L���XX,���� Żzx�<X+�r�ߧ�7x�5XNN77c@�\,�<"^���8�c�>ۑ�;����O�"Z�)�)��x�f���6��	�u*q���kQ���NNj�5���D"�z�4����(����elZ���)6@��8,�${�e�L����Y&Z_oV���,��1�������d�А���gI��� CzI� ����f66C�N��E�Ē�ee��y����)j�`�mu����d,J�ge�0$�It�Ψ	�g=��e2�|)P�(9���h��ɪ�||����T999�ۚ�]n�e|���^4��kU������04���Ke�W�����^�1a�B�~("�<�gD߇^YY�v,\ymm��~�K��ٺ�6��C���F8����ls״�}�/+�5�SL�Q�e3߹������%r
�Ԕ�VNYY�?3���	�>5�(BQ!Eb���p��Uq�ByE�����������ݐL<||�X������E�����v�FFMa���e
N�#�n6�ﺭ��Ժ���Z��ı���bN���W�e��j���Q6����Y1PHk�OhX$�AK[:�q^A���@�8]ȡ��-e�ð��6�h�i�i�XERN>�0����]��r/Z�5	fs�������m�DM��-�^$����+j�̗E
��=ّ7��k�����{���-z�Ra�7ؓ�jhJ�쾑�߫\�g�Q:�E\]|����ʖ�hw�}�|�Q�pu����0�+��2��NQ�t���kKwh|�P�(;��k��C�8is%�P���P�|�sy|+Ўз��:���8�	*���O����G���Jh��� �jO����1���S���(馏�hn�5�6A
w��ƞ����5���z�EL8��+i���FXI��Z%B�Q��$����m��_gc��|��"+���b��>@ɠQ�l������d5�JcrI�(�|*=|jj-v#a�J�9�A�俧f�:�Jc v9�Ё�O��a	ĞI-��K�_$D��jS~�__9.V\ ���r���7��$p-Z�C�^c���dQW�/&p}sbI������[��wSv��YU����=�Q�bRKEsx��8�����FY��GuQ��[����^����o�=W�j���+7�6�^�{�����".P�K�j��K�G��ίߣ�?yie�BI��PK   �EX-t:X ~r /   images/e121b57f-ec89-4d70-aa13-01e52b785a2d.pngT{XT��7!%�
���ҭt#���]" JJ,����������ξ�{���}taϞ3�O̙�뫴ȳ�O������
���!���!�"����������)�����O�;����=q���TA�񵃐���������!���3��������!���q�!7�[81�/
.����w�'C3���
~W��T�n�p٧��g�W�U��S
1H�M�RdI�"����#�bPrv��󞀔�f�=B�hjϫ��Ж��c�vqiO�Tpd�qιu�d��h��~a	�z��	A���G%�Æ�Cu���-���UUeKI��P%J��[�����ʨ�T��>j�S�q�9y�",g�(������r[�ח�0���#l�7�qr�ơw-UP+�(���OE��]B���1������!�i�:�!|�7��{��.$�g�Ǝ�ɋ�ظ;�_#J*�0�	���9�������7��OL�]3�_(�|�i��0��)Dl�Al�}�9c#hK��,�J�3�0�6����>��A�����򕟫�8��fp<>�������9�_o+C�T+�[)�	ߢ9����2���Gj�3�Raߎ|&�ǽ��@�nK�9�>�����A$1�b�%��4o����d����!#X=�y����	ꊣ8�|��&.(.������xj-�Ϲ���}�[��ZQ�{������n�\Ό�M�Mrs�����J��H�pUu��d�.����s��F�T�z,ח��ڿCs>��l�Y�L���d_�%|c$;���#��f$:�c��� ��t;��!8+���d���o���8�k�Y���<Y�֚˿r¥��n�Z߷pV��s�Ӥ�rj�Ké�����r���U��v)����B�A�E�P���%��ax����c��_���l�\8�󳝜�0���P�N��{��J{ǈ`�����Ӡ}�fj��>��s5?�]NF�T������(o����0����W)���?�F�&�Qf��5(�hr�C�@������	��}��ꔅ����j�R0/���P��xxx���_�������1���]\\���3��˫��ų�����O�O��+*z��ޑ��[_7����������������g`�O�"bc_�kW�3����������>^^�:;����(zMccc�����M�Ĥ$1Jrr�o~~O������{�+�78�X-���$d���=mΊ�ޛ�v"���O�lE�����J充��x�jd<��\��%�rq0���ߘ��������l\\!��1����qL~��{׈�H)�F�JKG��Qw:�F�bw"O��
�����1���)�`�r���<G{G�������+$�P�7���惪�Z�M�(���w�Jdll�0��+�~��SZ�tU�O���s��d��Sp$�LDxx���?被@�;������gj����<�層�MzV��?Q���{�ߋ�{ݳcs�,l�@�G�F�����<�mE���o8S�����]n6bpg��T����mW����Y9^鸿���!)��Ԥ��.LFґBX�u;~�6��<��B7]��;��?�!�(#B�E`�`
np�q]�Jm�y%���3�����)S,�BE]ۛ��is�-��������4s��������8��l��b&"��k���A������,��V��ݶ��H�G1P�`���H�H�Q���fU���:n�B�j����5�B,��\ό��8�����=��������ۋ��f/-E��V��L{2�{������"Z~t��
�d::i6�ny�Ȉ�:���#��C٦��)�k�6�<��O�rxxxl�d��_�QQ�B�G�o���V��|-�!`x�QQ�����0� ��'�C(��R�gXu����FW��W��@��8�����ׄ*(�����I}DGG�g��61�Z�w�����	���r��t���^IK�	�����r���6�e���Q�"��t!t~���*�2�sS�ڟ�
¥Q�9^��L����Fz�d����&Q`II���KJ�d�w���p�(�>��' �d����R����6ӥ��wK��KK�;6�MLƃ�:m��_50�����K�������A� �iII}���LF�Y�צ9���=Y|�D�&Ѭ7 O��αa��o�x�l�t�ge%tI;�n�p�q҅O�ը�7��<��@p5���ИM�?�؈'��[xݟ����:Y�`��}����#L�b�%�����u<O~g,'L"&%E`*7��p�EFC�MYY��:??	���vv
&&&���~.RZ������@��Nm�����*����$��)����|łX&cL�EE�7�At����h�E_��kk�2��zzz?���89㧧UVWW���%���z>�.,,,��A��~����gm�B�"W�`���}|vֱ�D���O�mF��pI8�#�5������>d�N�}���ɢ2����;&�]d�7���D###��? &rt\�M�@A�M�W0a����n���|Tb<_1H��L\7�󘻷��V�>
tsr��?�-,*z���~��؜��m0�KDP�����5�=�@�A�u�?U���C@DL�TA@@ �e�:E�	3��'_C��)���FV�,D��$$$ْq���w+0$��	������+,������4��$��\���&���$	: d�T�<?��O��O-�UTV�~�L�����,N������*������lff�"D@���i<W�WY���������޵�k�kRo�MN��d[�g�V�H#r?�yHr�4DΦ��lW)����mS�/A�a�8����o(7���������l��|�G���4ӱ�陙8���Zv��c�B�/FF�b�/��igUV�H�xد^�D\ �� qwy�6�&p�CBF�{ 5��ɐ���J�&W��8��!����z/��)��w[��ߊӢ��q��*��)��zޚX-6�}�?>�؟�`�J`� EI�E� �1���,��¢\��қr�d�L�^�p_%	&�l:
���2�<9�
�+��u8�FX�<�B��[��G�$h������@ �����k�VBlln�c~��������O�?�>��~�j 1YD�έ��j�ϓ�1�W*ʿ6W�r%�7U��rs��]�A�j��	��A�e�^�RSSK�Z�*�jR��T�@ �%�y�++i�9�27�����?0���?����v,��a��Tۣ.�����p��ߍ���S�I�C
\��i�/JTkm�(�鋇���k=aS***TP�,���X��,����\���(s������}Kˢ�=��͝�<׳6�ڴ�-�!�3M�5�SS�'Sw�NHTA�y+Vn�:䌒;��yअ*e�Lx���f�T��E�V����w&1�X��?�q�X �cxz���������(*5�E������҉�����IhJQ侉jo#���򼆸.83�\o�if�1aLk�V���;#�:�����
cpr5�3�:;����@�I�G��� �Y��N�.�9-�x��oa�Ey��4�W�Y��a���#[�PJbb�k�X6kbUU�Gw<��oD~3&��[溷���J��/�Onrl�����߁°����|��@G�O�q��\X@�b��_�_��E���:AH֤}v����Xq9;jy�S2���'zk)��l�>����"��x�d�!����֖kold�	�[{{�����C'��٬rSt�0�ŷ4�;���A�͍b�>*a/	%Cdl��h�S}F8t<�օ���3#ccXW��k��ny�!��q�~���.�2�šGeb�~ʦ�8Ǵ�������߾>� ��
v��'X/��v�;���v�~.v��m��B�*��`��2��W�����o�ٟU�S����x޾��u�~<�5/99�Y�+��t�NƉO7��ED��=�~�K�[$�vi��S�bc��.���n�c�E��e+��("x�������l
�X���C�P��=��ɸ���p�*Pk+�G�~��W�*���I�i/����'��H,K4��x��C0����z������F�H�� ���������kg�ƅ��1�8+�2[���_k�I�V�J爇=����Ԑ�߿��G�ce�"�I��}뽑��&�iK�F�lSY~�:�%�!��2�<N����
�[w�Qs�����&��-3�Q���`����D�/��4ZuTWEp��&=A���'!�+j��]��):�7��K-|�ْi��O�������,���d������o�hU�y��'��@�z�xˆP۵h�,AA��6c��׷G�}@eªf�+�WH�l#�e���ޒ'
�A)֯�c�1�d"�ch�@�Ȳ�)�h��^/#r:Z��b58�]�p����l���n�A{���S�,l8���uK��íp���͙d+L�&�5׷�z�5^�"s�k�l������/QSk��g�0����c������0��w�.�4g�(���/y+(��r(�B,��z۸������S4��(�B' Rn�3�bu��$�ˈ�띬v�'��ղ�E-\^�eLJ@JV% p$���ڤ����L��ύ�s�C�O+L�$Sx��f_�~n��˱��ђu%ǳJ�m�����ߢ�M�,(���(�E�l�ŚA����� Nc�R�k�!�K�6�YVE����*gC2�ѷ�;����MmN �y�ɰ�e_���W�K�RC�<^����/��~�no��g,;%<�J)�;����gmm�pH�'m77ο�t����(*i��1�|�1z#1�\��qω�RF{�3�F��PNF��b`�!ؚ��~a��?�(¿��������~vՎ���e�O�\^,�)N����>���L�́� 3E�&���	͵���9��7�s���нɴe}��G��l�[d�����E,��'V�-3���}�x�#ex?����cK���>�5} ���|���|�|A��+ǁ�\�v��i3��qG��qM.@h\ǖ!��E�yӔ3��F������ɵ����λ㿀���'G��Yl��Ց��G��&�7�W��W�q�sh�IR#��64T�v ��XYk ��qwP#��������pK�G��cqC˗K�֬��'S�^<��Ͻ-h߾��Za4Ra,��y��]�?�L�m����&{��%�k��#o��)���4<��A+��j�&8��t����i���"m�/<��:����>5=3�3|��i�:i�h/�����q�A�x�O 'F3D���g2�[��"''���ޜ�ͷ�Ϛ侹�+��#B�P�!��s�X$����ֆ�m����t���9�v�-oB�K~��)+�ֆ7�;>�S�$.�M������Q�,$����!���E�i(2e�1d�UU,4��˭>�C���?($��F�Į�Z~�E ��LM��F�ȼ��BD������ԣ���F��|�Ĥ����ۀa�X��8GEE�p��_'�[��x�U
|��aÑ����x)33��S4P��x4�|U���̾&��:��:1REGP���t��΍T���[[�x�U,�>�1���t�{�/g��F��rm��t�ө�i�{I"7;�7�F��
Y,5'���{������KYYY�0�<����H5��]sZr)#%<JiMP��uڪ1@�� �����ٔ	s�G_0�͏��~Fl=^�Z� VK�4׊@�����������@��z���u�g*��(�Un��%�z���_� DD�]o�<A�L�� ��:��"��+���� {nvrR0�EbS *1�S�|�|6�F���2�;'b�蔦�[p0��*rV�8�B5Y*�����M{��K��N�d!��׭$g���A�	3�g{�Y��T�j#�AH!��uTNG�	#X�G����)�&&T�ݼ	������ݿ��L���g��s�@���iREu� �]@^/�ba�S�х�1����l_V)��EO���V�))E��U�W:`>xE7�Ho7��@XX��:G$eb�N��l��i{3�2�J)��H�����ϋ; �����_��������w�ÅŤ����~�H|�zW��y�
]FF�ws�śO�)�p�-�U4#��]���ua,8�D4Fs��-E8Y���R\^�\ܮ�����Č"�p���'��&�����ry������`�o�����M�l��V�NVZ*��ή*+c�0n�Rѓ�v���-	x�g�lQ=���v�����#�PZ�2)V�o�]��*uf�U�6�}iAA��[����J��%k�K	����x@z$��!����ü%t��T��h�=DlVTJ���6��~+"�h.-��L)U��Gԅݘ�gQ�pǯ1噲��A�<nnn�*3\�z0`�G�)��,�n�3�N��KJ���*�|>�V�����{�>��}9�U-�K�q�ۛ�+��U.�b��n���R!P��0陝� ���PsK�R�ꇇ��V�E&<� PPZ^���5⎙V(�.3 ���D�7V=��q��4rP��_�4�b�@r�o#
S���*���oeҲ�EH) �h���6E��r_u�Ҵ���-���N�0�h{8�74k�\K�D&KnE~2)��ae[�g�O���YM�G�8`�m�5�*MҜ]�����FT\|�1�[u+^frC�ٛ�o��P~<#�^P�x���kv���[�yF
��ʃ�}��X���5�mJk� �(�/w�l��Q�9�:��?,AAA��rn�3��R�mPy�d�a 8��3��T밃
�����@��K�q����L�ᭊIs9B�
��������w�lV�1��͞�{11��w��SyI�x�Iͪ�B��4��tf*X-�@�& � ��U�V�> Ւ����[��r>$#�n��������6���-w�---g����i c9Y�[k2���'N�ݞ*xM?x�t��-?�G񅥴�z��������h�7v~@��xn5�w}}]j<D,V�O
c�g��㮉��h�~�k�|��]#t;���B�f�%{J\��0�&<�c',���1��&<�N�`��_��B��Ҷz��0��k
d�J?���ʟ�u�:,�zp3�,��\��ut�Z-ԗ�G��;��� ��C��-�e�p|���Z�}}���G�P������f����$��,�/|&��b�3e(��Dߖ(�8Ir۞�.<	��	
ʞ�T������Z�.�V�����k&�`-}OOO 	Ara��'�u?�h�e��?��������pkp�n�ޚ7����_у���T-���N��Q��B]�%��MY�v����^�s�^�.��VK�,���_^K|��o�f��U[ʛ��/�au�v�����`W����OI�~ўV��'�����������W�b5���*�&�5e���[���Pӣ��^�ph�P�%9�F��H�i�H�����~�r�<����/�A;���K�@���ўGi���T �E�v�'�����~W�;֯�@������}.!!�$i�F�� �)\Ρ�"c?�v���d�=������Rp$f��[}���o̘	0�8;A�r�Ԓ����Γ�l�;��y��m�,���u�Y�A�h����ϕTS�x��_���r���۟.rA`�D�&f�`D5��R	��N�5���l�y�P��c��֏����p�?؊$%M�`��;,Z/���ѕ�5�nN7 ����h��>6h�6O���b}BB��jĨnlV4�z9�����_`���~U�kmmܑ�LZi��%!!�wP�I����,[�]C��

q&������9�qo(|�����L�[	����QN!E$�:��K��������7�~�~����zѭ���p����c��K'
�vT`}����K�a��
JJb��(�|0�O8О'k=��4O��O�v��2��@�[α&s�������}&<Lg�ɳ:	��(������%�>҄��3=3���u�;q�3���������~.!A::��UGK#%P��Z6I��m��G��l�y@CCà����h��=�嬠�[=�.a:�^�ή�X�1O���3��G�]��a�[HHPP����7�*P�A�`ό{J����������:f������v��j�=`���� YWG�$yܕR~��j��2��Q�U(P㎌���~�?u�/S��(��%g{��x8����B�H��zc���xN�g�)��ugYd�V�0\m�	Z���[��(=����bG/-n��dddO �%M����l�h�m�'v?Qyf��a3�������b����ﹸ�R�s(/��n����2V7LO+t�HOi��f!��2�/�F7��pح�.48O݌pBą q��S��&L�53We>���oQ�q��?]m�0�/c֞ظ�՘rA�slEf�»A�D?T������|+l�x���L`�*h����ô8�2����o�e~��;�5���R�03f�y��O%���0N1���lg��J48+�Ӎ�T�1�e����/���7��N �B 5�<nʕ�YJ��� ��˃��c%��T�j�xy^�$$$�w���x��3KB��v�w��IL\\	�!'�m��4~_���$��nvvvED-C n�:*)�Y�3�ރ���)�J>3�����������|�8a\P@���\[_�gh(�ikk����~EZ���8�F���MN^� ?���~>?jdEe�Nocxס���6��sŨ.���`�/
�h��@R��E�-"<z�\�G���`���Q��{��!o��M�*� D�
2Y���2�J掓�,)C�+�A�֪͍�k�jF���k�V̷ٟ�ش�-$,<�.�^���`�����lyU>C�1V�o�ї�����x���o�jI�(���42#��km��XY*{��O�	����5�����A�oo���������/2�֪ppq�SR��́30ڄbW�m�WmU�XcqN�C����Ev >s��n�;�DD췇I�Xz|xC?h7sg��e��X)�ɑ�y��8-wؑ}áw�h��ϭ��O��9ۯ�s�n�[���o]�"��ɢF��g؄	�ߏ���ݢ(�
��ѐ���!�R���B�yZ�emn��y�SHX-����r� �y-�^ �B]{N�+f�"��!z=�Dn�s��*P�U��s�*'�?1#,�(Po�W���Uw��/���H'�##�	#�iT_�nt�ЪZ��I�t?jR69�s�B�m�hp:8ը��6�.�}*�p
B��/��;�=����ᱲ������mtHd���鸻]���t�|Gà�� &bUNd'uq������t0W#__)Fr��	�A��{��S�-9�\ӱ��
l�p��FҸ���H|2a{_T���r��O�[� �I���S(�l�V�rJa|&k�+D-Vk�C�bЇ�H�k>YH���u���;����V�Y.W���4�%T^�����􌕏���Ȍ�x�Q+��l�?�G=�?���H�ֆ���ɿZ�Ч�����胈�|�ljbbR�^�8_i6x|l�Mw6��L�G�V��n@�'lK�ƃo����&C��#���!�֕�G���X�4+�ĜF����s.�S޻�
��<��&{lD���v�E63�t�V�������8y�Η�W:8K�A	�r�RR Š�o�@�k�N�����|;�T��w�)|�:ڀJ��<���R�D.�IƤ
� ` ��3�w��/`�<Q�K��G2�=|w� � ::�D���D�x���pZ]�Cœ����_:iI����`jh���[��{
�`�\ogff`>��a'��^"�6`�k�R�k�D�2��$m����`"GdNXJ
	�����>lᮻ[|������*���텛%q,�g�Kń.�T����'��.���g�a��I���	�����mW���onʀ^���U��nE��WQ{v��!�R�n��P`{���g��/�=���x6qk�nײ��O�C�y�F�\�k��4@t �p���IJ�O(kO���=������v�.��j�p����ID*�����y���}�����������t=z����0�6����b��- �s����y=9�XPPP�E��6�4[\Nށ��/5{%р^�
�ߪk�����y�f���M��V
�)b>���2�����7�	pp��Y̏/.=A 1ް3.U�a�S�.�kr5g;����i�p_tA��#abb���J���v� o��TG��/P�8����U����046�p��=��B�ssq�q�rq�'���[?������jQ��M:��ڲ����@%���f�k1W]���z#O�D���������ѱ�Or��*��Fǘ���9u�MMuC�!U����"HRQQUUH��/���^��x�ɵהH�I��0c���O��D�'"�WTp{p` ���2���
d��[r�.�=4ҧC��_2�3��}wPs��bdh(P��o}ټ#��u���!�/Py�fS�^������$􈁫��7x����\���\�k>�@Ǡol����~̼����z1�z�����c$C��1����"O��~ee妛�q�`�a���}V��3���щ9� ]9@9c{��@��L๹����Y�]=����O,.N5>j�<x�2x<�<8�"������F=Cl�䫺��t�a��:���37=����[�gp��"[��r	��**l����\�y��C�u�m�� |��l�J�py�3e,�'"�x����6f�Q����ncIe�/�F�y�$żϩv��������m�YVx��k�g����h�¥F:s��L�?��?g�GWA��,h8��+*蝴��_�e��[n�dܛW%�a��:c� `��b�k01���]��
ԛ�q����e2���%�L<?ꚽ�C��Pr]1�G�f���y\��	�Js~����"�n<.6mx�Հ�d|{���^#U2�L�p�k��		��m�� �[=��F�o�N

��Z�٠V�����o����Qf�pf6��^����N��f�;�D��R��a��c�M:��L\ЕH�✬,��+�z��|����4�{�)¾f7��K�Z��X��%$�ܹ�>���r�E��D���x�g�+�6����.��Un/����8�������nj�N�c��"�v�9����]8� Y�9����� ���+gq �}���Җ_��M�;,�3���߲^����j�S������Ϩ��������,�Ġ�!d,g��� '`�5��[X�2��A�̕͘n���r>d&S8	��<�ed�\���X-�l'�ArY������������:~<�����d����b��PȨ?:���^�d��';9)�MF��_��n@��pQ033O����4{�)�i�;����O��4�kp�gdT����(g?J�2>�`ah�:}���w��������	��f����J��"a�r�k/�s�r��7JG��nIt�b��帨q	T�k�y<-ݹ>	�Wfp�̝X "� tq��UQWǻ�G�V��|��ĐNn��^����Ra:F�$~�A����0H+3AH�������y"ټv�{�r�?f�m�qL��W�]a�7�;���j[��J��?d�Y��u���e9��bt�Y�����ٴ��P�K4,���$8f�.>�iuugoGg�P���e40z��z,�644)���-=�z�;FP�T��}KA�=l����ΐB26��, �־�����*u៫�3r�߽�uc�Blc[�Y9���*ք�����ǳZ�o�V8NT�P�@s��Ve�Sc�����t�[P�@����� 
J�}����XJXf�W#�珥˧i]>�A��rl���vF�Z	�PC�x
�dIn~��trb�9�^�g�mi�Z(��N��y�EO�he��^�����P%�2]��ܪ8T���J��ا����U�f���>	��� /���*��?�j֩��:�R%ߵ�����ʟ8�L�����ite���?��	i�]���s޷,,,<{}\��E�]��p]��Ъ���}���N.�i	�*��ڤ�.v�5�\1.	k�{mO����A~H^b��Ҷ�#<�hߝ�����_`���u�V�� ��m��t��!"2�9:)�r������4������p^�����Z,�:�~���k�?�����j�X]�@"8��n����S#�q� y�h����78�qtr:q�b��f]|V;<�U:��}k��]�`�$[�$p̄Yp�W��aw{���yo�]P�#�d�����St��� �%Z�ꊍ�R�,z�����wi����*��92� 4�V#�;c7'=$�Z�����Q���l����D�CSD���]��I�!,���_�����
i_�� a��/��]Y����RL��KV�18�fN�{��M���Ȼz�_�粪5PC�v�z�k�Ov6��ų�G�@�0��?�&��dg ��W+�*��y޹�#�R��$��&���Dv��/pp`�=o�]݊T+�J������[A<���ucS���XI������ ����j&'��x3��u@C!_ag�D������[KR���p��� ��j����`�TT
�*3�l���Z b*�nN>�=~�d�ܓ�Z��n�Vi�Ł�{���U�[ڃ����m,�׶�h�0|���аm{���`��p���xt����h(��פ�p�j�ݗ/_�	�p�z���V��RHNt�瓗�V�t0��- �@�7����E"�ǭ#�O"@��U�I���[��l�����b��Q�f�̱�N>I���	}ΐ�S��4+�R=�虷��3�ҥ�$�8.�����$�+�c�6 �����`�N���(Ȣ�:�����Mc
�,��F���ǙT�v��p���� ��km���Ӂb����+qM�q]�c��nT�a����l�"����|G����2̏s����(dՙ���o��D�R��(0!Tk=a�K4�ۋ��^��"a����g��zW;�4��ZxO�Z{/���\9r��x�L^�����x1�Ǽ�nd)��!O!���y�m��[Y�S�`tL��m㻐�����u�, �A� ��sl�-�v�ô�ﲞ��0��y�:=��������Qn����vTh#�z��]��z~R�K��F����a�zhF�s����w�ϰ�0�=暂� <�Q�J�" �����h�Nk��O�hJ��~`� ���x�z{�Ԓ��l�"�k2��:w����ץ���Xuu�B��ǩ��\���F�3�ds��9=�#>=n�z�0b���v��\�'(����)�@	�$�sG槷���0i���>,_Π�A/V��5b����UTT�����7��j���fl��8V=��{d"���~=�~=��=�/ �����j��lG�ұ��� ��	V��� ��C�{�B6��ؚ��x���o��c�K����)�{7xm/}7��Oiy�1�1�}u�_��� ������C�N5>�7�k�ط1G��	�h��ߩs�<�U���4��f,�F�&&w�&�-�W����:�[p�c�ZL���VRRJ�<������G�`gg_�+H�����M1�=p&(g`����˰r���3�t�ՠf��@/������W�$��D�i����ka|���@�%�1�h$�b)��A��Ƕg�j]���%Xа9] _��+-��h�?3�3�>�CgS"�Ȏ�ꕌq�ܶ�A�ݜ����\����K�����whW�np��e�SRH�rd�L��ػzz��J<�F�w;K�����P>���ཱིآ�Z�mo��%C��,�d��-��&+�L_�ߌV���k�N������e�CF�q�;>g6�a�3�>s@����k���e]���Z7ɦ+�RVa���q����Gˡd�!ϡ흝�-5�J/.����.��:?��y[�{�6������b;�OF�$��S�@�e{ܩ "���lP��6�r���_��,/�K�h����JK��b����L_�g�/�_v�L�.���_���}{���G6�竢�X�y{B�|އs�7o��P>��n٘�)�"��a�k(�"����^5K	۲*���ox��P���*l˒ޛ��jF���j�o]�!Ļ���u��*//o�U2�fH��ۯ�%/��S�3F���~ã�>�e��^�����+�H0M�Y����	\��mrrrgOaQ��s�.$��A����踸�;@���,��A{�b-kv���
SW5�@�������>��qz'ק;��&#���~��=lO����u}j��I�J����4�M6\蠄�A\���[Z��vC������\���=�)Z��rUX�xAdt�S�l�/�ߜI�"ء.[�w�'��?j�/+�Ӿ|�2�L3;�/ښ�f m���ַG��e�b'���a��sZr	��P��z9���;��U��rTG\��݌��ִLI�x�p�!gl���۷o?/�?�����gJ�b��@�^p����-�!!���F�@+H%�E	P+Ꞙ�0�*�mmK���
��l�]�كcP�a�ѻ�����[ �]���5Qek{�%�ޖ+y��@z\����d�6��]�-�Y���ƺ$%T�N2C��I��]f�����b�1'���)9��[b�b+���"k];S�ό���{v�����c/@��c�r����ʟxCL���7��.R:��J�Sp"��JX����~��3I���x6?�x���5�`Vi�����^݇�����pܻ5' �}������*�0Y.���r_����Z����Ϫ*����d�zֳ����L������OH��X���&�����z9���8Is�-����6�A��:��zƋER4�$~|q�+fl�_vz��c�x��oؾ(�ʜ��,f�TI)��uv�(X��5a/�XY�*�#���AUpe�%x6ߺi����y�tc��x�,���FVc����vp����MW�7�Ȃ9�l>�֬o�j�r1X��~`�܌�KDۜo�x�E1(��I�Ѧ$��Wي��uU�ig�$��HF�t#�ii�1F�vuC��q��@���n]��s�;d�J"ǵ��H�=��i��|\�M�r{(�~��V��{��n�8�)�$����~�#�Nc
�W�6�#z/�� M�t�Z�wvu� 3��b{�������c纄�2C@ٿh�����j��=l�>&�m!,��a,[j���h��{L%%%1")ek�ĳ�l��-,����|�ozd��o�*��3��F����V7̮g,�H��U�L6��_��Yb�ʀs��ظ8�ghR�ɭp�tF��5�5�!O�H��m�v �_�~�-aMbn.��"$K�X%E��#��h�\G�FSͲ��j]4�\<�0�E^������I%#�wYMM�|��ʓn&�2a$�����ɉ�r\��9EI38��p��)@�r�t�/5]|��G
�K4�޽{������A;MB;2������lRT ``�P�[B�euk+f�# ��36��?��g}����gʀ�p�m4�4�}?^xh�;u?����m��N�d�����O�us/8���X�O���W8�#��6;}E�Yڇ�����c��~�;�b+��&�ɚ��;��z��<�Po���j�9a�G��k�[�<�7[���t�ޔ>�A#��}OQ���ܤ/z��qWtgg�ǝ����Uϰ����k�+bd�:7���O��n?�/�%a��68;;2'�O�GeE���?�
�Z�w!8�1N1�[^���f���'�=��H��l���R������|�=��[	>�=t�ڱ�M����u���p�%��		����˿'��H�t2���!�����%.�f��eC�褂�W۶8{l}?ۄr<��̛y>;U�X�����;�.6%q9����x��γ5���.�Q��_�D.f��J����ҶE�⅛";�#d�3>%�h��@ճ�ͻ*.�} w�[<A�
�F���ձ\3�|D�VxyZ�b����?A�B��db��o�����;�"�D��g��i�7d�C���:�/�ې�>/�l/Ǉ�%;⍨�-�z'��1�w���Ot� �nB�>�s5�m�Z��.\zkF����7vVǰ����.-����K�N{�DI7�zi��>o^�v"�ݜ�|���,������а��V�#��u1�y{��	��p�?�i<�L��+_��ꦎ���Uw�ü�+�݇���A�G_��<<Ih/(@|��R��w�.�pƊj��v=E�B������6r	1 �6�{om��d;q�s�����u�VĲ�GO�U�O�v���B���{�g�C�ETy��#�ǄO�}&|44A@q-�F��al/h� ��G
#���78	ͪU+�sޏ��yxd���
_l�A�ѷz����	��442�d:Jv�?�q�&h=����D�����+�i����v�Y��� �A}n�Y���;�����w>Zdq��k8j��?Sqָ������"�W�|��I���������	��.���366��[�y�/��+Wk[а�����Y(4)b��4�>-�h85��[��m��g�X
����|	DM{��)����Y�rn�w��E흯c�ߚ�3�t3��J�p77��9� ��ܷ�D���ybIT�z�/|�\۔�J�~ߟ��i��VX�8�˙//�m�˿+~�rSRY]��+�.�y�͎8ΧO�5�j������U�����"#1��"&�	�׆Ǉ�����c ��� 4�}���R|kb
H�~	M.��n)X�5�d��x=؇�[�pƴT����o�/4����~�|د2�/�u�و�����.�~���|F�k[�qJ[őϑf雽���u�Ҕ�������?��2���ic�%"]҂t�� �%]�t�����!���ݍ��t�tw�{~���|���gw��ٝ�A'`I��a�
�A Hw�	�x�A����,ø�
2C1�DG����=��^_Ȳb�
����h@R\����ЎJ����ZF�����d�ׅjT]n��q��i�It���s�.�t����Ov�	�h�Bi>e���R�&��cg���.������2��%ե���Y�|�h�3��@���LN�c�������b�({���{X�$��@3�;�j��D���5�&I��;�C][R�Bv�H$H.OY�Ͳ�^p@�Wk;�-����)�!�ߩ03 H&
诹#�����޾|�x��#����1r)9��1�G�,������]��+7��s�բ^!67�`,�iD������ϟ/$v'��ﱝ�k�8�j��o�?����f���?O��@U"	�!���)3X�%��P��ɰr�/����y�ɧT�L�#4�~
d7t��r�A��ӳ���L�����F�dV���-I>���Φ�fF����eS6&:f"��9%2���E	u�Mz�d0	w�ˑQ�a/c�D�Kc�J�Y��&�q����]i��s�P3K��ѡΘ{�L�����0 %�<nk2Ŀ|��t��gO������r�rj:O��*F��|�%��$5��� ��<���2�u�����|�+**��l��2>x����#ߐ������`�<ŭE<�=-��`���+}��rTˠh�_V�S��xd�!
RIRneFn3&r0�-�;�w�nt��49c��rx(�d]�N�iij�؛k.5x��=�yxo)U'YP>}����S�W\�q�B^^^5H�$��t�Y��RY�U�l]������}g�J7��Қ`�c���5\�" 7���Yv7�r��a�ڶ��|��HM�D~_�!_�����V�����q�5�����I�3�[��E�����∰�WW˓�(((���*� ,��AB�<Ua�m�Y��`����=6֨YE�S���OX�{����x���O��X;H�"�H��&KVQtk�}'%#C�*�:��	����ܝ66X�:�yl^YT8J.(G��r2�y�8��lg����՘��Nm��C�M����^�� ���ӽ��{��u`k�q�B�����/�N�tR4{�؜⤳�F���<��e��c3z�-��2V<�cl�L�:�Y�h�#��3�1�3�����A|z�7�z�5���.�}4LnmkC$s��u�a�-��lw&�0��⍬����%.�I&��[���LTT�����;;��~�^�jhg�T�@��)B���x��6�`�=&?��d(l������y� �`��C\��L{��f��A�n}�ܓ�{O���eee����H�nϩ�Z�,Z��!ե$F�l�N�	0TJ1�1VYg311D����t,�����a#:"B�Āp�hb�	�+�}�D֍�������Sod��#������7g3	pT?9Qn0i���g���23����]U��t���u7���������lQ��PQ�/Ԩ`��,��p�ҋX aEDD2e���k�A�j��a(U8q����η��/!FvҲIK��!��X��&�cb�_�]�u���w�}:����!O]���1�@ �s�+�f1[���{w�:��뙾Ğ����-tob��;߉���Vk����9���C�u6�����o�H��[ȳ��]�s�pZ�	��ׯ|�L�Njt�3�p����&�臵�ϻ~}q���=C���OnL�`l����'+h}@�!��!:  �!DS���ܦc����B�U��3L`���Nn�q`�G�Y'�m��$�
}:D�e�А,M�{��n\TTT ��E�<��>�kN�	\��w�]��Q���+�V@�i�}44LS-ց�U��@�yy9C(j���f~�K�eN;kӵ���%EĘX��WG�zW�t�1�W�WS��~v�#���'�����v�z��]�YU�v�4���ܻ��|^��=��] y��Q����$�t�v��nk��KNbSk>��J�On3��LZ��C��x744P�cQg�6�ϼ%�>\��;BGG�.Y�
��5w��$�ԝ��f֭��e�{�����=Z�}�)omB��G{_�x����ðm�;[�Os�(P������\@,P;���µk�T��o�R�X{/I����y'

B��Ƌ��\��߼y��}�ܵ1QL�����*,�Tؠ�>��f��Zg���Y���L:��QP���(�c����ϬM�J�V�%%��[��,�i�Rj%_i��3��W/�
l��t��>��U�����>�wi��Q_Q�l�i>�Ҕ�M����H��[Iz�����^#���w��?<�c��"�Q�'U}^("��D�����TP������4H��t�f�Q������<�Lsw�M���4��>`�V��釵�^�ws�3�e����������2U��c�E6v��?a 6X5�\�po¶�C<�xJI��*�`����+��w;#������e1�ZS��3w�wf���S��K�����B�/�({���,[�vx��MX�R�Į�{NO���;���Ԝ��1E�>�-�C߰_�l�Gwo�ԕ]�`V9z'a6S����o!�j�� �<�USװ`�$��0.�%�)�x��:_���r��4�6q����C�?c�-7RV�FI���y�(�/��"�O��^�2��қ��13�ƛS���Yх폀&V�(j�ذ�m��wLِ����n�����������Cۧ�M�س$�hfM?�O�g�


jeF���|E<�G�K�3���F��lA'4)I�"0�8)���s ��C�'ۿq��W����n���̯�'(H6[�(Ze5����Ɔ��Z\d��̌	ޭ�-�у���<Nۄ@��G�ɩ�C������vZ����K�E�<�SA��^ʙt���Q����m��j/�T�1��`B��NK(	VAjk�F�Ftx\��X��]^UD�g���+N����8��L��ή�6���t�������L����@|FD��F�z�&�\�&���
y%���]0v`��ϵ��gR^(�V#�?�ƽ�|}��տ�"[����_�@��EVm|�	">�ѷ�-1		���̺jZ.ss�꺺e�sD$8�Fs�v�C(�BVV>*,Cb�ϟ?&��FuA�*��q4@����L��й���C�E��aa�H�]/II�������℮���$����P��j�yHH��q�˛��+�R�<�)Q(�]�� +#c�ټ� o�꙼��D/&B�G�s�����������1�V���3==���Y��D[E�/���
*�'��`��*E1^�������d"i[c!Y32�۷.Б��'��<I��t��cx줰�~}�B�D��C�B�:W돊v*�q��_����m�aN-eٲIf��ŀV+�<�D&�i�Ħ:�3V���W �,T.��TV�͓it�zyK��湕��Xb�R��|��2� ? ιp2�[�b���ҹ���r�6�A�3�q^D�0�|v����:/-WN7��q�" �ɳ�����9*s�i�R-<�R>0d'����wy����RLDDԳt����֞Q��p�V !#�osm�6��N_�jiy�w�x�f6��wMh_ C@��Q2��4����{�R�]Oe�	����l-^(�ў2 .ϟ�E��D��d�
;�4�⊴�Ի�; �k���5Yc�����٩bN����愈FG[�����n��Zw{�Tt�hw�!𘅍��ޠG"(."0Ԣ�:�T�.����5������/]T ��y��)�f��`
VxM�366%ü:��> *�vt >@f7-�)�����f��Ă�j���9�}����}"L-�+�$`w`�8w�?ڳw��P�x&GRGWZ���/U����V}��2���`8dd��*�����qccc���<nNT+�*4��өY��
瘞�q�"�����g>�pp<33�[6`����dj-Ү8��<g��lw6߮���Jtn�3::�BU頲ghhh�+����Tz�I�ɭs���!g��6{>`�_�>ޝ%����h�푫�y)HNCC��-�B�l`n(�t��qujI*䮵^-�t<RF�k5/SS��i�L���Ԃj�D����$ku��������;�7�V�>PxJ�]��5�<����#�������ğ��x���^����[��A�:y\���iU\����>���59F?����Q�V�u!���l��J�qqu�H䅪000w���(+����\;����_BC����M��<��G�a��P
���g(���z���IJI�GE��R��s����|068��}��#͢�ݾ�0����<w�ր�����k�n�n��ӯ��0'-G䲾$�����f7��,u����wd���{4�#}��,m�Ćwb��&���]\��߷�;� z|@��!�Z&�V�'���+����L�do�RTE�����;�>n�H*�4o0�
9���[�޶����#,�I�u���9Ǻ���ώ���6�+�Hy��S��ee#H�e�z_S	Q\����7��,	�Nı�mgE�яM���GW�NՇk㔹�pO((�'��7 ��݃E�rO�:>�^�	�逹 � ��6)��{��*�p���]�$ϟ��s��x�����@�&.k�U~V��)�L�p�)3�U>k��P0뼱t�@o���4��MC����jo���S4�BMm-�H�,�@����p��{����V��d?�{�.��������w�����JeLR	�PO_���ݤ�{�H(�j�+ev����`W�c��z���*Z@��8h^]���m*�4�����}��|�e��{=q7)��R7�8h��S���n�B{n/G@��X���pŦ�W��z��B�r�$KL�fPM-��H7���\}
k�X�,�_Ch[𿑳���<��m�LɲV2��e��=�;l.��M�
v������۫,rW�D��u"F**�u�WT쮖�ʣ9^pU+K��dA�ar���	�����W?�"�L�/*�3r��iX�+�/�*��e��B���]Jd������<f�JL�����%H_}".�x���
흰�ڧ��r�O��0��=�필����`&L$+�d{�&)��+���?�����d���s{�N�F������H;X��3BD"s��}5���͞���Œ��UA J;��d4|�9�_�P�h���[�lq�J]�������ۺZ��m尾�����y�=Bo�����vm�����F���h�
�� HDV6d���e��	��Y��q��ۑ��f��X�2�y�U�C�wW\2�]���{Q������/ӭ��$
��n۞حV`���j��}|]�b�;�ͤⵆ�mS,2�t��!ڹA-*��S�-	4�0��R226��OS娀pr��+�o t�J����a���_��|�ٵ����}���b�Y��?914�����1iFg�֦�����_��II��t��:r�#�6ŢA�r>a��>	HJJ:� sz%�{��F8ݴt���0&�}Qe5҂H��"V��e��I��`��m���-TZwc�ƾ��V%���eM��˿�L�)߯��u��{��P��XR/�Ϭ�z>0[^���^�|f�ot��@����o�oi�b��~��)����&��{��)"�E'�=�D�g'*�&���c��x�+�@
�����rٛ�����}��EM���QM��O6�Ka6h��R�Y)j�v�[�Ė����Q����W�HL��l���xgzb��1�=���؈0�ϕ�Co���N&E59ٟ%i�{��3}�tm�����q^��5��?BH~��	!�m��[��UU]7_j��#�u֟�K|z4
�ÿ����6F�p�..͘
5	c�m4��R4y]���bcE�	)	�Z_�gLǟ��Z�%lfưwR�c��
���D<I[���\�� �������z�����
�ۯ�+z3�b�i"��꺰�q��z�_�d(,N[7�M=��v�.t'<�,xO�^>������;N��l����c�6�c^�Υ 0�Cg�|\�$�sK,j�؉�̵��6-k�˭fc>�����mS�E��ϓl2�v^�_7�����"`�Vz9���-�0���L�ۑ�����-��R�(����վ�H��/��(7Uz��OEI)��퍂�V�K��$��9�ß_�g3?~�__���u0�ۊ�yx&HC<J}cG�����ֻ��`�j�17����Y���ϟ��s:!��{�)x|2�d�;X Yd,T#]�&��M;�|{��gU��i+pl�H�.L�?؀ٝ����(R/�A,P+����5Y+��ei���93�_����������9�����l�,��rgF&�Z#�o�A�oC����އ	������y�#E�:��%\�AХ���,�'h�M�rI|Y��,1i.J�l��d��������Z`Pi��� !+۹��1�W߃��Ѿ���� 9X��L���'T薐��Mm��i����X%f�2'�*��48�89�ZvioK�pC���b������ѡ�e���V�� //6ū�r�J�4���XTY��6�fRq�!��	�cG� =;q��"4=��?r^>5�-��W\��d�5�q���'����N4��-���PC�H.ۥ7���G�y*�l����S�K�fR���0�8hr܊��w5���YXY9���v���W1O���~a��I��z�����ã��ؒҝ�.G��F/�
��U�|���x�)��x��QT�8\!$��&O����w�1iP���a�]��+�独6N�E$�<�r��}d���\A҃�[��%%�W���{��@Vq��TtW-@+�zSq��S:v�f6�\A_�p�!�
�.22��F7���oڻHZ�V��(#�7%�U���|JC��M.�ZD���L�RV��zb���g���4
�s�R�y�M��Zg��Qm)��Y#몖��q�>PE8?,�����C}��'���i[M�Յ�8�a�9D=o�l��!3����@�2������|t��o7	���vG���K"��=1��	�<�/P�V�[o��;!���\���S�B������R@Z	�ܷ�����..��(	�_hTZ����������૜dgED<֪�C��>@��hI�п�b�`�����`ء䂿x�	�>�W�ef��5���M�$�%z����������H��y�!p`a��L4��I�m��N��=;�f���&y�i5\I�6����3��N��Y�0%�G��454(�Gl�b?j�;�躝��=����C��d9D�J���}��3A��;��eĘ�.72���C��
��P�l��x�5�SS�@�8�'��Rv���O(>�ߛ������z/�Jӛ:���㼖���G~��NhfO�� ��%u�mp}?�n+�E8����D^�*����|�x��;4Ml[.�}�
���'΅ ���\��{I�;\�7�[���������`��"{=z�7D�B6rE�<_-�Yi��Hp���������,T��ݽ��Al�l� � ��/��B�㙘����R}BJ�FF�"���+W����bbY�?�Cw� �t�V����ĳ����S�U�G��pB�Wh�E�r���[�y�[[L��?�Y�9�:��ؕzgYE�W`�hT�h�T�7�)����w:kBx@d�N ��+8s�?�+D2~�'�ni�� ��ꬠViA��E�BBB�c���Ũt�|�a_t��c��e5I|�SzSޯ�D�6�|-/��J�Lx�&O�7�����
���j��T�@��Y�4��s��V'���HY��B��t;�s6S3GC��XN7���I�9�|ܼ�ጷ@�N�|���9+++�� �����lJ��J6}���4Q��,\�J��0I������a������s�B�ߜQ���.UX��s��k�_�����1m����0K�m��e���V칳����kk���'ᶲ	٪C��<a��f5U�)D.�rW���=���_6��s,?�$�riy9�Xa"��D��3T*�����PƠ��R������b"�=��DqWk�������9�Xр��*��r�\������*�f��c���3��"׍|f�:��3OO���VR=K�%�Xf��^~����|6`kͪ�������]]�(I\�a���v��M���W/��~�G��e/s���.���a�.�Y�W��T�{s�;%�-:YiI�-��$$$�����Q\��/�[�.0g���d�^��]Q���)i�3�UHI��&)tB�WQ����АFD%q�B3�V���O#N���z>p�-�Rӻ�5"C������s���Ǧ��x�;�]+�?k7��֯�kh?Yߝ�C��� ������{ծ�|�! ��Q��������7n
P&�����NVF������"F����+	����&y�H���Bӧn���dA1�/�)�����)�����Q�ΨJ4~I�1�K
R�|�3����C���Q)	����ӑ�[^��+����x�`����$ҁAg��ƃ䐴�k8#�*7}@�W�[2+��fAG^�.�(~�ob���r{v]��@������!Qy�x*��c͂�h�ƫW�������k�^�0����͖��$��|��Sﴷ)Y���|D ��W�=3���61��b�|ă�)�������������X&��ߐڞxquu��_��۩�����G@�>ᑚ�_�|ʣp�h*�5�� �i<V�d`awr����TաXpg��\�anײ�w�+�}s�.�*���`V�'"2����.Rի<��۽ηm~��X,��� H��.�C�"�]h������_�e��n�)������:T���9��������;GTm&���~D>��<�{�q�">�`6��A�V�x����7��z�XY��2���v5���0������\�ڄ1������yJK��#��
��p�6��_�l�F�+�h����9�d@�cV	{����eex��Q����=OY[3:��(o�� �X`Y��w��d�bCf����x���^4������t�/�k5�l�.>��ؔ���܈����b�����J�,ٯCMe� ������x��9�V�1ld�'e���]V��w
x�N�`:S��{�b���q��_s��{���!nn@�_��������F��_�\��ZnAAЄ Ц�..D�	�y2	\�rR^ 暧�/f����F��71���T<���^j����nϴ�gz4�X���fk�� �&*Q��̈́��MC^���V�xQ�$�_�us�����G5C�t��6�V�7�k�B F?[������t�PRy"���}�s=��xr]�~9�7����_N.�:�mڵ���1���$'$$���./���^ ��K�N�mdΊ�1�Qh����8��A �xx a4���u�X�������� y�2Md��������6ڟ��w�9 ��4թ��7L�q�����NK�JўWd�W]ؔ13Q��l<\�� �5�UC˟�'Yý������Uz��5S|a����26�~����Qʝ^��{����׀Q<��-��sGxI+U͆�{��z�ؒ��>Sy�d�wYNK�w��J_��6�ZB���t�EQ��J�����r-CK˞7tt�o�����˗sBr���Y|�69d��3w�xxx�����@@�G��UbP��!ʰ�9_���Ne���G��U��O���A�	�}* @
@2��nNP@�x��X>�H�#2Y����J~i�$��-PWx/﬷����u�z�j�T�,���q@���,�a��Ɩ>m:��ډ@�ۚ9���dy�3q2�*���A��ʖa��5ݽ���^�z���z	w��y䔭#�&��?��t3V)-*5�߬2�=|R!Y�O$�7���
_#y�?����kT֦����`Ȥ��W^���l��~w7bTCg�_��^��7��(m{�����\ư�e#9�\������U����G�܊����H����bN�ol��!�y5M��6����3?�z���V/4�$�3�0Lc�H4�ŏ099���!��긩�=U�-:Z��1�Ň����)���b��p�mdT#��ǡ�ȵj�?���x����n�8cf�)�(�}���I�h���^u
W�(�*��X�F��D��3�ˢ5_�<�ra=�=����fn^I7|����b�pڋm�����Й՜�& ���n�.Z�x�$>�o�8�,,Xqqq�9���qUgk����ţ����UW!���q���T^ذ��j��(U�*UZ���y�K������O��븖�qkW?-�����7��K�կAg�S�I�~-��1{�Q"��.�֥���e���������c�V�bXp��(�5�TlG��-��8䗩>����k�ʈ}��t]
�urI�P�\IXߎz�2��s��Q���܈����f����'�&�T��ռ���:�|��@���ܞhni������RR� \B��o�W�ש��\\\�珁�+)-���~p��}�D#�CEEE�WVV$�����\x�v��
�i�G��WسO&$Ce�+�ikZ��o^��ON�*p��b�h�Di_��jݹ�:�=�|��˦���k������h�0cUTQ��pW��KH Y�266�.g��6:*�W���**j��	x�6�\��ׯ_#${ܺ�﷢�����A��?\y�ω^SS���o���^�z�8P��e�mv{�s����a���x3�_Z�������N��q��Wv��Lz��� �q,�B��a~qck8�[��筭�P����@��H00`�_�E���F):T������m�	�i�������!!	��qEɑ{���pĉ� �JA�7z��Iٿ�*��}7H��y~4KӖc�}ɨ݌�L/�4�>�<]}��O���*<��RE���Ϝ4����i��`UhWY:\���6z200 F��׻3�d�5	|�B�let���O-�7�HŰt s�x�����&��>[�(�M�8vD�Q�w�_���5
Ϊ���K��_�hi�Ӏ���8��� #��ĦX��z""l6��h�	؇!������@fU��IRDH��������ԔP���7�v/����^�W"�VWi�/����o���̘tI�=ui׽a%�r�yN�"UD�&�"����8�_Č	��Ĥ����jL�Q�d���>�-�+�4W�%�>�������3��>��MY�G����T�E��*��/��&a VZ?�;0p�~����������ɕ���+.իW�`�F���[��u�	HJI�2/$X7z,�����m���\*/=:�{����,�oGT	f����-�nNMM>����ްİ�j�j��/4�g�ŐəKcԞy��v�e��)��j_�:V��c�M���ݮwwKhA�m5���l�/�gj���v`�3���yZ�������h��s@�����j���<�0CJZ�]����dk�d���?K�d�Z�(j�U�6s(�r�q��9_��t�]��0�������oX`�/g{:��L��b	45󑘖m�m"z>���.6����*�ȃ��u�լY����'����c=#"?��]���z���DZq1�T�%�������`�`z�{\ �_���������1��WR����ߡ��YEw_�r�U����L���St�x�"T~ˎjLM�a�$(g��T�8\��L�%�V�E$r�x1���`UJ�<�"�wr�髣 ��JGQы^){��U3cq=�ۼɩ)*�'iii�
��z峿1I���S<B�]	��*/C_�|��)��w~�h��5�y�]�h$���U���!>��G`aG�U�8��8����͉�NQ�-��F@@09=���X,�����1��]��{M]`~�`�Hٽ���g�񍍍^�K��߁{�� ���@9}�H���*�5^(�=2=MB�q͆E�J+'`�x ����u����z-�$6?�K�aL�-BO��.,�Ji��߼3�n@�ޚ����|�l6+;-~>W�:��rC�ޡ�}�x�Hj��2�NX�$ٚ�������<p)����p�7�����������D�l��z��e0[ۖ�4�R�Y�����(U�,�2��l��R���P6
�b�߆�I�2?z�̛����쨚}��o����ɍ�a|�CSt����h��ᑑmW*A�ͯ��
;K��ؿE�o��׶�45Di����L���w��@����l�����䄈���.����X~���֙���,��]ޞ�������-�蔍��,���Q())M�+�EDD6g�r��E�v՟.~���5d�ԋY떤�Nq8|K��z,�ٷ��o̾X^R����m�*���33��)~��]��~�C��R�uk�8S`��l($ߒ$�6<W��x��?�y�dO���A�� odl�Õ�))��B�	�_AH�R�BGG����_+(����4�gam��${��Y��.��<gЇ��D'�@�4�T��}��6�NMHY�U ��<OD��$֝-�z�,�l��tml����gZ��z2���z�����0�J[j��::��Ʉ.��@�ޙ�\�Y>�q�����d�������
��xxP��XA8�����o��.oU���lK�0�/�8�ܸ��YK�T��	;h��|-̀z�>��x�{�r�j���lF|�&ܾ0��!��Xg4۾LvU�⟐���状{9�-����v�b�?;�c�8��k?]��ayi�9���:	kj"%#.I���V�M~�<�d�@����ab�ߏ��������
RDP�V��_ ��~���x���p����KLi�h�oJj�hyjadj���J�$�7����l/�M!Fyw{ִ���ͬI ����WF���2^@@���Nȏ�jjj����84,f����1�-���|���Uf����2粿p��s��.
~�u��>(ГD7���?��==���E��k�_�ݍ����}��\�~>>�:��U$~h�HC�(f2���P'���z�.�=d�>e:�+��<e��F�[��(9ag�����<��6?��#{��� ��3ԥ���Z<C�Q^<edDgaa�"���MA� |2��D^jG�{ߚ�����o B:������"�I��aFn�F��$��gC��k/mx{�a��!FK�f��t'5��}�^GBB�J>�v<����5.��Y轓��B��wec�i�?�ND3-g��do�bcb�6�XY�(*)uHH���EƧ���>l��ѱK�}H����$�fb� �goP*�Y@��s��o5��kj�����֢=?D�����YG`&��+���Gr]l��хI�O�ٔxj��)��iڎ{*.y�b���5�΃*ks7ҢJ��s��|o�hhMgr�o��v��:��{H	m���}�E�~ T:7a�[�� �a�����dh�ޘ�h-T�7��.w~  �102vH�ma��*��t{��P���^��H��^tK�~6�ةg`y�t����s�f��]�Ņ�xz.5������N(ڮ_�.�$X��&�읩�eR9iɷ&6�l����_��� 4k�{=�\Y1�bي��eنl��d�c�Ӏw�aS� ��:��}Ux�RlNXX�s�&::�u�Tȝt��h@��C�k[ňګE�V3՞��`����dAq	�ҵ�y`T^CCc�|�y�e����_.��zt؅˛�+'�M͆�gl��Hр��%�|)��c��I֝�R a
$��cKJ�W���h� d:ly�it�n����L�68X�ܙ�t�����7�I����w��}EWDD��D��volB�$���o.Oy��DلEn+����@eC�X�Z2��3;RB��Wܼ S��<4h���H/Ξl���̵\�ʜ�3��<Y�k��V�����yq�8�	ʛ������&�KK��7 ���� �0u�d��;W��?9u(4��~�����6h[]��CԔ�J8�a�W�_=!�as��^�f��ع��o�\��rZ��;�l٤ _t���z�M��4���K(/����0$�:����/�Rl�~}7S|¢}��Q�z�	��l"O�H�Vt�H�1DU9�F(Β��x�7��8�<���|k�u3ȉh5�ZZL���Z,]P3@��n�~�U8�ݜ����
��dŤ*o�a�hi����@V;X2�.0�m����2��&q0R�\ʚ`J~�}����S�F+�8dZ��ع��-2�N����(�}�J���a&�阹����P�.�glN��*�u��?�\�6��4O�:�;{��-�yߜ$^{��6!<4���M���������-�"4א�`���t�c������P!�����7�nl��t�8�`��I'"QZl>Q�`6k�z�`��E�C'��4<������W4����U�w�6���˺��l�����������6��䄱�6��N�:��.zT5�]r;;q��C&���J �Xb��g̫w�Grl���&߰�=U����%8�~B׃R�k���I���KAh}��^O���}�����Ϩ����#b�����l�#��R�`���`"^�5i/#��"��p��#@g�g�����%�я��m<ð�Ow��FF�֝��:k�Q�kxU���yD��wF^��^��=g`�kt�ω}|��I�x1��q}���`rG��C�b��@�[lpZ��T`Wn�`��h��P� �o/�qpq�����ufsa�����ش\�c�TZ���7�KwzbL+ѫ�i�T��o^x�����S?�8�S�P!5Z!�7)I��nܬAII��zmkJ��h�F���a�&�u��V�Kk�xi�9/cb��6����w�;f&<XVZ���ޓ���S���n�<�/�4q}E<E��(�����j�=_�5ϏG�p��C��U�O���m�V.-�C��>�u���CUS{n�=φ-�,cLc�3�qf�*�pe����@XBe�}�J~^�E�!**jwo���A������Z:�_al��a��U箟0��n�د?L�Ӎ�o�'�<�I�F�Ix�<��f��=//���o�����ζ��L��~�+��z��m��\�-�履�v�����ժ�Ƞp��lp���9++����&�۷o�7���B:ڿ�B�{~y)����1gT�$y�P����Ϝ�әp=)� <1��3�'��{�����Z�p,o�b��%z����̞[�>�8J*��h�+t��c��3�ouȄ�3D�� !+��t�Պ���xW��jԜ�Ok�\l 鴹�5�и�K�����:���@t>��-0+�]@X�3?>^����aA}�@rȇ6?T�d ｼ�mo.u�T5|����x�B8��d�֛?��9��'�?C};���""
�������� $Yz�~�d5[k(���%��5�����#������C���-�����^�;	��_YR�b�5���n�>D��ٹ�0.�MaccC��(8���C�9*��I�J����'X��
N�*�WK+�'�A�؛�b]�SZ-��_F=���50����e^��a������D��.��n�/��RHM��AX�KF��kܵ?|<_����u��x���6����h����-k��`��P�9S���ĉ�ď2�b�\
=�,x	a6�����A�R,\}�%�R�_7�H�E�6r���51)ɼ��j�dR�!<H���d�3��V,0�um����V��p8��q���o�4����\l�1+�������Ã������~ee%��3����/�x�6��"o����^ƩJ��7�(:�u���`Q���������{�`�AT)rZ�����eی��z��^%�j���Mul��g����Cu�G�7��"Y����[#i|���D������YL�HB�!�o-����Q��n�����1�8b�Mq�-7V{����q"�7��,-�oo��t�}��z�i4�(�����(�~��n�
�ᗚW��CW���;/\Z����^R?��A�n̮]H(��FMMlW�О�����:��\����u�fX��i���?�}FFƹ#n�I=�z�
�ߏ���s�B|5
��+P�Iu5��<Y�ȸ��d�9J?��V7G0��� ����� <a�#�5p@=@���Q�,����L2�*� �pa|�?~(ʛ�����گ� /��i�S�TU/2"�}�G�iJ��Wl�q�U��썄��6���#.��7�.U��@'0��m�B�P���XG�,�2n�"��������C�Y��Q��"�TWW�ʥ����n��(�&���_�����w@��s���D�~��Ѻ(��j%�?�N�V3̀a\0ijj~:���h��-�⑯R(4�wy�ϫ}1�2�}	h͖I�N�<�&�̤]���O�C�����6���C����U������@"�'q�Qp���|Lg&v�3��o�BMǇ�����k��O@��O(�)�6i���~�-���ϓ�C ��ۓ��]��8e���7L}��b�iД!�7������L'~��������N窝~W��g=��io��b����O��&�����b'''�z���d�K�.����T<�d8�����k����P6ZZ�ъ����]�K���M�B2yIɀ�3�Yuyn�+<<�=y��*���rr�2#L��`U
� �+���>��������kdd�0�,�����&��Ă�/����7F�0լ_���^�g��|�̮�6���Й�b�컟�v��I����xm�uHC�6UiI�6�2��e3p�����41ĝx��)M��T��P��o�.��G�W[��;�A�������hIۅ���`�J��'77�
�H�æ+�����@4I����h��>�:���>�͘�ܟ��UW&p[s�^:���w�=~�X��3�	�[��~iee�(���xP�ܬ��*\:�`�x��.�i�z+��j�&8����L�51Z���i�E��YEu����{$�%//�8~���0����G�aA��h�2L����{��^���m�?�?��(��kF�KiP@@B�K���nPR�S����F��;�A:�����~�o�wp��:gﵮر֥��]������wb?.f���Љ�Ud��
�|���/��Y�z���Hǻ�Z^��%	�J�%�3��j����Ka.�{���M���s�I���إ�;�����T�����F2Cl+Ҽ����g��u����9t���|���z��'�i��ǻ#*����c����Y�lD�Xn��u����5^Ub���m��"��yz�)��P#<6��N��'[Z �*�:_m���]?�'�u\��P{�d?�4v7�H�Fz��ڿJjB�Ix�]��0�>9�/?k�{\��*-V\]t:����ZkNU+�I�B
�q�2[��Ѵ��Р���*���Z���K�Z�ϳB��l+7_8���p�G��:�^�<�M�?+��K�2����|Q�䋶wCؖ~�:L�ө���L��|/uۯ�1\�U�%�Y>p:p�
P�F�v�RSS�����)�������G�ih����cz54)v%��� g#�^#Pw�5�/kD�Ѣ8�u_�ng!Έa&��,���h���F6(4dXo,�ؓ�eH���:!!A/[����B�]Q��-���?��at~��>;��XHZl�*Nb6��ňR�q��p���o��঵d*w3���ղi����&�I~V�gϞA�K�肋��62:����~�',�zfa���ϯwtt�i���C|V�F'.!Qĝ{/!!Q�ب�D�� s����5�����.� D�.aY��j�7�:܍�?���s}R���n^�s��vB� �"�A��2v�zzo�5��\�GSyƛ�lR�i��EBϸt��@w�\��aSL�zN�m�؎-c7��`�-���ʴy�M&���!얓�X�&$$<��` ʴ\E]}�~;r�E�����ցx���W�Ry=��׳�ox�_����C bRD((�DE��Й!����cg1�ϟ?��&���BP�=��5�^e􌄄�O�9ds�SZ@@ ��R�2���M��E�la��}���Mo��---���^III����D���KRvV�a�&�pǣyָ�m`lLvf�ag��$7����Ȟn!:(�����I~��6�金�j����P�d�B�_㫮��`Z�� PTBBV����Eo[y��ɍ[C��Cr����o���(�~N�g��e��a�z���[gyC���>�i�vk�R=��Z��������R򋐐ψ�]Re��λ��ެ&�Du� w����x���'W����񕕕T@~m}��/����l
ڰx�K[4����hЇ�a��W�Ó��b�"Ԓ���v�Ԡ���#@_h|zz�)8&6vm�@2\5��b7�{w}��{���6���%��O���W�Z	w}(����q����ȡ����
�5o�����4P�%'��q�70/�Q�q,/������uz��߭1XBW�e��4lo��<@jrXöE]��v2B<����o ���_?��8�\5�t���t�T�&'�M��-�{�%�0�y���<,�K�Ȍ�җJ��Wn̪�tvp�}I���γn��`�WB�)�G�3����#t3���ɍY��n�]�7���ؓ�t8\lBҙ$[FK.M�33�Hp���gl�z�Q۝�g���c�� ��֖*�4ǀr�UД�DP�X�shh(�p	�Դ�c�� :eM�n��T��d�����q�ǽ$��X0��?��
��<k͕!�����\��{3e���+����D��{O� Cǯ[[�e�d]�IA�m�60�0�F��<,�!���Ʋ��.��[�j-�œ����˴[�q�&[����iα����4���}%'=&66�;�K(�<�!�F7��os�g�#w&�v{�V9�b^��Ż�%Ҧ������̬ױ!�&���䔳��o����<C��l�\�w����&,�����p��i�أ���I	Zh���S�a;�S����r`�ӵ[��K��b>(���-0$����N�`�9���b�P�o��		� �v�&=��WU1��}�.9��8���� o8m��'B���da�᧹�*��<�b���h�CCC]Gc Jn{���ב�U���m`f9����u���Q:dg{C7Q�㘭�."yx<9ժ�����ٙ�M������t��kie���]G��r�Q����b��ă���W9/�k(	�w�\��y�|ܔ������Ǐ�5f��Mwtv:-�ұ�`���F�mlx[V��M<��weF�cS���lk8���~x}bB�3���ۋ=��=����2��ڲ�؇�<Tz�J&����ή{���Cy:�i�-�W*���]���h�jF	�ͽ��������������YX�tu�6��H�+���Q2���u��jR����c����������3����q�w)Ew�j�2A�d�a}�z:z�v{��Q���A��UuI���Ovv0���&���<lfz��+ �)4 TJXH('?ixVVD!��]��F���5����������ojo�%А�1���:^SΙ����X�O�Q���h��n��əj0?�N�'W*K�wx��߆��,�㳳��P�)QI�. �>��X�<�ѱ���UQQS{3_k����Pc�a�L�&Z�"��D�6C(��K�q��϶i�	�����Coh�kP�L�%��5p11���SSd���2^nᑗ���y�3+�`-��b�8z�nq���a �uW���.)�åH�^,Xm��O�e
����}dDz���K��O<2?Ezۑ��X�$/��Ǜm����$�0�[��2�{Ɋ�Bǌ?�����6�i�p|��l*fX�)�������������k���^��X��6<T9�q@5�%��\��ty缤S����q����#t|q���89��8�����"���K����L�Q,�`��Q(
.������	����隥�����O�#���Jk4;c���j��A�ĠC����s(��� 2+��P�sm@ �H�K}}��u^������ϓ
�Y-�P�MN�� vvvf�.��o�4�v�ӡ|aa�FJ�L̴�?bQS�G�Wo������[�899��1��0h�� ��X��0mMXY�L������ϟ?P+�ȝ(2�"�������F��5��5[UTTt�{B f���l���h�U���&���R�:�ߏDFF�������lT`e��c]�ONN�F��$w��k���!ccí��',�L7�s��)zR��_��X��d:�IJ"�[툝~��e����v|c�����uv��nuB3�_BLAY9C�e���GB��:e������ԃ@țo�ݝ�O'������Gl��?L�
{�FzF��ך�v�>����Z;��&OE��~?i�{J"&:x��`�Q�{�|���i�������?y�S�[�  ��EC�;h��
F�H���b�F��$[��$�sp��i%%tP�\^�c����W�>�lI���ᙓCݴQRH��i�30��~f_������@G_����o	���LL�@�o��3# (������^2�3�������p�t�X�$�����w�pؚrWHN ��@?@{��P=-�Eu��&<�?�Ԫ5108�h�#z��j��Z7HNO=5���ps��1�áF|Rҋ|��R��JJJP�<N��""" jHii����""Ҵ�� �%꽌��'߰iWG�sȰ̓;DS�}2#��d�
%�A�����4��:�u�tx�r�����m�/�ff�ZZ>'�Y��\PH�N�6��\�� ����)%�j�F]���=Zn�!`����E�x��az����#�#Gl��vvi>U��z{��''nl���\�		�=����NC�Jdn�֮��\��,���ܲ.0��GU��^Au�����.޸� M��ܱ�W�X(Ne�zXUf���*�^���1��&5o%(����\LS3e�T(bEZJJJ�?��9"B 2ƫ�
R�����j�@�f��d�C�4k�`,w��$S8�G�!,������6?�8=23���7�Ny�u�miYr2!����Ě��t�R&����i[��܄U0O�7+m���m��5�d�͐����K��/3� ѯO�!l/�f���
�c:>Y)V)��[C�a�7}1�}p��l�F��6�=�h�T��,��6 ��.W��%���k��I\���۳B��y2i��7�X@{ ����4��~�z,S�kVH��?� �mŧ�����Ά��>-K�*+�
����mrb��b�ebbZ���CxIL
4���ɭ��
_(��tu6ۡ_Φ��8Xס���F����,@n5,Ʃ���"ҫ�L�^l�&��q�#.��@��_�đC@J���$n�2��cR>�B�3����Ĥb�����;3�U���KMN����� ͖�+<�I�H��
ό���*�_d���O�ntx9��4�G#s��m�s2�����2f�6�3O�gUS�Iߜs�:��L1��z^v�֍���x~��|8� �OLL�45//�=`����~�=7�(J)L�g0�����=�^33���=	'�	��u�� ﬛%��ƀ��V2��Vc����g9}�C'�z��\��jX�l�t�P�W[�0\�T�־��t�᳹��[��KMZ?����M�g�-�'����C��n&&.����T�rQ˱�݃1�%]��$<��"s��DB'̞�@h���=��Czr�����5CH�ٕ��LC#�/Y|Խft.�;>�zw�vwu�[�Z	�Z�׍���4usQ,�ny��`�Y�2,����������S@"�����ω�j���76��D���CC�W7�[��H�{�?җ���WZzV~v�Xe暼F����`nNA�l�P��B��X�.�ܷ��%7���0��bnA3��:�-���_M��O�j~8/JD&c����h9�Ȁ�� ���b��q\\\��r��60�A�|||�k���__/[QSS_�<�=y���r�7�
��MZ�G��*� *���;�������g+��_T��5��7�F�)�UUU�'���uV/���]{A^�e�� ,��"�f��q�#y�"������n��k������dF��뫅�r�9����(�q�Z��n�6y
@...:�r$���|��(��:�J�j�e��"*)�V��y��e#�θ7򜊈�O�UZ�%�/�ֶGR��c�0{!�������fVU)�� �t5�p��������kT����Q<��\Ÿw"^�xo�p�+�4����YԤ�c�@��m2�{"���͙a(g�קO�:ZE�`��]�͙�kk�


�:���CBVG��;|P��x�МM֧wf����Y��hj�sr��# _l �s�K����=��7_�v F�����84�fm*�0b������%�l��("D�{x��������E  ���(�UX[�j9ͅ����o�9CEK+��X�W.����NCC3���{���|�S��Of	
D��ӭa�d.��	Bw�d	��������ױύ$W8�$���F&�tj`B�^J��0_gen$U��(�l�I���i�O٩�QsssѼ���ޓNAl�1]��[��>-���%!���X��b\�=F�i�0���ޠ�}ݵ?�i��h�o�G����9Ձڋ����.�^�Kğ8�$�:��b�{וe:SJxΠ�D5��h���ו�iN�����5���/������1p��y$�ɠG��'�*,�р
>���V߬����+�k���ߗ��S�Q�KRb�ԻS��[��YN�ݷo����΄�B,� i���������I����¢E*0��R�k\��}rD�p��~~�P4�j���}�Lo
[N��}�4��e{�o|�����l�M�vYX���^����܎�.h			��h7;C�������f�������sPC[��&ѻ��M�(��E�R��ϭR��#�������X�����O�*8�Xx���#��:��9)��o7���}���
��qy,����"U+G�;�+���tc��@�twe��E�CnbeUަo����SQQA5�������6�XPP���/�BV8��im�I8���*�&7�r$�g0�trl��������Yjn��/���b��6}_û��{���p�s{���TK�)d2��td��V���5cζ|�ɑ��ׯ��6k�Ճ�P�����"��ed�K�4�Uou����
/��Lab�Ǘ��X���#Sz���?��9��w�]u�X\ƽ�a8��-oL0GKKK��K���u���Mx/�awtt|���܆����u��"2���(e�q��c�w U�Y���"5^iS������uӇ*yP�Ј7�1����6Zj�S�1�,����A,�8O ~竣�����|=���Bz��OA@@������l�a�i��$1)	�[9k���2 �q��h]L{y%�ѝ]2�& ��4n'/���r�萀����r������Kv�h���j��P&8���׀K��`�z�wZl�  Q$x��]��x�2�pu7�@]����|J��\�Q]@` ?�w�͌�=�s_�D$�M~I�I>�ɋ��-l<����F)����r5ͱ%��kQB\���rQ����n{1�=>|�!���4|�Q�ؾ����ޱV9��KEǜ-��6��)�pO�����e�{�ly�_ed�,RʁTo�N�Ր��w�+�i��CQwGΓ�4}�ǠxEJ����@!��FvV�E���3��fsB;u��S�������:4��Ya�%�^�3�R��E��^����Rf~���6_NBl����w���l[D3�EQ�XzMduu�}��&��F.���y�3,�w�B�m�0)�Ā���Qc�w����򩪻���32껬+.F�_�m��UQq�/�Y����3		��u�#�Ѿ����(R�LF��0[[�����
���E�U�9j�����
/Cc2�ω�BZRi+���ǒ��W�k'��ܽ���Y�(�`,qwޑ�G���x݈�w��������.CǈK��.q9�g�#58#��<��ދ|d�g�.FCi,E���19��z4��C+�O�����U��,����۫�d狾o^:-mΝe�)(+���L�M2s*|�v�.�밦��d�ȑ^ZJ3??����j�$)-���Ǵ>	��R[g�|||�����T߱�G�Uk>q��Gw���L���c�Ӟ��r
��w3J��E�Wc����Q���o�V__�V��{;�H(����1,�V��Ǆb�<��@\C:V~r�^���ى��5�U�J���
�NW�
rr�����K�bc}��
���{�=u�
m>�gP�(#�+&v�{Nq	�ecf��ₛ'
�mI�w��]�n��1!���*1<��_�ޅ��ulœSP02�ʱ�u��>X�9z����4
Ok��!������l���b�9�L���ثˣ`�<fvL{���CB����5ˋ_S�@ B^]oN}꼼�����G
	�l�OO�=�/�8м���;���+R^6�%~1���f&O�$>1���ݦ����h��9{���P����baE�A�5�)B�y�TA@]A5��������ka����گqN[�Nֺ����r���5��kg�%��F:�|vM�x1t�f�Q����6�*C�ۧ޳<&g��S�V����T�J����ܤ�L���m�^�%�>M`��{?�_����"���;|���s�ۭ7�����	b�=b��9����h�/ᬀ������Ԅ���0z*))��
�5W���7��"���^�w�::mJj��e��!pS( 21�W�%�A�T3��'�7.jjh�'���ܔ󄆅m��y�"z]{�2�ڎUU�s�:ܼs:�����cPw�*(*[x�k����1#���7����gýD��T_���[�#̊=?1��[y ���e����h�?y2PD�Y	"��A� ��;:������.��MM
i8��OIl�N������ybݞ��)I�WVP����������o#Y�T���PC|��e񈰞W�ZK.Y  ����ª`�ɵX,,,c��`�B��(_�D��ˇ���
���K2���/�+\��c� 7l�y\b��NEU淵455��&,~�eg���Z�uxza�e��������05Щ̃=.>X0�X�����w�N�7Z���DJ��ͩ�J��3�^F#kf�0�ܶa�mM�F507����Nfw	�~Ù
�z�b%��
рgJ1n'e��8�Ĭ��wc�Yyk�gR׉3��Y�+c�ZK3�X;b\��m�����J�)%��{;��j�,o?�2"##϶z���`�~M>�C���sgB�e���T�ź�-�o�rT�l+g)ɚfʴ+yrǍ?"ٗ�!]e5 ��)�0.aj�a�r���t���.�e��2rRu(�_TR����J�Q��d
�!�鵸���VI̶�p��𿧪������cb˗��=��l�k��sl��7�҇;��1��by�Q�� �F=:�'�}{�kz����7����o��7-��ͦ��x��q�0i+�?�XV�N��-*zV����e6l��Zoe��6k����L�,�3�{�RM��0���>?ׁ���v)\���L���Dtv	MBſú��5s6X��W�X����J���ǧ.��5n�F�=�C�K�R%+��*s��{��rINa!������<��M������a�ѽ�f�}�(�i�Nhي}�\_d`����#c��LdT���SV�E�Sy5�����z�ʗ����� �>gaa��&�� �2��������LHP����uIZ5ﳶ�)w���aff�m:Cߒ34�,rkj��_Pd������O{C�/����h9�&Dt�����?ז�����p�d]j���A�4B�]P``]�/rr�ϼ7�Q6[����6��*jj��g�n������FF���I!��x/Ҹw�-���U}���IP�%�m�=rz�G�{�c�>Jk��SS�-��� ubB�V����c���,'4���N�b����k@�9!r�^S�����?��{�e	�qs�Z,���$����ZYѱ�Qpus�QL{��9���%.+;���۱��l(�1��np` �b/ն��Ƥ	X��c�8�5b�w�ܧ���ύ�~�"�������|g|5�W�y{0�O����&<����"E4����\���g[ۗT�7�����6��Ͳ���Q����S�sf���x�c�ĸ+3����:*+Ѭy0u��1�Âw�CXN����j���f�=�g�kRqG�p�K饿v(/���Edd^���ޑ��<J,�]�P��T%&^
^,�k1��U%s�fa|���:��l��MLr��AWܽFFF��������1�9����._:t>B�B)m`��Z��=�\|Y:R
����6������@!O^MDHN"�V�+��8�� �,Z��We��g�)��Rt���BU���o�w��wǳ���0c�n��jff�Vɷv��=<,�r�������P3��h���*��䛑AF)Oz86k��Ɵco�������
��7��}�`TL�XAq1�TN�M���̲| ��=k��w�-w��w�����t�p#o)F��h)-��.o��Xl�|7J����/A����e*�	4��]��w�L�>[k�%88�U��[�GK��m@hwyX�����3jl���~�x4���= �[LLL�4�'��3��Y����ߊ+��!�ǜp~�9�Ӎ �W��K%U+ᯎl�R���	���j�_"��y	N�h�����@�R�6�Nd�����|}��%4===�[��}�+~�u#��}v�wt�S�ޤ�}�A������{4�dkkZ������ڬS���{~�����=���[�W�����
"�`���#9�F���~]�������?a��̷�B�kq��Ԅ�k�0��ꆔ2<���f'�����Fo�	�jp���i�8�dB*�ʧ��'YMm���-�K�U�{�̿?ᤉ&Ojӵ�88Uz�T�寧:�(f�0ih�~��W��tW�š�I:!��%�"���ADF�䶸9�t�X.-6�Y���NNyo�x10)8�t�#ѻu's���L���,!�K�8vS��]�ݟ/2����[	9�k��DN��LoP�R��MI��S�����X�@���T`��#_�Y�.Q'~P����`���ǟ�@D��c��.�0hI�'�	|�1��=b;���^�̌v�\)�p��QY�bF��j�szrRPRuT����ߡ3\�i�ш��jʦ�X^�'�t'�����a��r�0�	����*�c!��tЎWuuu���G�}~cc�5�@\\_-{8M�Ch��p�a�&!~0�=�!�#ސ��S������0p��r�"Z���������A^�� kR�tnin�ʾ��_Yj���:�'��l��lI���揖�
~�������N��������8�{w���A�T���r��,�[����S�>HgB14����E����@��4���,��z|9�K���&e��.�<��Q�)q�G�,��yc�\M�HOK��W��)Ee�38�6ܽtҶ�1�	Oس�ۀ�;6kP���,j���YYP	��u��̀�ғ4���c%y����kˉ�LO�t��� �^I���d�
D�u���컺�D�͍Q��;�h��Ol%����
-B!��������-(,�+��c�84�
�ս� z͆t  	���q|y�^�c����!�B��׉ Q��:�صL�n�����,ml~���q������j4ڣ��8�~������P�����a<!!a�� }��L��^�xq}sCFA��ð.��{�\���4qA���	��c2[;�F��˔��O�P�`Y_Ɠ"fF�PQ�k|~�o�� P�g���c�W�?
�������;�q��������a��cbe.�J��rُ�污�� i�7iD��8�>��%�|y^K���+)����zK��G����� �6�	�d�
�s���l��{�D{��7R�sW�0��4s���CT��]�����Y��\��K�ߤ��\1�����M���}��q+>���9�����WZ���<��U���%O������P�#��2_����t�S`VTVB_?�+�y8���4)�������r+�������Ơ�5�����x.�R��J�q@�ϐ�/T��9L����������(txLc�zAA�ջ�@�<�߰���#��h��K���3,���w�Ƌ�jsss�CB|������)���L/��~��m��~��b����.<ꛟ 謚Z�**>9���/{<�8=��[����`���8���XxxH�m�f� �Zש��N ���ie姷7l�i
�r��֭Fߡ=��q0L��'��u���Z�^���U�^E
�2~e��i�L_5�ׯ_I��҄IV!�d��}�V��n�wƌ���Ĭ����������*�Ó�e��pw2�DE�yx��x�nm76Y�MpO���m�^�|����ކ�}�N�r�?���]磤H�U��0�]�1a��X�rw�l#��̓!�TcU	��G��P��^��ɴ�[cL�+J�o��H�[���>W/M�C|�ȕ.h�������]ez�
�kVl}�~���\��u��0���]���W �Km��S��/Q������C�������vr�RP�1pqtd��<�z�T�������	�ؒ	���t�ga�4t�H-�c��u����@d���L��f����Ғ�y��b���g�{D66���n����̷3i, �|@�u9ԕ�V�nݵ҇��>/�*+���pĒ:�r���F��æ߃:�	$��b��Gf����LLu{m��J�Td�!-���AY����e�iO�x�����&9���^ �����t,�$���a'"*	�gc�(�̜$=K������k[�����}���?wl���|nN�[f��T�I\�=�x��fIܱ%�w���Q����� ق���?v���[ʝ/��Z�4t��~ĺ*Q��&%#�y��4
�����K�-�q��V�0W(�`���ur��9��w8��	�l��v�P�V��ΙM|_XT�	T.�i���5t:��	˯��uC���GR�J���+)������L*"�_���@̇ l����9�����p���5��c!�0�z�;T���2��e�vh���nm�A���������3�>���+?{<_,���vY���+ ��ή��`q��������IDBB����*�t�f���A���4^hÎ{p)��01o���ީ�t�X������"�@RDqI���,#5�	���b��[|��#���*b}�W��]p�G����a>��_��U�قC�Lf�k#9i�������[��R�BcYz��t�S��%��k|��Ѽ(��7�G4�F�f��0���c�1�LL�rp$(��)**�l�o���`�5�0�V*K��c��9p):::oۈ������������<�M��y���ݒ�/G M�
��tKʊr�,<�������+���}J�R#=�hdŘ��&�J���|F�9��2����|PN�ͥ���~��k�`������%���b5�"3��P�C�� �ݻw�Uh7�������m��3�?�k���ud����G�0����I��jV�p�gCD����֖ػ��iFQmr�Q�c:@&..�72",/����Mn��YT��p�
���53��#�j�tt���������,D���;.���[V��q� �wS�n�ONK�R_<<`D��2l�E�~�o��� �CWO������
t}��p��m����ݳ���2
J}���>$�{���	Cԝ����ԗ}"#1�ss������
Y�lllN '����сg�8S��` \�?]�L��������Dt@W�`2����"<��t%O��' *Zi.����"611��8<7�,��� ���IY���@.�=.���a��͙e �yEDD7�
H��c�rYO�P��B�/�Tb�CrK)%,�/��Kq�ի��d����l�`G7���^�ms�}\J��ڡO�N��LQ��9ř���
��5呑���Tz�0X�.���*�O:/*)*��E��Z|pya}��nd�� �3�������/Z�������n�Rֺ�����͙9P���WYy5y�Xe5�m���o�Uu��>�`�/ZI��2�9��5dVd�VD�44�������˵���;��So�������%Po��� C��b�:|׿ր���K� b"l�aL=�ƫ�!6s�7��0���0��X$��B9�vK&�����v{Ӊ�xxx���c�	�`a11$@��б�Q�
���;���`T��[�ov���e���^�ľ���������U�c��~HOa���B�<�6�)i�*���4Tohh�w�?������R}����k���`���҂����í��ɀS:5oඐ	2���YG2K�0���\����v�0?����\퀳=\ăV9.�R���z��7[4~=�����*��·IΟ�UT�"�/� 00]��@���[���ӕN��6hLL�w>�!���z��Z��ÅڗPs������h�K�p�8�,����j�'�H���^�~���%1�N��$��Rȉ,��j�l�_�2!&r n��fz/�����ä_��#���}��i��s�t�z_�;~��2��@4VD��dd�)?~�C�Qi8*�j�C~>U͂Ϟ55ץ������"�(�_+�t�Ɯ
`�2��Dn����
y�H��<��F�s>11��?�z��10���A�o���q����=H7���pV@3�@@e|�n)��7՚��1����Į�[��u�k]��i�⽓��C����椳��lKC�:N9�Z�C^����O��#����j�jj�x�懺F�+^bb�k�g�[x�K��bIn�� _��tD���N���PVVa���Q�mm]��A���U�:X�EDG>Zj��m����!�ׯ_�nW���PH�'%�yp@���h+�����4�G1�T0o `���!�Y�P?�����~>����g�v���`ccjWW�����������\P5@6\�����%;��{%�Ԟڦ�o1fK^��Ry'���-�vvv �Bb���?ˀ(~�Wp�L
H����A��T9�_���9����˗P�#3)}� �6���݉�ȸ���8A7^���CKI)љd�^FP�I$gPB���XN=��̔/^vF����F�0Z��C%d�ƖS>Dav�9�T���)��Ȩ�(!J�T����G�{�d�S�Q���F��Ō���ֈ��V/a�#�3��*2,�������O�%�C�������W�pwww_���u5m2�P�7t��]�Ztbb ��P�U�����P�w ����%��J%ڑ���_���*�ys�MEE�������y��š�*  �?((J>�#%��k�\?"<�'��Ģ����#`-��=; |��Y��U�Rq�Q|`��o�e�&���F�^p(�5�l��^"��哐�ү�0��w3�I�*�o�>��E X9Z�t#��zA�{����/�g໦��Dȃ� �������$�^tS��5��C�wQ�b�����s[�[���Ǉ���g��ۀ��(,D��O ��uYv6l���5�܊�Ȭ&T>X2������s(D$%%���ffz[�Qddd�))O	���2,���~�/'�Ai���Ͻ?K�S<�� ��V*Ӣ��2�ǣk��_t�1p��@u �� �7>>>6=��USUE���5t�YD-%������{s��k4���	��p.�ߜ����R��ۙ��UAx�-�1�{��i��[f���w�3��$[r�A�v/1C�r4��v|y)leŸY���Pg��F�`��ۙ(e~V~Z��zRY�R}����A	1�LF\���<bd�)�d$d�VC}=T�޵�B��y���_��5��a�wlG\�?8��NFa�-�}����[(��`�� jhoRJ
D�4���F�\����q�X�W*�ˀAds�Ą�d
'6`�X{���@ff��}|s}}�n��\�:������4���}��鲿R��/<�V�?�ld�GMa�G5���e?�5�.<`�+2�C�4�^�f��;h$=?_4�F�!r�E�fV��
<�p���ZT�9��4���h�e��u�ݮ羙dF^�d�7���-�����%n{�1�`�jjj�S@������`Bw`�٦���6%v	�Agw"����L;f*��")�_KK�p{v�o߿���#ya	��+(X�W'��@"E�����J6	3>���j��'T�Y�]��`���紴�٭�������!]����&vL]R4��g�|b��W4-�W�����H^?����TT�Pʤ�N�@��,����o>��W��ur�цS���O*-��Ί)����x��ֶՖM�ڞ-�?�����۶��Q2D~�;��V����/�<i>�|����=�mҒ���/T. �E�x��9b��0P*)�S���;U+����~�u�Xn� ���%43xE*�ӃA�"��� |�ʡ�oooD�ޑ��Q��:m��d.�<N!����.:/��ܒ������S���a�]�bU,��H����]�y��u�c��??�N6��A�chJ5e���w����w	.��^����2Y�	��W� �Ο�DF�$���C��Y�������m��K�� �|�&��]��ru-����g!+��JCX>��KT+��y�������"���^�ǁg���t��WEŵ�nخ���GЁT1��ȑݦ���	�o���/}�����&_Z'Y"�HHH,69a�����w59�A�j=��>dx,_[Z�7~��P�F�ڱ٘_��8���R��|�0��GK}���f!�;���ud��񒔀M�+<�Ui�Xa��Vc��Z0Ȳs;ü	���lB}�`����un�w�ˠ%�`BL/g�M� �N~e��3�ȫ�a�\�/�*�L��ax\.��f��>�180��r�KWW"K볈A�,��$���0RI�P�t�I��EB	�'���ML�[#�~%��mS���������Cg�C#"^����[�ٙ�����j_XP��)�߱^�k�F�������o�����0������)�����o>��UuB2
��ߵ�
	��u�7�[WTZ�1�!�}��0%�x�`�Z��f�0u�QX�?Y��1�b�f���@��ڦ&BE� �}���6��{���U����CB� 	zk����BW��x=�AʴU:��\�D���=������~��i��#�ς
���`� /� vڥ�y>�B�è�LoP����i�t�͟r}��%%�:�����r�z��+�?3;6&;�ʣ��200�����|��D������������?]��h�Б���
��.�����Q��Ʃ i���C	������>_m�?c��sqQC2�����&�šȌ���m���N8FD(2�WBꌘ����/����n�uu�P��߿ewX��ơ�8���ŭ/5�@����i�N�D���.{7��r-22�K��W����H�e�I�]jrz[,�P���3ΔP��l��ُ>UX���e��N��#��I����ۦ�����4cV&E_`}L43�Cz�$��3"��PP~���n��I���*�6�6�S:۳2wvŎg�$�&��{<>#ȇ��6~��g�b���o��iժM�XXX�&n�A�unw�k���(G|������P#�蘘�:��KS2� ��SEBj�7_\�(���03+2�U�Xl`��G�ցn<�=�$i¨sE���s��� `rjʇ�C��cNz������y*�0��y�e�t��������8h�(;�|��HMEo������<���	mC�#.=O���6��^>�/p�m��/777ߖ�}~��=ԗxzZ�f���I��PVn�:�3����������� `3����f������6���!B���es�kƙ�WWo��c����u��OO1�}�strZi���ϗ~�����i$0\�ri��B���\;PH;v�hh�����䲷>�,y0����CR�t�z��I����Agq�k���r���� V�� >U��H��L��������%�B�JV!�	!\{�QD���3#+��d_{�MV��{�kS\[f�������ϣ�#.��>��z�s����K.�\ii��Ƿ۱qq�F]�;�' �>>�I�������X�,�d��O���̮���|��۷�I�JJ!���ͭ��qj.�^u�ƛQ��+��1E��/�8-�d��	���á��К��ʈ�)ͅ�G̖��~�s�O�h�W$=u�}���D�H���+o=����yrZ�K����FB7����֓���ҒM���y< `-���Z~&�@�m�My���|ݛ��/�َ�࿴��C,z���&V�������"}����i�,��f)S�X��=?���5�Sz����;i�BB|�AW4tV6o4�▎�_�~�+����/���Y��){ڧ�2�3Nfe���֏�tlC|AŅ���Y~�;�0f�[Շ��VO۲z��O���� OR��OA�(�=PO�_�m�>���j2Qk�𑃛[u��+���VT<WQ�AAA!��ܟ.�ԩT!�����(�@mʹǄnJ�������|���U*�b����V��L�>P򓁨�y��ݗ͕�&j��&��wPMû��!� wRg||��lۅps{<虉b��{Ж~VfJ:����vJ�4���n/�SD�=����k:p*H�WKTQ�*t����]�EE�2z���=�z>|o�(� �ٯK&��B~ ��z�5��]BJJJ_߀���_y�N����#���d�	�
�����]��M¸DEG���d�ߺ�.�z�9qw=g�[��ʛ���D���*�Nl�wc��!���M%�,0���y��	M���e���)��b���^2�f[�23�?����N�Y*����s?�l�te�=hckKTO/Ic�v^��j�����9��
�j�3xt������u�m������ڴW�wʀ*+j�Lz/oW�D��WXܡ��!C���Yǧz*�5N����ؘ�f<������WAA���y���)|mMHQM����;�oȔ�w �[�%!-�(�"2�ȹ��Z<�	j�
���.6��TBnA����#���K��>�y�Al�__<(~��Z�n��b�m���mm瀱�#��+u�Ҋ�B9u�_��7�?����Xc%�=Pgө&�a׽���V٭�s�;�:"�~���c� ��IWt:�clȑ׽�!���؋4�º��Y �g`'�ý��qC��q	�];x�� �(���ͺL���$h3Rii����s�l�	�F����p��,�Y��<u;!�On�����0z���$Uss�-^[Ԉ�����U�<V`��K��u :�o���
�Y��8L֭����t�	�=t�
�*Vl<�h��W���㱲}0�e�����Y��hä�oL�����	>~����������O{� 8G�H�;j�E������o���Y)��@dooOHL,�Г�^i�_�_�6���׶X�'_n.ɠ��K�K����j��D������tܙ�@5~�T5.RR`���`���a��=�]��C`�H��bs3KK��	<����ڏ��.@b��ßYTv����V�zV#��������F�N[�#C*����W4S@�c�<��]������̀j�ڲs���L�[��Hp�8n �
0��}�����f��vS,����p���@~
4�PO�[�B�(��k�FFFO�~�A�dP))��ֿӽ�텥��K��4�n~T]YHe�h"�����Ej=�&~��Z��[P �?�ŋ-ي�m�&Іb�$�-�8�`��墦6�������4����J|vK�y4\�c*����顳I�8og�8H�e36�i�8��@/ʐ���������N����gE�ןn�㊄f粬���1���Ћ1_4�����[}�����/_�^]���d��Tg84>H5@�m���/���=��v���Ùy�g@�o����	�9��z:��f��1%�o���A��?^ٳW���̜�Ҩ�է�y ������ied��Ϭ��l���"Y.9��iσR `�����			I�_�H P���+#%��� Z�/U�a=��>E��*�����-r�V����i�g��7#QL,E���}�j	�$l��6�J˽;�:::z�����}���Y����A@o���2�\�����A������$y�����jt�������HN��z����u���3PA)�vPZV����Y�SJE��Wa��@�eg/5�L<���2�؇F�#Eax�66���0@���SL��ƃT���O�0�	����p��.d�y~AA{���� t̫n���L���~2����϶4x�.�� ��\S���Y��/:##��.?�%� �52:�S�|�#H�O�!��#j**#�u���o�h����IW�<�>zU��~����g]���-]y튊!��Jf�܂l�K�o<~l4u�)|���Q�z��Ǖ�o��?�u�u,���Od.G|sX�5��%7�3�-��0�~
G�קk[�<�s8r���9�ꯔ%�7�)�r��{�N��C�(�6���v���-$g%�3Wa)ÜZ4-,�Ŧ�{���5v?#�vYo�J�n��������|v�^������z��������M12"b�m袄�A��KO�� ����[��� `�}(Q}�E�U��y]�Պ%���<q�H��[}��͜D���ļw�h��%NN���]��'<bF�_lk.��¿��~S��ێ##�&���h�ݨQ�������O�ܪ�@=�ϔ��qyf�Ͽ
-mt�3���5�-T疡�Ýo�z�富P ��*}@ƪ��<�,��o}������?z"��=ҳ{ξn�h�wy�e}�İ��cy��/c1�l��n}e���kO�����R�6U��^��4�0�jeU���{�O�QRJ
ɤ�hƿ�X�Ů��6�ǧod���8{*����Qx����Z`w�0��K�������ܼ_~tAm �!���M�4�YP*�Z_�t�c@�6�!h�3�74�3��M?�]�Rڅ8�e����s����z�����C�����-��t�V-"'�U3�|}~��˝��5�K���&��"�L��	p祩ӓ���e�ՑZƭ3�%�� J&s�uk�{2e{��C��������=\����rw��3הּ,�,��f�G�KC#�][�7�u^�ٹ\�	8��X]u�@��5Z�u�ˋe��|6�:��m�d)�%@�l}�o��G@d�H�SU�t��������}��ۏ��:B�}.\����4�zS�55�x�5�P/>�� @m�v�����Q����ҳ��|����O|hJ��ptG��.���.r�����k����>t�x|�����C��7�j���T�E����#�98���i�7��09yE�Z�ߛ��_щ:9�<�C�3o}e���7 �"Z��[_i��;������f�_��]&���U�۝�-�VM=~(u;�d�K8�δ7�R������9le��p�y���rPΫ�5�� P�Pꤋ��v?�2�d+.�U�?��`b�=k�x́���1�n��W�|��U(/���v�N�ra����o�����kp��_�, �k
�v�X�x�bdrr�ё+���0��v�C�8���0�λ+9�T����=R��Ԕ��$������E��uk�KPۄ��c����kf�K"���ʭ�:��������rb��3kz|���g���U>\�[��=>�+**zel��]eu�����ԯ,/��A�F�������r���r���E+�����p��/S-�����Y.j슬l����R��턩#q�a�>�ߕ�%�6�\�ߒ�{�`�tͪJ�+�3U55�\�����ccoe�P�F�:999/�dm������K|p3���`�XM���+�g�-.x��rܪ��C/_��M�E����w����@��mu�,i[sIяY`+e兎˓�vG������Ğ++�l<�5UӍ����f�M�A1�s�������z��mo�#�|�K>A����~$8��,l��Q��?}������E�?���|��r�K���Ӫ�rz� :��������J���~`<G�xs�lO���Z�<=����� >��bܓ~�{���I���C���1[,��X�����1�f�^��B�DO^��)���	�k��[\��^�{�� xCk���lG�i��.�r��e�����cJ�yȊ]"c�3/j�1���p`�������1���22p�w3RR��B,����q!>?�>�'�%��#ᱝ���}d��g�O�Q4Z��h�"�I�=](1t�oBb��`�@�D�[��H� Ƅ{� ծ������~�o���>�10����B�p���^��x5�O]�4�^\Vrni)���^wY��9YI� �k����H�L�E��]F^h���5�%F�^Bf���F��V=���δ��lz��	x�h���61L	_~v�$́��n���:n���031qR�Nd�X ��D�N&r!��ϡ�E���d�LC;Y�`�����&\d;���׏��>n�>����ɮ�����qqLYS��ܼ�
�C{ˑb���"@��;�0L�6��Q`G��\��a��cb� ��������H�u�/qRR�����ݞ���ͬ��C�?h���ۀ�<�x�����)WMJ}%�4/���X�������z�+\��V�*���jt;q�K>T���rG�ɂn����K;����̌��M���b@���-Y�K�LMs��IE4�c�g ޔ ����F����%����ܽ��y��{Z�XU��O������}����#kW�@��MxEE���9���M�{�FU%�{�JU}�3Kb��`$�SVP���))���B)�D�>�VxC���OČ�x��&�1~���x��x�
�$��ׅ�sR�ߛ��S5�rl
�ҳ���%g~��d���kH��4�;���f���|�^h](k@��VN,6��<�M���wQ?Ր��v����ܤ�T�-G9�������2bf* �2����7��v ڐ����������@X�b����q������:����tNN�;E��PXI�S�e�h5/잻۝���?��YN��7(�Gm�ُ��!^5Ꞿg?=9��_'�������.�;��J?z�3 ��0G9�b�(��V0| |��:�_���rP����@�F	9��	�+}�b�r!�-�zTt��☀��b7�� pn;��oL^M��E:�og�}�j�c��XoY�a�BU��Ȳ3V~��,���?Q��`�U�@	ąu�y�A�/홄l�
�/$:�����uF�D%&��9�?0�;�w~�k�)����s�b���Zpe�[�6�)���u���I6�	�+��x�2�����_00(1tդsބ���B�Gc��O�����_��(�JM�/��݉���G%��k;����/��i�?;�t[��AU�XI������\0��P>��T�M�c����Y�W�L����N;;7�S�t,�༃Rn��[�㓽&u))���)�=h4�/�@wv��=�}����T/�VDJ�Cy׀~��Ox�2�+$v�J�*װ��j`1� ��Wi�pr01�g���Z�}��|��y��JY�go6���,W���2=`�3`w֧��>c��>�mo#tm�I�*-�˖9�V&��(�#1���D�f]� ����	iH��o��wX`��XU�Ѯ�Z��V
������#�`����7O�;Y�����z�\�&���$��ߎ`�����=F��!��Y㜲׽���s[x���tB��fp���/���k����uHR�X���$�nb�uu��k� t�o�v��2���]+Q��-����5=���L�ı�H(n��<}�]��3��F��;�v�����L:���i�w���������d�荭�P�l���;�|B����Wp�بB�˹e]�
��Cʋ��Vy�W���rGͫ� ���J��c�㹾�-'��a����ZSccc���]f]&B1��H9���/�z7\�N�x����
___ ��~���[ٳ���������5�>��[�7/�HIKW������ �2�x�QN?o�h�A5D�VIDD$����o��YYY.]8<@~���?<��1A9����Va������Ũq	70��袤l��"d��_`�d*��}B�Յ���qD��$���
vvve�%%%����vW`n�����[F�筝�J��"M�İ�z�(�.L죶,D�j7���w��[��L(4�`a�2}*�T��'-��KB�:,����7��S�\��~��L6��d��r}���Ϣ��7��1�ZHʑ'/)N�t���e�z�QQQ�����Ti*9��'M��w0��C�v߁#_�$������>ꆲIOkFK@ԏ啐���$]��К���~1�8�:ŀ��]
���X�ܳ���2�e�sfF�q��é�Ƈ��s��ZH.�p�>�.�L��Z�Fq�r|��1*��.B`�ۣ���=����oAf�m����>�Mz�1�4BA$��o���A�8�0@�I��n6�u��Ez�z.�LY�@�BJ�R���2�c�������_	Cp����Y�G�#ʝ��!{� B���l��1f�����t9�J ���B���^��>Q%[����27����gVV���Z@�p�%��=������>�|�~�Ϥc���yb2p��eƦ ,�?�J�;�N����^��SĠ���_[�Y�jj|T�a=B^��Y���N�6Q.x���ŝ�\����iI��.��fH��}�8鲮���;�a�@��L�������}�@�3$��"4b@M�����0���g�#��p1MGTG6���jI.��(��&j�hiEA��5y4A�c�,�r?��[��ҾS�����q����N�ƣW���]ɫ��E~��w`�y�%�ͅh��NuLVZ&����D;�)	���U"ኜ�&���߯�3���O/�߻���][,I��_�C/�Ic:u���Nx�V�E�������}�aϛ���-�Q�x$�n�m��B��ލ�/5J!)ٟ�E��mmO�B�9)񐂚%��|�_�2.�=�"�Ȥ�����7�E�o�5N�0W�Mi������5a�l.����l�!�߈��~?ZYp%o*�8��Fgp�ڞsJ����מ7;�BLU��ƚ^7���v\ж��� Z�Sg9I�j�����^�k�|0��M�?�x?�s����&�٭���h$����3�[�W����4p4�4l�����"���D�'?���6:��[y��OUU����I�J������ϋ?�e�(�3��T�q�;Ǎ���~���J��<��<}��q����t�ߠz*Vp�E�D �(+�=\*R�W�2�g �%ǔ�暶w�'.��
���R񌦵��tF���Y.?���}�Ҳ���0�P�OݟӉaG?�	֡���|����e�/:<ȶ\NF�Xiv�`(�R��F֑1�ku���uF��<V��5V����B����#�dO%[���e������8zSgK�q���hD"%o��l�}�xe�u石��QX={�M�^��(#�����ƚ��(s�y������'�����v�� :J]��F�`^���1v����GXN�_Ļo���U4�Ӈ��.�ģ��ڮj��Ԡ-$�)[{���-K-�/��c��2����LC����3����D99��ڕ{�����,�U��M�1*���rT@�(�n�8��/̈�V���~�
��s;�:ݗ������SYp�M�藹��5B~"?Q z��]�D��'�N��O�@|�U��tz������b4*�Q����#W��15�L��Nr 1���}W��tt(>�%���(��U������R��@�ʆf��v�����畢�~Y�+W1$w��[��\�=��x�䰈S��8/2im/�M-���m��&�0�7$�Ӟq��Q$�a��1�e�F��}��a}�?�9>�m,��ȵ����m�66���������H��>�ی�� tq��=o��+t�����k=�&�\Yp�U���@|i���Dz��	��8TK���PP�: ��KL���H$����mFFƦ�o*���%��ޅt�a���0l&<�w3�ƿ�[^�ɼ��y?{��r�
�����nj>aY��s��s��l��;ך}�F���Yna��m�tf��Dk;�u�\�V݉�C�ھ����e�,lC\k���4\ibdă�XM�- ��'�����,�.8�.Q��4
���q{�.#4=vN,;�:������ѨE�@։�-1��P��f�z������������J�Ʉ��f�j�hD������)�t��u�J&+4g�x�99����� �ϧ��ӳ�khd�&�����v��=|�'�|Y~������]}�F�Vi)[�J����{�kɃpV#���T�Q���5)���5jKٕ��.Յ�����nų����<�ᨏ)�n�A|���d��s������Q����#l<N�i¤�����ӌ����ٹff�T���<��s�/����\B��e;+�H�hDQ��si�,U��y�okt�j�f�nu~��:���а�V3�F�s�%ܘ�,�e�z�;���׈�C"*�;.�G����^dgKz���R���]
������R]tH\��@zGe���{���ad/�x�}��HS��[��z���k�V���AÁ��_��ΆM�����>�em��K�ւM�hF����JW����s�@Z�?��jԖ�����O<��N�k9<а:�D�KF;:��;RNN������&����i�k�"���C)�>�F��RLW�ϟ��'`Rْ"��S�ukMp���^b[�����G���[��%�ߑd��^<�{b�u8��#3%��\��%v����R	�*�<=�R���$���v K>�x[Y��了���Q��O)DG��������ȌxTxh�u�;ڗO�En�2V�����گ��0Y���ѭ3�j"�� �ˍ�ɡ�)�����e��<ٺЃ����	��b�\��⥰
~�c��d���5L�)�2�@2�	�i.\����>�I�A���+XH( ���tTJƦ����߃f��+���a���b��h�x�{(O�����#�~���������_��H<�����]�*����M�D<!=ۍC�Ao�����~��򆌪j��Ta>�Y�������8#��0Ry����Њiz"���ȷ��	��.���9�E M#AA�a���(���t��4t>��cj���$L����W��<< �A�,<��(5���^��c�r���j�0��B�:�Z�6]�I&��6;�5}��#e�����<��S &�׼e������6������ٛ@���Ѱ�q��d	���ׯ��������}j�h�V`�d<���;O�o�|��|xLN��Y�ٌ��{�le;@��(g�����i�����L�*f����S�3$�"�0�1�8^�_��8#��h�s����֛I�e�Nfǽ�4���i,�_1�V�R��z!�r&���в�XUh�&m7�T>�L'�.޼r�+� e���1Ɍ��ɚ:xՉ���x��z��m7��x�~����� .��b+-�ut�z>8B�28Baw�3>	��Ho��?���n�6�O�Z�:C�>����D֯p�艱�Q�ߋx� \�,�����fĹ*�PX�l�ފ���x*���0���2�d!�򘮭K��A���.&|(i�i1Q;��Z��*'��B	�t_aMS*�I����;�:�T7�G�Q(��5��t����(�ܷ���C`�H�0r`�<�pH5>�ꀈ��as�=��T�2l���<^(���WRRc����҅8�ߏ�n*��r�".{�QWXM���O�ˢ|Dy��[�zR���<�Az��q1�~���4�ۋ���s�X�V�ɰ��k:�4,�)`�N6Ck�B�e$�x�iI� jx8m�������o:�c�mQ�S�ܻԹ�%��2��Ȉ�9�&O|Q���e)��`��R����5c��7��1 &S�ygP��ƦEDDċ�a�b�I��P�������M�
�Ln�kٸ!���f&�˵P`S�vo����ٹ9Y	X=2,��ٳ�~�����Z��Ӛy���w��@@p�Cʻ:���<nAQI�]ג:;�+�����0؇� fNN���M)I�G�R::ǽ6���8h�匡fAIH��o]̘Ό�=��OE7v״m�$��:�;�I��)�=1.+2Rn�C�9B�s�-�Tw�Z\����ᨨ������#q���!�"eh��%�~z�t�X
[�����J'l�}oj:`3:"������`_Nᑠ�P��>�N�1����}e�pS_�TIU�n���o���{r���y�����FE�3�(�i�r�d���ɱ��P����9ػ��� >��-a�+���US���;wrA�E�"��Lɠ�K%�}��0���黳W���4� ;>ͮ�����$#�l�vV�� �k��I�
�<nA܀�3>��L1_��do��|�H}Ftm����� cO�}<��S�|����I D��|j��6 ��E�4�L�y{��V8	]1�63ϲ�y�QI��m��~ �Y�� ��;�S/�R�u�����M����0U�&a�%%�+���x�B���X�H3�$ۊ�-�S^6Tk��j>�2����
���A���Ը�('������s�2#y�������@/��).V ���cJ&ԓD9 .s ��T*�k0Y>��X��m�yzv�yS����@k� ��hhO�j2!�.* #Aȓ�J�<�A�����n��=�'��Т��?�>��˜�fiy#?��9Gz�9I) �t	j��,���%fU��-E�n�G5 ����<,����٪�w�Z)Q�/��2	���#�n��S�T����"��?�S��ж��V���������\~F������Z�����Ȕ������� 
�t�s�n��ap��%�5�����3��W �Y�z�'U����4���kW��fFN0�s���L�sY�VU)/�!�;ڷi���/�V{_>��WH���J{[�������^( ��Y�l�Xj[9,���u!�4K-�+-y�1����������1]�Vy�@�NEE�+.-$�P��������_\K��Co�h�r�������T?^ϊ���f�ΡH��;i��z�J�eob�0#Mh��p�y�]��1��,g�jqx����)�TUTr�w����yy��K|k����P'��L����k��r�F=f��&V
�'����?TTT�J<!�xO��eNJ|�xS��^ʷ�������t.���+��:ޱ8�E�|������b�z2cչ��pils��( ��j^�r֮�Hq%Ȧ{�.@�qS� �xD���<�q�4�X?�ޢ����e��I�m1:i��qyd ;�s��Kg���Ebp���d~��?4���m�&���϶O(JY�4���l���6��Z�Jh�TMm����������%�,)�Ph�6s��^�7$�~X�~��m��r�=���}es.�j�ʝ�$c>�ű
����:��nϪ+Dʌ4w|�	m�M�׆e��'��r����
c�t�������cQ^�0�W�zc������'����.��9����=}����5��ڟ��3���5�B��n�/wn�<X��9{��;�Y���%v��	8 Ź��VfFFg������+(o�%؛nQR%⤤{OS���}�=*U�K�rim*�>]�=P`��R큢z������Օ�Ԥ]e���'$3++%m��h�4*�?��ME�Ա��\��@á5���Es��<S�|�r�Y&��}�
�:�%���B'�l3|_X0�Y�{3�;��BΗ8�����VW� |�[�(`/���Ps������B��po}`*B�/����Z�ϭ+�/U�RZ/�dv
]|�_���,d)���� ش+et��c/�ٞ���a/�sIu�ƅF$����}$�gaFBqΏ^�}��zNϫ�m���~ Sa1Zz�C���>=
���:
us�?Ǵ�x�ӫ�����ІҠ=h�j�^;��s����鍲��w6G�5��W�ł#Td���G�kbbf�0��}��i�T���6.��t�cG��W/:W�Y��Ԍn╦YU���P	Nz&��K������e/*]K��ҍ�$!��|��^k�������&�r��e��_���������C^���{�5�������z��^6is���I��Ӆ��.�['�N/!z��${�y�#ph_յgCy����(�Y� ��ā����7�Z��>�}��ǈrc��LJ/�f�{��G/~�sҼ�y�9Ek�
�h� �e#� l%��O��Ĵ��
��da��$��4�s�����Թ�aT�Q;"0��ƴ���w>�x��lR��\),%}ܪ�d��`u¡q#���n��[N�C������O�'�S������']zAy��8�.�L�΀Rs�8z�����;jؽ盛�������s�V��Cd���'��p[�u�-�
iu��֦���o@¦��&���A�F!�G��3#��D�XX����_ʰtxp��Ắp|��_�TUӫ�]s&�3���
ޖ~�㦠��*��*N.�m/��>t�C�n���aW��3�ܸa�l.���.���p�]Z:��ڇ8��z�Y�Z�e��:�Hk�d�s�f�*��cŅ"�X2�נ\�h>I�	��^(�g���c�iLn��L2��y��Z_�u��' # I+��ώM�5��	�e�0�����C�_��\F�$�e�WP>o��܁=�e���Ś���@�$�r��\�	��y�[,������7�����܉磰��z~���F�ՠ����fy:���Kt���hpY����P���,�������<��+��������'�X�z+�Q�4�َ���zyB5�7d�fq�̮�~�PO�;����4���/jh���+Cr~~>���hf�n���]�j�F˲p�0׵�������u�&l���%�AR�u�r/=beF9ߨ�+��8H�j�o"�q��\l吀	gKĿ����d�wE�A�$��?s�#4��~Qm):$#30�t��+��C:���X��̛��ԛ��}�rIr���䌷=���i��Ve�ǘd�J�71��r��C��
�C@>Ў�`rn�t���� �����Ј�Mԙ��;�n�	I&�ܫB-�W�|��v�j� �v���C�Ir�VcNK;��O�ӟI�^�
�k�S����[�!v^f3m#�5�'�{�Go[ó���.�����PP%yp���=�rR�w
;�.��І�h}�6.�8���/n��W8���)7����pX鼧�ҽ㣅����j�ήGd�l8Kx�v4{k��+J��HD!J�L��r��<?*gIb*��F*Ga?bj"�{��9e��w(jtj��E�Oފ��2.�Ѓl�G(�E#���[|A^*d�����r���&�Z�����>w��dg��ĩ�h�ǯ�CéF7�����c�2�n%�|����*���~p�M
�JY)߸�rE[m3	�
M�O��c��
?:��("�ZIY��T����4_'�w��;�M��7h�"L��������ڪ�U�;-�1ъ�ي�H�խa��#�d�H2�h���Ԁ�qz��=[�@k�쓋%���d�4G����&�!uN: �buW�έ���z=V�:0�r8p4�p*, �v�G��2v��hi��Yb�dd�ǯ1�u��}�9�G���H�؉a�-_�-_"��g�iXYհe��ƮF�Θl�w}7�.�=����x�[ +Â-���u����M5���ֵ^u�ưJsH9+"-�[�xkǣؑH��!]-��Z�(������e�sϟ8�����`T]�i��,�_�Ykf�-�,3d�)'�g�@�>��0&�H�����e�����p�&S B����9�$D2wM��L�̂�J-�5���X��A��"��T�������4����,g
3)&�����s�@�Ϫ�ȷX��<�����.:6S
�"�1�(�UֶU@;��ݕnH��w2:�W_�:Y�	gO�rֻf��~���Stq������L��g�7.TZb��+�J�vo��.u�rBf7s��8o�xx�a+����8���*emo+?J�0��S�b|;��j������[9��<����o(�V%�a�pEBk�V�̛l mkt,�&�騌EUUU!������)+��K�{|Y;J1�n�p��2AE�	�{/�EfĎ��w���}�,h�/Ԍ�ުx?n�uދ��~���.G�'���ii�LN=e_��g��[�ꏳ0���ͺ���oPMRt�L���mg8B�;�K��P�8tF-�tn�a�
ܦ�'ǂ֕�SkY\3y��FWx����3���%��/-���"�.�1�ҙ�P�H*���ߠ�����; D���]3�ii"	<֏)iW�/�y�(%'���p��f]�8r�]�
��`�Q����g���y�e�?P�7���(6�HH��CN�,L�Ȉ����e�d[[[š�˖�����V����,��Gj��߳��,�u�����NO�^/��6?�;!��ux�ųl�@�&�VE�EͯW���/�u� ޡܩ�=oB�$�3圎ͼ��-=�KU�����^��/.�77�>�7�eH��3��s%*r�y���2�\���"Χ�0�+��?}ԅ2}h}�� #f&�u��+%�>]��#E��>u΍�gAM=�dJ?/��[�kq�����^�M�r/G�>H6�8�kQq<AB��0av�:���<�WC�F���3�6H�|�)-�%��˥�d�z7&�ҟ��j�ܿ����p�쪣�Ÿ́�ȵ���"�|�\�4f����zI��,��ѣ����3Yז�&�-ߌ��ޡsc5-A���'� NG��=!$&7��) F��K�3��~n�#,DR���t��p���`���n������3�[_g�!]�?A�����J�Ѱ�����w���K9.F=��V�ǓCue3�.ܗ��
 �1~&�V�YM'�n�_i~��N�m9����;�qq�RcV�6���[����|PFFNr������r��d�Xcf{��cu��	�'��E��X���#�K=�|x���q=*���ps�����i"�i�ꪞR֓�I�>��ݗ��M$j;ϝu��v�^��s�K׾y�t�R띪��=.y*JZ/o�Cz{+C��7<Ξ��#�"��>m��_�?�B�|"Ȅ�c��ɩ'tt��wZpy�:��O���fa'U;'��pX��c�q��͔�����L�y��m����h�!N�˝��<=}]��ht4�3N�\W��Lu�v�o͐@������#�H��R��z� �G�����TM@�˕B��7�����G^���K?�_�-��:7�e�&���zg�E�ǹ���f�X�]�.�Ex�2ҷ�#�$��t���H3��()�H�{L� \�l9h�0����Vba�ا3�0Wa�Cn��v�j�r�|�A�yT��sW�TW�tL�<�K�D��V�xt�Q�J��F��F�u����P6�jóxj�xA6|Q�)~�[��rY�qx΋	�.��b��UE�!�46��F�V�21������ZR�~�7�НX����ܘs�q4'd�8���RCo'�H�*H�S���B�q*���ϐ��	�~�_Y� ��g`S%-v��W��H��M��6���ꂼ'���\��n����ݠjnn�O崾~�y�_���6����,�V;w�Y*�_���KC�CB��6�.�ٯR��;�A�\t=�y�\�N3Z�@n碖`�S����>Y3�8C�'ǀ=�];%��� �(w�u!i�ش�T����+����@�I�����񭝘�� �˭im��ժ[�U�٘ۂ}�w���/����y_�*��~������X3�622����Y(ߏ/�����QTT�X8�!���QŒ>M�o�7��y)�~Y�����P~*���D?Z�"�:HD	I3�\=�o;8X�}�<�
��O(�x)��|k	�,�P�;�~����c}��h��廽t�M�|`��B�~2�ȱ��S�؎�̬I%�|�U�{6�{�yf��n1U�p	���^A�ΰ
s���}�B_�w��k��A�hdR��n���ֱ]�܎Di�P�Hi1��B���O�CI�*s�52,�顪��졂j��c��,m��s�$�.��{��2<T��Z^nW�y"�D��}7l
n���F��Q����K���r�'z�HCK�jҺ}� _��P^H�,3��^OV6Cb�7�yua�V`2����q�2�8��zt��k}�o�� L����D�Y���=�}�Z!�7�ʚx�)�#����{�[7e���q�O�2b��J�"H�u]����C6�Ēb�ԪT�����d$JR�S�R3�����^ulF�*�7�����a��䎌��΄�,���ox�Cs*�/,=e���5�k�c"�ƪ��!���kCk��e��!d���zOƏ�;ie��Cts��*���̯2��%�O0��V�S/�P�կ���$~��V{��:Vƪ�'cڇUR������,��x�*��v0�;�eV�ϦA���.jf��{d�����%�Q�2������a�	�fhfv��$F�FD�E��,����%X����io���,�p��J�#ʻt lw���al��\�Mp�Rj�]k�<M}�P�Α����{�aM��g�?�m��l�&I.�'�a2`�<��C�m���Ž:z���'/rQ@�u-�2��)y��������2]Mł�\3�g����C�3��������yE�U�u��aɃ4\�= ˌIl�ۑ��Ҷ�3�n+�j�ǝJZ�����=�AФ�(�77{{�ƨ�X�a���4D�'�W�Mƫ����6���f�;_^��.5A�fK5��Sր;T��*��xM����(�:a��qJ�-�p�=�=j)>n��/��h���>��F�.�i��WU�v����⚰?3r��;�^�ǉm�<|��T��h�%����}7�q"��qq�����N��~$I�t�H��B�,�;ZE���l�.E���Aƴ�}	㿽 �߇��[/6��SUQ��7:��.g��.�lɤ�>z�؝wI��஌��Z��!�6S��ⴠ*���x�
�(��MwH���!��� KK��t-�(���"�� ! %ұ�HHw�"]KI�7���7��<�;�ι�{���sff>$��f��������v@$��վ�W�
�L~N.���И����D���W���+�u����o��+�g�f��85/z��U׫~,��lq�n��r���K�
��U�����	�}��z��9!�f���ұ N��1T��3vv�^�64�4~h�>��1�I�]+�V0�3Xh8Y-r��e{�V=8�Q��U䂛L�t��aZ�{sUٵj3^f��:ф��[�_S�R� ��C������j��љ����=0��!s�7�����sR��ˉ�����[u.M��O�=�a��٠��k���8C�y�
�;�a��m;?B����W�����
��0�4�x��Ѿ�������OO���Ǥ	�Z�>�IN��Z��0��.��#�e�pU�U|o#*�v��G�p�L���ZR���3q��J"�و���M;p�x���@L����Xe�D@���Ŏ��2=וWa����n��P�\Ppq@ȘvƢ�ل2��G3���ނhy5Z���M����l���}d~?��<�M�(ɳ�Q[{��-��$������1 ���kx^�o�zff&�����t��wdVϊq���uz���;fY%ױ�=�E".��_3^1VJ�f��F��G�����ίF��𚋙9β�C������{�4�{��=�d@x@'�ߊ�3ْ,6B;#�x��4�5+�+�C�a��W�2�c�A�� O>}�3V�N[�؎�߽:�3,����#�MᰲV�-��	#ԫ�i�"�g����@�߼I&�O.��E4 ��X�l'�m^�����%�ί<��7/��6[�m�I�U�m�t�ZVG���F�u�7&+¿'��o��cT�9T���s|{
}��)h�"�Z{L����S��� ȥ��!���s�WmNNDAA��I�Y=��o���y���ݷ��|��<O\G�J�Z�+c�6U���q���ĝ�/�,hArF�(����)A�\����(�GԞ��W�I�LMU��q������yy�夽�W�0��)�0	s�f~����禯��]��Ș��b_���S�fҖn�Jb�|0�n���E]����c��et�G�2��46���t�
�[�����K�f/��i(m�)���i�Ǿ��:n����n�v�.�-�)�n�&�9p���F?<��[l�vu��?�g䂜ZU\\�.E.Ռ�_�DB\����bo>R��z�`���܆0WxKl�D��R�aƍ	$�!Ѓ1��KPkH���f��>0YoGG5��3�>~��Ҁ�n��gEY�I�G*j��Ү��]J�ǷZ0�r��so{``��h��wߍ��C��K����s��Ԁ�=��J�`�#
�YN0,:2�x*�J[:'϶7]�\�A$�I*~ ��	Z�v._3���}�i���	)��#�������ck35�SJ�E$p�ŷ�z�7���۬�^����A5�TUUi�qꜬ��u�����i�֒2ə44�AN�5���gb�}�Y�vv8��A<�2��ܼ���4�=(����
��(o�	�����b��"�ӳJX�%���n�@f�=,()�캰8���٦���EARC�Srdg��Q����b����n���ƣ#��x9egg��P�O��|eu�BQ0O����w�و�)s,=�g��{��s6�nh��!�4�O�Sl64���`� I�귛�%�I�_;2�~,�N�����ut�$~E�2H��8Ԙc�a[(���馉TW!���<R��b�VNf�L�����TJ��6��wH�8!��Xn�g��*鸆&��_]��^��E0�q�<�/�C����1>N�-�zb��-��4�P��wwxx0�1vy��+2��-�Q�d2�� _��/7�;�Ȅ�Jgb2��f�弮w�1*��}%��B�K��X-{�uiȟw"OZ	�BG޺
XL����j?dG�W~Q;�J&_����լ?��	k�(�p��wY'��l�'�ı�Ə&�T���S�c�gX.�{�QT�u�ؕs�I�3i�ќ�\�9���x�ʢ�ѻ��<r�^�̸�דy>�zv����N>�����vx�V��6�G;��5I�A���\	�W�2(��lA4�HN z�}[��}GTԸ��إ8�z�g_O�0�>Z�H�d�.MZ_�|Q�d{{u��b�{��Ǿ����,���'�7.{t�J�\0�ػ��; �&	�\Rw��a-�{4T+CXJ��::Z|7d���x6��x���镛gY�0��[����,�j�e�pl�����TC�y�r���١8<_�.DT�>�����8��|DX����{̋�����4k���0����pg��D}��{<�ii��n��"y�s	|?6ƽ҄	�U!~�F���>ʗ�g&R�;DZXz��g�ps<8�=�t�,
6��v����c�t�cb��q�Q�_˦=��d�6��=8��c��l72��{LZ�[������5*��3�戳���;������=�0��鱸7K�[FU�S.�.57EQ��˱���]��n~�vvHɊ_H����}���V��}���/_^�H6������N�t�x*��8;oI%絞�XqJp��C�td1ou�i�!T�H@��Q+s��F�k�j�v�[�A� k���&���y03<y���c��*��+�;)fX�ô4n����,��P�YV�Wy�+�wn�1�2<7"���טC�=�.1Vϲ�30z�;	�������.p�F����TGM��Z���6s'��(�Ďy-�1��.��h�[�V�Y��A(�п��������SA]FBD6�e��o�B�Q?�=��0��	�1
�K���g�@ �v�B(�� EL��%֒��Pw���(��궒���j�E����1��聤�P�������W���t���>�Ñ����D��bZ�����P���Ow�-`Aͩ�Y�T
�/�n|�3��t6e��>Oß�T����I5�r�\�օԎ3nG8<��~6^�ޛ��ˏ�fP��0g�)�0���'q%���?"�1���&T�S�v�W������=\�آ|�=xoD__1m�%��@%�d�҇�L{R�����!�ARA>(ޅ'����?�9t9\E�δ�h��M�3oz��8K֔~y�����G[���ng1��zq�1�#(]Onv����^[��N_����i�"f�/<�z2�%�{^y�h)u����@�R�b_C�0*�U����XK1���՟�7i�˳n�"���+�d� Nw{#��o���qf�F�=�8�y�	R�{���Aj���'�Ȑc�	Z<מ��C]�0�8����l��O��A���:y�&xM���������}����Z�E�	�� >��Ι�R��G�����H,�*�2�\oF��T(O�sX�V�G_gl���Vt�Ȍ%BoTf�t�W��R�wp����{�>[���^O���e��p	�`���,=7c�>"�d	O"e�ePh�R�|��x�Y�q�\�hǬ~�Q��3'����sQ���k�����	�G0R�)"T���
I-`�׸�z(o��g� Dm�1�3�#~�M������ZR$ K2q��A*��~(���L�a��wEHL�m<��2$�K�����/b���2qo."x(ē�_�-���m�`��@�/�gX8SK>�@D�Z�2��c?� 9A��Q�5��_^b��\k(�p;>~v �ɗ��*����3Ɇ��;�U�!��~��ȅ�}퐓�Aݼ���g�ɷ,��������L�%C�8RY�p�z�I���.&X.�پu |��f�
��i9Z�O�_reܹۇ<:S�w��~ׯEW��,��A �]=N�t<�vQ����Ј�lf�g���"�l^��a�aۻ5�`jm�	�D8D���E\D೭�wW@{���5糛,��<�u:�-b˸�����;TdL��	F.{Ɍ��b|.��٬�i#<y��Un���3�N\"o�}��c ^XQ�N줻����R<o��1,S<���y}X�8����Q(�V���IB2�0J&~x���{��ӥ��.����M��k1�M��iͻ���_0�ޥ�Ţ�����'�!����[X"@��|�oL#�a,��e��I-�X)j��V1L:������
ŜeP*�C`�o�kr�I
��Xˤ��<��EI�IW�V
{}���_�B�m��H��HC����^dWzu�G��
k�u��"B����T��/]'d幠�ÈT�:����r�[���g\��`�GM��(�xV�1n�����(�9�W(�c��w�E�?�d �
�8Z@P`o��Ǫ�J���r�P��AF����=e�E
�WW�W{?�M9d?��$9<�Yc֖^�y���F6V?uzfƤ�N?L0��� ��(�p�I�)�%=>����[Mi�7���!���>"��,{���|�rgQ���4�o�9ɾ�|]w��7��T5�f?��<�l��]!�������:0P�/S�$���P��W��a�[t]����n?�՗���;`-ӈ��-==]f魘��~��Ѩ�Jg�f7���}��4� &�7���"������Lԟ*�����Y���@�&��׊��#P+p�<���ܕty>_}��MR-f�/eO9(�Y�~Օ�خ�'��3���JDv�Nw��]6d	���M�_g��Y�m���k
q� ��3"�5���P����lf��l1�9lsvo��~5����#!(������2���ŭ��`��7D��� `~����>�<|7�Ω� ��z@&���El
�^L,�٥��K�_"���d�l�`�7#䑒������º�C��B����Ϲ�����2�}��#��a}9�6j�ɥx�pJ�څ2g��h����A���Z��AIH�U9���^{����edd�5��S3?v}0G��3��C�O����E��)yN�����5!�rζ�F8����A�� ��K�c/F��0�=���#Yi����@�~�J\���m�W�T���ꗡ�&���;Gt֚�ٓd�s�-�ؤk��G1���>b��t�ߍ�ͯ_�+mT׹��3�3d�5d;�S-�e	K��zM��(ed�j�]�v������i{�׮����#�6k&[�1S;=�q��T���8��0E�.�!WkN��N���������c�C_Ԫv[.��u%JKK��7׀��X~[l#W�`��f�`tt��m���������1�p�T���ɱn�>�[�>���!���{�j�BCf%��KBq�_wjZ��FG
� >��2x��M�{���.�v!�}���BX�����P`�Ӏ7hAT#����4E��}��ɟh/�����3�5K4K�v�*�w4��C�&9�{)�X	�0�ލ���7���,t�	��wYRUv���R�����	���;w *�jK%jYjH�+�����5�����s�B�fԪ�OX����VR-7Oa�tI�w���f�\�Gw�}����6�H�C h���vv^;�t�c���:�]�����碦��d��M�s�:�{\Y�l�>wz)7�D�;��U�����[.P�g+zN���[D�$_>�g�q�*��������c�#��_�s����@��7�G
�̡Е�wir~���t�e�0����Y|�Y��چVW@�<3B���?)��ᤧV������Dԋ��&��"�Y����r���85�W?9(w&nv ����� fO����	����<Z�
��L�X��IK;�P��m_��Yu,�d��G谛�<��E��~�����?�q���]ܬ���*5x�Ir��dpNI���>� Y0˰������c�p.\���*����n����Z������D���+1:i+6���;b�"g�|��#g����s鱤��s=��l����1U�W��CS�C�B�g�?ԇ$ԋz5�X�%.ƥ[>���&�����|��_��ʱ���z�w[
;+�R:NN8�wLjzzz������3�����k�b���L�E���-���}�v�F�Z�B��?A*���d�C��)�Nf�Z7���7b����T}��~:�|>��:�BN
�ϵ��lX�H�=W�J}X��줮V���)D){�ъ����!�.õ���R�b�,�7�ѣL��T�]���{N��Hx�_���"��Y�.�Q��^~����g+
ݏc�kͱ�X���y
�.]�)�����j��
��KM;y
3�MMM׹��lS~��o�@�|�A���������C�[���z���,J�3%=��D�PL����=U��	פD?*�ٻWD��2�:����8_���9̈́�䨌(8���Z���I�%ZS"o0�^�3_VJ�iH����g�ZW�;����3E,ԄHm�ˉF�,��9�����D\?G�kh�����������O#��C��Ҭ9�׺ߦv�
L�(`���`gg�ucl�Q]��aM�J��t����I��v��K�t��vb��0�7\�0��:հ���:����TĊ'=*f�r����~?x�֓*�6��Ĭ�s#��Ǧ�p�]���#��",d��"��o͗.`S����њ<I?c�W�#|_,�5�������y&b�0S��I�'����Zw��	j���E��!�wzy(�c��,�S���QQ�:�Hs,�ɝ���u��a���i���|`��,���F�J�"��Ѱ��Ϛ ��g��Ok���P"��s$����D e�::$���ʟ�8�|��ϧ���8�!�yo۰r��}��tQd�8��<��Z�}��(X�/ԄAL�J;�C�dvP�����Q4���P�!W�:�l�T_B>MB
��xI�~Qډ��<u�f}�1��dw9���#�)c�T�\�l�̻�Ǩ������>Y�C5쪈 e�$}!ʃ�����/����;�k�[�U��'\5Sǝ�a+~�wߡ�#��g������𘵬���!ƶ����O?#��<��0װ݉�0�vS'&M���V��d��`v�{��*�"�1���Ўxr1Z����dq.�F��9�qO��i��3�IY�`CCj���6F5��0@�g�/����Ѐ3R)Tϝ��Z�p��`��!��Q�0q���h~te�������q��W=s�K�B�}�W��b�]��o��{�sPr\������o�.�*�W��M;�����rpp�w~mT�4�%��@���GD3;VHN�)�]�����p�0��_�J�z#/3鞖�T�O�"���߇�=ۗ���1��|��.�Q�0���(b.����#�ou����B��%�NnH/HʜR��-ij�+�f�rȨ5s���c��ߺ`7�L�%JK7},�;g����,-���gM1���k�9�/�Pk^�T�	S���	�y�_Y��M���qp�<e�/���$�J;Q��qa��C�!V�r��Ώ ���>N��5�����1�WkF�f̓��s'G�̻EӍ���Ni\f��7G=#������X���L%ໆ~V.>UF�:hd���Fl�Jʡ�3�=A	��ʨ�yp#��o�N}�j5nzn7F[��R_#�Ř{]�"Aly�f�_�r�V��㽷�E��Uwp�������ُ�� ¬ ���a+�뒙btv6�=>Pg�_j��gǲn-+�y�5�&��f�v�=�"�N�Ǣ�?��� �n�:oY�"�Aw��߼!V���v�N�]G>1�g��J�*P�'<d0�j�-j�ᛩۛ�T�6���Jӝ�c��!-�4��>�(}kU2�=G�T�{��z�pat\�x�o�Ҕg���fxjʤ�Q�����嵂/_�h9r8��q��V�����R���4�~�2��	Y��ؚv.')�p<zE -�5e1A��sc�6#q��j������sI�� �ez���?.�?�o��h��J@�_�:P�~k����{�e㋹v��N�Sg��l��Rk����7c��)���!@�{q�m�8���/]o�1̆�U�X�;��ƙ�G�1 e�ļ
���A��=�����Caؼ��5����j'��DzR���Aa�H��e�(�Un��)�쿈�
�s�(��.\�hg��#���dS\�Iǹ�8�O|%q�$ �-�w�"q�|��^�̚�@�M���Ml�鯞5��[^���K#wXF 2e�{�Zb36\�qZ����l��-�����m]x�R-����.�Y�����^��|��4;�9T��u(ő�QΗ�?�����O�5��tuuEgT��1�1�c� r����!��	6�wq�-����k�,�3������ >g�o]$�F�.������xŚ�ċ�*7��>K�Wz^=� 򉦇6\�Y&����D?C���%��H��_�npl����T��]� ��1��`� �:i)h�t�鳰����V�[��G
�x�=R�r���3��FG�8�O���Xs����%..���SXc��xmK�K ��;u�
�|urF`x"�um�֐[kn*�$2d��"��-ܙX��\�Y\�_���Ҷ�`f�z��ɋ��Qy�G�Wb�w�]�&��S��c�7�JL��K;�=U�&j��qP��w>� l?�?��C�/���=,��i��kj�¹ݳ��nM��E�L����.���"�K���%�^����y"�6�.N߯!�2����fTՌ���wQc7zr�5�2+B��Zn������z���/Y�!���2[�ˀ!;5=��
K�9���,Qgra-K��6�dRa�����p��2��|�\�k����o�a��ȸ�2��{����wy���A�U� ����(�͒�J���I�f�:��b/#�Z3��a�7��2u����� a��:����=Y7y�s͋�ꉭ�]/���'OH�+/ �9uk�%�~�҉����5�����I�A�I=�f=�W��|��r����r��y5��HY+(��fY�2�ò��qc�X�_.$s��&o/���b-:�/xڑ�oZ)yt,Hh�h�
5[K��^�F?oCz�Jq�e���2��W�ŭ��
�V�g�P31� �7���2Y���#	.~O5���E��i��U��^NT9�RS��pa�ɚ������|Fe�gk�k��KN#��z3A�n��"�t@�<>P�b(0���|�o����ck�=�]CYwJ � `M�[���j����C���`�=J�!���okz��M��[�H�ҨSb�P����s��`DB�Rݥ.��zs�+1(�N��>r�����b�s�KJ҉�߲�
(�޹��3hC���Aً��J\;A~�|�e(�&�.U1#���������-'i�c�<�����R���f�q�9�/.����,Er�2�r[uST#��HR����P��X5wT1���*^��E�F6@ݜ˛�%!4��u�p�Z���$!��7�^�u���\=!�'���w`����7$�����������
��6gJ;r	��L���":���֠��Y��A&Mjl��N�#�^�U��+EǢ�hR�?���^��+U���%�i�\��x�l:���{;�|>��MӏT.���?�&�G�C�Z�	%l;H�/�r�� <��3��^�]aڅ#�Ƈ���7�k|fXBIU�
��}�֑ϻإ��g�ݴ�����B�~U�B%z������F6R�?@T.�:`b|)�ޤ�K�>�T5H�R@��K��
U��yAy�7�U����T��Xyt�nz��ۢ8 ��{��Kw�ƚ'����~˷���U>(v�v�c'頋��De������D9�ӟR�0�YBa�w�f4�А��7j��I�wq�Qe��#D�A�ޟ�<v��N/�/��8i}:aV2��`��F�%�sI��׃�c��&�8�Y0�^b�/�M�C����?t_���XWC�!��؄��	�rZ�X�n�`�+G�=�y$>T~ׂ�L�_���8o��Y-�!� ��LCAяf�ďǄ�X���4gh3�	3��I���<9s|�o�w~ޓ��[%m�ߖ��� рf�w�߇\��d�׆I_L���#�om�tT��*���;�k�K�V������s$�SBR[� ��� l��$T����E�#��h~��Ǖ݃�nG=tH0'�A�!�'~����>�D���c��@C�4��o���z���y�mP��!Q��q�LՅ� ��M�m}/>1
W�ͼ�{�r�`P��km�c�P<����DSf�۸���wx93�f���x�G�YNM�\�{���d�w<��n���F�+��a8`�Ba��=g�w�����6�����*-�-�	,��2Zu�?FT"D������E!@�n�*=��BZO�_��^ ���e+P�].Yp�^���8����d�D{A�B�8X��I�n;Y+�
Z7����S���� ��R4�ӗ5�Vר �|#��&F�~Rkxp�6!�iO��|��Q��$��.��@��� � J	N��p��m�R+�'goV��
�U0a�&ΪkÜ�g��wԳ�crAu'�%ַ`��n�f�y&���w�o�KFVV���zeHU+�2��ȈΓydj
,����9d������	W� ^�>��0h��7��8-��E<C&,�}��^����}�a`v?����4�傺FF����DK�e�okJa�6;���R� ���cvc��g'��D�q3��O��N�~z�O�&����KC� � ����/Z`�UO>M?�\�U���:S$�% V�zA�2K*َ���U�!�[�����È],Ż�-l�"j�T���������,��9��1wMg���p.�=X�8�t���m[�!��#O��d���$T��6-����X*u��3v�&��5%g���$U�>j
���-<�1�='�G��!�_�R���2�)f7���,���K��]X`ƛ��)
���6]��/�j
�I��ra�S�F��(�mV�V�j牄��w�����D��L����&��a��d������?��j7f�H�}7X�X
��F�/M�ISbT��t�_�.S�=��	��]�� �:̝��k����D5SK��8H�E� �ܷ���C���7��e���k�Lg���nძ�r������ �翺<�Ҿ�	�w���n�%m�@J�h%� �a�aD�������/��P��#�6-��!�0֋�%�/��Ԫ��&������-x/��Pz�w���NM����"!�®k��n�3d�MoRz,W�:��l�ڣ)g�U�E8U�~P�g�i{6a|�
�
�
�����ḟDg��&HL+jk�o�)�E�o�LBvt
G���#��@������g�n��.�7���7��)q���+�ґz><1���M���.�ή�CR��mD�@�V}x ��w�вs4����\��}�^���r��R���}�u�G�7,����`�*��݉�@��a T�)��Ɋ1O��Mb߭C4�3��K &>�������>eѣ"�ؚ��bAȮ�۬��Z�hd���)��h�@2�$���*L��Զ��"��ŒݔKP��ް
�ˆ���v���f!���ڼ*do����t�^h�F��O$���T�%ʅo���Z��-y�Be����;y�g��Q�1���B���
�맄�9�4bv�Y$n��#W)Wb��#u%}U����^,���q�'ake*�\���X޿��RI�#B�|u��l��	�D�\y�\:��n���8{?ꖊi��Sea�m�/��m��t�'.#�x*��|�ӵ��N]j���KB֍�h#[�
B唖����d	\���xr��UhD�C_�2�4��ϱԳK�x��#�����Qex��_�_^�	x���)�I����te<YS��h|��cU;��x�`y>��U��1��]cS��@����!j̞8 �Xz�7E�B��S;�E̕	�T��S��ӱd�Ow��0�����8Yx
D�O�_���\�zy����x��G��QuyȻ�����:�{���{��b:�`���m�'�#� �=�j��8?� �Aj"���@�|{��}�H���-�,���߶�/9s��S�rn'��x�a��-��ѧQ���2*���?m�jܩa>�4TE�N$�j�Q��H��&&�<�Βh�*de'2�[�K��K奄����I�T��6zt2Eݿ&�L�b�j.a%��	����?Y���ｾ݉&���YHKS.����S��-¸X���X�� ���:��_V	�|�2�n-�LU�t-/}����ni�-M�����v�CKl<�*����K�C"���ڶ_or�������a9�����uF��<��<䄃s�ƕ�[A~):c��)��F�w!qo�w���3dt=���,w^��i���O��\I�=�׷�D�>�4WSS['�v�A�E�Қm �iϝ�P ���D�v�6�X�t|HۿqP?��v�O�nҡ�Id@Ybj�<�������*W�{�F�VY~G�G>��f��nu�уNsC����b`��q�K�FP.^.�.�&��&�����῾f��lr��n�!��w�k�fZX��$�x|Eԗ��4�9 !�R<8�	��%�_M2F�f�{INn0�]~s�-�yp���d��D����W�&ś��v��y���c@�X���������A3�3�����Za���!<��n�''�m��8lk�t�'�~��|�n�W�#�����rIO-�=샫�M���m�ua�~G2-��K �F�\�Z�=���+B�na�|"ڥ�W"i�5A���w���{�	�!��x9��7����!ǌ,W �����b/��`�$�=���2,��%?f/M	0,�.��Ƶ��:TÖ�D�|����.\�i�/٦�h�e1��/q��)�+^�@�˻ف�E�kr�ߪ�s���g��%�l�~3��ltJ[���=_*���=ǖ����F�:Lߓv6��3�j�w���S:� "����1�w�4ʾ.�촿1�q���)Է���6�=�Bly�%f�k�����"#��R}��vku�Պ	���tb�)���]zRҳas��U�m�� 8sp��^��%��� &�N�z3��lk��c?����P�����)����c2�5�.S�#���Ώ�7��� �Ct�P�ac8���n�<G_̬������I~hy(g1�0o�V���w�d�+lv�o���c���E����ʦ�L���W�3f��O���Uė2�l��skh���\���(_�Q̞��Q~Q�=���s��Vc��UGl��J�����E�4�Y�i�2�w'�˂���V���9~����f�t! ���~�h:t�9nJ��5"@n �k>Yy�9o��.0���8޺�&�;\� �-O�Y.%߬�͸�˰�$��]�l}��kZ�q�A�M	&9�ּ��ۡ\cW��#8M�bO�BÃ�|�1���&v0��}�9��#3�=g-�j+b92 �\/jy�Z�FrR�AU���)-M��쎏E��ڠn�{��4	q�D��8Ɖ�g�Љn��Di�Y���k�_�EM��_�#��ѢV}������v10R��R�����0��l=��r��8��>y�hg�K"/������@Z����;�e�/�s��>�:��쎠��i_َL��G^<��?��2��q���0�ܤ�>��P2HH~�t��0`��@�v��ybS�Tx�:��^l�CV=��e�j�������b1��b� �b�0���d�_:ˈ@J���1>:�����÷����j
�nR�&;�8��˛����g����o9��y�	��UVS�]kXظv�z��c~�2�n��W%�Q��c���nh�R���/q�v>��+;Y� ��i�NH�&wD�'�� �QLt��R�R�/��~M"���?��W��gdJnf��g�-ƣґo�fR�ܙ�.���i�l�+	]�`/I�<L�6��X�x�Tֈ�)o>&�o�d�7J_�.�mY�0��s��c��U��9-Id�pی���頛��c��)�[�W���}d����i��e��j�~�'����6��U�'�o��d���ln7���}�ce���d�����k�>�T?Y��%%ulh�=Y1��4�rb��/^1�7E�-%(f%�(�@�Ʀ���e��ަ@x���ժ�齬��_��B��U]��TY�5>�Bʂ�Pe�r��GG�ѓg7d�G
B����+�Y�~�����@XE3CO=1j@���XC���bn��d�{�[��Tޅv}cx���e4�$hf2$��4%r�]?`�yiッ`kQ��|��?�T�ѳ�һ��o��D���;�Af>�-=6ַＧ�!?)(�����1ʹ�:�*�f��Ǜb�ҝ"XS���Q"���T5�<mRU� �V�ٳ�Oҡ/h.�kܰ��d����\�����B��f~;]}yR���U����r�Z�|^����/��o:���i׼J��+����]�ˍ�A��ɠ���m\ \C����zI�9׸0|ҲW�ɡxF};��ۃ&��1L([5�u���ae����2"���M��G�������J|Ҋ�a	�M��hj����sA�>����>�M��4�r�Z'��ř٩��ʚ�#�����&f�a�Rf'��kYB0޽#�"g���4~��EM��Z�TҴ�+����{�<���y.zy�	��|"��Lժ=����5�0��"��+#���U��Iv������?{�죄3m'ȏ�=�0�����Z����:��ck�����pR?�?�*[Ћ�4��LEn=�u��(Y����n��M|�]�P�E6-Zu3�������?]��?7����0����	�*�_C����Ԥ�Q�Ը��s�M���ï����"(5�E����^.V�ǥuL�a/%?�װyn��NԒ^O�)iߏ�OZ*���*�ye��\6�˛���
�{)Ԙ���y�RF�Ѻֿ�˵v�1�ч:��=I<'�0W6�rr"���O�й��O�,�Ŧ��-�H]���Zg=���t1^W�v4:4�hŕ?�b�Y�H�cf߮��É����/�F	�#����-h�jk�*��3���i�^.��P�����Q�1��Q��ժ������.'ȶq5B@�r��d��H�*3��#O�'�F-�o�&�xծFb����o*O��6�E3�4d?�j�
��Q�a����j�u�[����h�c/����;^��N+hFxI0���0��c�����CxYN�7v�'��S�!%N��Cx���o6��okuv<��s��
�W�3J#O*��/R�\����Z.�Y�;�|N�4��gk�s��AsǛ��� ���u�J�?�����,)����";ށ�ct?�{�ZOx�V�2���27�ds�x��=������l_�簑��DϝdQ�����b��Xn|�+��}�:�ϵ���+��n���h�Y�6��}�P�v�F�K�`�V=���诒�\lK��mys�2"A�����BJ�����p8�t��S��ܥ��������r��o��:��w�i9�xi<�E��2��b����J��0��������@^�s���ϔ��6xW\\2��Qі5?������F1��
��}�{���s�w�bhh1&�?xQ���U�T�X�����:."����:O�������O]JG9I�Ҡ tඑ؋��Y�4�xH�����	��QS�i
��A	��^������~}�֜�&(����Tc�Q��I�8�������q�J"�4�4��&�wY?H=��1��>���\�wX��&ȼ �HJ�'�|/��\�9��+L��8�N���nӱ3��G����cI9w2v�d��0wh�RhWw��	~�4�/��}�*���n81�㍘��?
/�j��S�#̈���o7\^��@=�#���|����1 bc�64\��j�Tzs��7OѰ�{���������PPа|����Ga�� (D���M>��b����U�ڟ������������7FV�C��.���u��ZѤ�q���~un1�0Y��?�u$�0��N�zY�C����1�"���$ȫ#$�mɰ$
	RR�;�<Owj��t����>x jii���=R4���O���!+^���)]+�;��D�7�z�NNDTT�ñ�8�SSS�`�R��M����gk2vN��n�����_6V�{Nbg6�DA"�Ş�rcMcJ�~���ܙq�1�=B��B�h����4�!�=�:c;#R����R��k��\��=��#p�e���@��Uo��ƦGW�Y{	hg��X����w�	N�
c|	f�d"��-��^2#;�5p|�(l�k�f��Oߏ�W{?I���-����|�� �� �C��8|ZF�,��v��*F+?2|���iK��=�ڔr)!~C�@1/�&�o���o۳���F�%R�~?_+��Bu8l�a�a�b"1?on� ����1�;z�!��
��Q��
�)��i�H�$L+�42<�?zB-��(�qz�ys����?;������.z��~���ֱ�m���
e�H%��ӿ3����x�N\�nހ��y�'W��'�����s1	����R���y���ɸ�yE���j=y"�Rط��)zT�4����j>�S�+���aQ﹄���L��h��.R�;����gy2�
��n��>q$�%�V�s�XE8<�N�m����>�QR_���ò����	�/&U�ML�w���G
�o���Y5������ q�q`�u��ߦ-���'�\���O��BCcd@�:;��xW�I�:������R�u��)�����Z��u��ҋ�ņ�G�[FU�u�� *)� �!�Ҡ�t#Hww7*��4(!���!�-ݝ�}���������=���3c��֜�{�:�>����x���q����鑌�k��h�J��X�����=B�dћ7/)sm'r|{�i�gIŃY���_��'���R�fk�
�.�����w��?RPR���bz\�**F�/�����f�]��dD�F�}��Z���b�c���%�<rR����{�H;'���<�ܠuo�Lx�9((D3M�i|��*a8+M�P�J��
���zR)YY�=V���b$"��ήא�4���L&Ά�C\��f��Xm햃��ޞ��<^���<o�K����I��r�\�NC֤��a�7�0�I�_? H�r�/U ��m�P]�.R�� &�@Ģz���9�1�����0g�8�b�>@:�q"��k%���0������Q>��4����'��^n_9��|A��@TB����
��_D`ba���ో\���-�n��ڐ5���',�cXJ�'�Ϛ�`2aĽ�`ko���w"�qD �/��kRH�n�R	?�HW���Wd+�h�qZ�3�察�@�,��^I��J���;�l��bLu��qRSzr�'�*��z��?�>���+ ����젳c�;�����P$���'q�G��J�"�T^>�aw����)	����OkPz��G��c�a�0)�tVZ*E��X�ВuT���H6��X$�|B�L��מLT���WA_�߬�t������h�~�ЃH��쏸Vx��i��<��*��_	�w
(�ӗ2�%����f��^�Lu��e��L1�Ϳ����K)NwM�wB���up%.)ٞ�����7�jc=�u��K	��!�/�a��35��tے��d��ҵX��U��B���yY������(#����J����zK3�?X���~�ml�j9�b꧿ۣ��:���T9"����������� ����H�ǣmG��R�O���_=�u=��&z7��e��8��b#�
�\:�# ��Z�]v̕Ԗ�F˽�,��{rJ���՞vyPG���s����2���]ok�<�fVQ�aM�=Q�5j?����[�z��:f.]a<�l��|���Ɠo��(�ڍx�{#���/����:o�k2����;�&'��I'wa��@K�۸PT�Q�������W��|���O������ 6��8��G�=�D! ��w	�����������1x��S�2������\�� �mru���^щHV���Ȉ��Q�oH��ԃ��7�m�f��t|eȊ+C�)3������?x��	�Jd$�c�����D�t�!��$��'O���_B�o�e�����s�Ǝ���c^^��ps��=���!�����Waԥ���<��9v�^����"��96�!����#:::�Ma>66�ü�R\^�xzꘙ�E�Ɔegg'.%Mo�/��ttt<�Dn^ޫ¢"X���8f668
jjr::��$$���0�88�/��Ao}�Pz
<�r��������oA�d<�w�j��479����r�G���"����qu��D���Q��ɿ-�Nd�U+�/��]n����@MM����:8(�yUQQ����������a]���=2&�bE���D(X8M��d,m�V�k��grrr���m�XOBA#�K�p~~~$����߂=~�����)�IJNO ?��a�U�� ���bsBgcO_c=����*��b	��u��N�zX{{��ΰ�L	,v������_y�())����!��v�#��n�R�|�$��'x��@M*�h�_^_�KDS���&�e�JYpss# #{|7@?������� ��,�!o*�������t�'�L�E ��%�D�j<O�Pdt��wN���D6.�5������3�N3��l�}h�H�J���3{�*P�?~�z�'h�x��\��g1m444,mn�

B���:\�|dff��qN�J,�����s�C����2SJŉ�;���#N�������⡐�kp�
D#�$i��~�<��[\#����/i?�v�M�R�~WP���g��L#����<��K���D�]�E������4y��/��5$�I[�p���'�:29��I<s��aL�M��eY[�����N�7�z�r���U0����f/%�����Χ �ޕh7�\��d�708��i��
'��e������*����Ơ#�t"��!��}��Ze���<�US��cݽ�Q��#Z!�%/Y�_��#[XX䵳�^̷���	:�f�����p�!���R�-�����M�H0�b��#�0|N���N�����N@����[�͂h��<N;��#=��m���K���	x�C����^!����)�4yy3=��E��-]��rۓ��EFd�+�����;j�Vuml�����j���B�ޙatt4u�K?FB䟆%�0��O[3%����_9q�IIJ
9;�~�����#�7Tэ�6 G���^	�K�ˣ�1j���\g)J�����Y|,jY�"~]ssZ�PO���$	%���a`,,vk.t�ў����گKޞ������$]|R�����m��� #
!�s6��7WֳP�a�~�
�7H������,(8���&�����o��&''m�����������F������{/���񔎮@��m`���dc��`�>���LeEH� iF�D�M9B��C��:-V!cg�ʯ/8xCyʴ����s�𴍌`dI�~��o������ X��\���Ǖ5�0u|�8�������XXX(/�a*L���N�����4Y���THX/��W����/EȂ|�σ�Ӎ����Fu`�wq;l�.6y
����nnnz��W[�e�ʴ|�G$���a�hh��YY��㹟� ��@&����FuD�����b,z]���R�v���Eɢ{�s���s��ҩ2�V���0�Yk���
�2h%��r�b0@���Nә�W�^^�{{��,���/@[��B���Q�`4��������L񍏊�L�ZLBC� С`��c2⃃��LD��H���x��}]C����x��ˢ�
�'$�~P'�[�u,�K�l�WD�r)((�~�x�OU[[+���_��(  "}fv6��ӖOpB�*��>���U}QK� tys����O�����Ϥ��1�L�n>.���yk@��Un1U�F����Mv���DDL��� L�1���n��T�A�����yHw_&@���B&��LS�:*����������/G.�����\��|��	//o�ar�������^�
�OHHz����0]e?\c����#�ǃ)�}�{�?k=m�A_(�_г���s����� D�o����N;ʤ��u������� k�䛽�z?�P���ߋ\��,��*!!p�Ar������������������<����:�]�g�n�����ӋG���8?��⧦~7]��j��ߖ�ݯ>�����0�>���}y�^��֩�x�Ev!�˫+D�W���Ă����n�����il`@^�V&�����}___���O@D-��Y�Ҫ`b3j�����'C���.y:ł�����W^Zڂ�����G��H#�h���`ʬ�y\��N�N��[z{	&�o����2s�
��ò���ǊK���n�~���O"x��8��ڌ}�8�BP���x��ӫ��ѣ�)P�w0����΋�.b��T�kDFF����?�R{3UP� ���6����V��~7Q���e\6k�1��od�����%�4yf��I�$z�J�����Gk��ի-�1��~H�3���
D]�h
A4u6���q�
O�;�-c���+���q��Z��Ϲ��zc�>:�`��W�g�2$X.-��I!��LJHʶ������ �(�/LX_q9Y�!���@ ��T
ާ���@Ȩ���>$#"��53��g�O�'999�44��_~��ZP@��^�?M��fj[ĽR�'����+�n̟jx8_$n?�?���<�>���=Q:��!��� �����n�6]����8��ׇ�����#����_D!�5z� ��r��z�5^������!%++��=vTt���%�6�o1��O tWݏ�ȑSS�t���mO�����n��Dl9,�9�/�<�Y��d��i��.7"����# �\�2E�����i��Ĵ����(,��hw��q��58(X�c��.(D⣤������9f�[W�>AΧ&x2:w�>h���i��X�����-&�\�LI���u��^���،lx���A����T���7�I�\���9S^qAG�2�7^ ���=3��p[��<�T*�o~���b[t��� s�ˍ�H�n��0"[���=�����c3���K�<�=yے%-�A˂9k>���15�����
�<�۟�(�쓲���i�^ ���Q+o�*����I�@e V�<����	����ɝ-%���_`�p`�����>�5���k�rq��:�%q��nDm�����r���p>\�w9��7y��H�_N�N�hqq�����,8��t����z��:�$���j�!�db],���|����ǝ�����[*�jf::x�Ԯ��1.>w_`֡ߎСM���-�&��a�*���������핃�&��X��׽���/\r���S����G6�%$ZEp.�02�V�������B�Ụ�U���/5��hi�e+x�{�v�\��+�ff�����~
Fc�r!x�2�&�}&	8Tϓ�\���Q�% q����Wm#���N�9H*���$�����1Q@w����r� AǠ�I)��1��u�l>NS��O9� ����	aq�\�fP� �m\��:n�� ֢��T8�37�:�4�y��o=}�c�%x��[���9�羇U��6�`���eͫ�����v�o=>�!Z]�5I�\���@����fb~VZG2��߾��kw��0��.p�&/��$K	��dfz#ktJJ8�h#��f1�
����kd�HݘGĤ�cٞ�ϡx�_���I=P�RiK�v.�YP
	i9l�7͢�ANFvU<�1��X�����D D�8��]�/�Z)����([r*��@l�I�b3i���
y���p���eJ�����b ߛ.W���+�Ok�o�v�4j6�L�' C�յ6�̤B����\�0�n��n��8�7��<Ql��B�94��_X3f��!�WUVJ�5�lY�����C͒-�������f��#8�c�NN�<�<��M���Q��ڃ0�E��@�&�0��OifgS���5�fX�$��5[��idlL�N���dgdѦ��y��p���R�2�YPM�;tq	�dQ�ˍ�ֺ#�,����|	P`4�������32zbbbR��g�V�s�BF'o����'p��[�^ވ���@�!�ܝ��r�E����LJ"@�e}�8�SP&���F5������. J�'2�~�����.��=ۙX^]�շ��X0����v�X��݅A>��h9=��@�W��^�*-/w�����t;���/h��Ԩ�qɝ���q4��i�k��`�h�E=*���Q����H��'��z�o�ؽ8�m�PW����b����J4����%��y��ġ����p ���~��f]�]a��A��[k�ې�n	a����JJ�r�������b����@��>0�.���pw���NSF�犞��S$1"(�}���x��,Is����`��V��[@"#'د�"  @0���~�c��0��K|W�s�$����v��
*C_"^tEg8���G�ȧ�����ζ����L:Sm<F�k�,�4���
�TQeϺ�zrzz�}頣#[�d�7����Ěح�^"c�w��y���D�v�[^(��%xH �"p�j> B����6�.%���s�"��ᰘ�n�IgF0�
�4)qCc�Y��_��l�X���pp�	�r��̖N�\�t-��ʤ��r{uR����!α\xL�ciU�I8�
E�H���{%͆?���h��?i]; �0���*�#utt�p9\�rډYp������k	��#СS�Z��Γ�ЀS�p��bJ+�2�N��`',.>�,��9�1j6�-I�D���"�?���䥵�Li�QИ��$C�&P�@�x����T�� �jeLNp"O�mG�׍s|..������g��R�e! )R�����D������ɓ.휋��&��kk����K�\yd�	@È�$�'\ 9n�K}K���r0�'%��n��ZWץ��I� �¢"����Ix *a�3�צ��>�9���\1���i��Yl�.3\�ň<���/�0htop�e���<�s���#�7q(4�?�A�e�c�[/�oc�����]s?��ѻ��CQ��Ȉ��d)�&�10�N��¸šW�W�WR�F���@sc`!���t������t�Y;�@L�����h}�w�����'E�'m����\���% ���������5��\Ek� q��Ǝ��}S���3Q�`�Q2���T�->W�8���,�}�������3���L��E�P�����L��� j�a����8���53��f$�a>>|U�f0����Z6�+r��A��=h![��
 K�u�&OhO���Vr�X����啕?�6=Q��Ś����ݏ����g㍻1�����C_�\��uXW�U �`[3d�����w�t7%�i5�-¡�[���M��|�3D��K9����3ӵv�b�=?ľ}�>�4�}���xy&[���25���s_7��(0SE�߻9����9^����,��p�³��%�C��w�<D���E����z����t��XQ����ri��>@J�;^�Е|��?"(\�����'n��iJJ�%RQQ�.f��!	� ��{e~��O�}ڷ""+'��=����v'��,������K�����A�3.�����L�:gjP� �#�]p0 c�?T�~���	]���2��N����̯J�1H�%G��:o͟��cC'��L���R|�ҍ�l��y�L�,��"hZ1`��h\��seF%@᭿�輿	@t!7��'�u^���4l��ҟ���r��>gB-Q�)�a~�`q'�MD��iȺ���F�fX�@ I��ݯ����ըa0{ʚ�_����K�m�0�d	10֭ �/�.6z�V��.]���Xkd)��5����۷o%@}��0)@+O@���E=A���*���QZ
V�#&���޸11�^)���Op��=Q<C���_5�#�|i��Qc�R�]��XD���t� �]�����U0�Tq�ҝ��Y���K����3�e��㇗�	G�ޚ�A�<���i�WPPxɬ��r
���B
�s[�lU𵆗	ld�r٭<`�5���x.0>��<�(�Zd�2�zp3�1#��,�/���O�^��O��NL��<����4�*N^�և�X���f�Ƞ\.`J�@�N\��&�;|�q�)�6��L�t� ��S�a�'zJ}:Fe�P�����)�P^���,9�:��6e�C���̡�S����%�jj]��'�ʅ_��y]'j R���Ϥ3x�	>���Jd�#d���6��������Ƞ=���:yx�W���~�����N����%H�eo[az���N��Sɜ�{��+��O&1�;�ư������>�?n���	��p�V��Ȟ���w�NE�*y��lp�z�G���<��s���	G�c�
��K9���䩢�׻tE����È�v�8(z�@v��&u�ZV-�|����!  i(!������j� ƭ��������4EP����i|���ل���6?D(-��� �K��`�}������o�p��V���\g���lJ�������7y��6�^ �׶q��Oq�V��W�:g��Z��W�e[�F?�TX�?22�l|&-�Q鞋���+�̣������J![
���<W捡鋍�q Ɩ;���'0���h�uQ'wL��&j�H�7GJ �[t۫���F&		�'h���bK]�>~uuu����>D�<�o����1FnV#�������3_� Ɉh��	��T���F^0\U�|eDN빏��*ł>A?�C���&�]l��%W]�nv�{-S�Z]ߑ�����9Xl��,{�	޼����M8M�a�1,�������$Ôl�֖i���T������5ĘއE��)���Y��z��t��R�mE��%n�5�A�3sr,��Ҿf vr��~��������2}6�v�S���u2��w�J�m47ʦ
�<��[�^��Ҳ;����?U�����J���WԘ�8t˵hYQ���?��0��Q��:���ADT|rM�yZ}FM�4�F$������j*	�riE@�ٕ7�\.UTJ�y�Ѱ��/{`k���|�M�P�C��Ύ����쉦��Z`|����%-���Ey�%)3��V}��>�>�i�'���0qy���m�Z���u}%f6�Y��QP�{Pٴ5qG5K���D������}]���SТ��4���V�nV@W!�Vd��KD5�Lm�7��s?�X�m�.���t�Ѫr��os�����җ`�����5��Q���|#�wܟ��#�g��m�$�	22~7���QVU5����!���xz�.����i;�����0s!���}tzCCFvL�ݠV441�Z6	Ztb��@����/i�W�-Ш)~�p{Q�s(]�61Ԯ�T�.���`C�!hC���q��,\��G�bW'��BTpx�E��خ�&���RR�[}�n/����9�� �fٶ^J��gdd���7��d�ro�8�� aF]M���a6�{�Y��.��#y2�mLv��ާbB/�~���V�<y�Vn<���5�a�$� |���͡u��,��@��s����1��{�cv�����{%N\o'��?�����6p�<"mkk;�wYl��_��ֽ{R��+/�����g�30�g���n�>�Gz|>�|�:%ڍKKK?���(���D;��_W�A�Q�;N��C���L���\�j
�.9�ͪ���>�t"?v�$F���'���ɝѧ`��r���VIDGG��9�j�)��Xg�xH�T���I�}m/q��O��Z��t��g��aG!�S��)f�}�=��+-Fd8����|=�[�k7�z)� � @K�Gr���O\�M15.>~�&U��8ϒ���?D,[0֎��U ��Jua�k���/�E坩�ʿ]=��������O�;�����j�Z��%��NL�*DH�\��C8ՍH,�2���H�;]��������{=�:��S��W'�#�
�sM^9����7���6�9���B��� �g9��ȥ���7e߷�u��������I=:S!�.[fHAvo�r�1*(w\��d�Z�6G�9���ҬGB6��'j��5�ύL�F�=�`wt����� 7��" ��>�u@v Zz#�xVM�О���7 ^�IIa��	�v�c���PT�RO-*�\��I�66���YL9Lh��}�4U��ZSs�*Nxt���Vl�܊�'�$�1y6�TRI��+��l�̸�(�'""
�#�K��22��q1�C���t->:>>>�=Ő� �	� =����[��Rx���׾�gi��*?,����VX�٠�K˖9���	"���H}�0j2w��؆;3l����V�As6��?�fI�z1}&х*Mb	���O܇���Q�T�"�@>�t������]��	��())��T��-E�'dK@F��E֧W|���%8�A+-eeeW��n'��n�������&�&�M��:���e2���/N��]��$YW�M ~>ބ��$����L�����U^�q�+::���f�*�Q3>	_D�4y�R������\\/�-�r����f� P�Iǵ[I􂉃_���ަ��,N�����k�o&�R2���wԌc䆶DX���a��*�������Rf�`�_�[U�	�*�;�#�%%%4ϳ�(
�i�Hi5�<~)���K� N�)A�_��X���+O�Ϋ�K�v��12����[ơ�U�uC���9�%�*݈���Ǖ/onș��3v�
��|*��mj_�j�K��oG 8帾���~�pw��VeJc#8w�	w�2A����wwN�9�a}~݆uv�_�7��3�;�G��`:�O��zYU�3r-HV,�!(���u e�܉��j&'x�g�D��(�[lOPDD<	fzzdBB���������#�O��_h;�����X2��@׉�LJ��3�?lQ���/q		���,*�y#SRR
J�rdi4��V��=�+͢g|�e<�0A��:^����qo��D>�s酵���-���'& ��|M�I�ݍ�SE�Z���3��lb(�zNt���W�Ic�Cy%s{��7�4�vȉUe0==�z���_TT4��d��q;Jv��ݭٚY�����`s/7�@�`���13�@7� �������;�l�}12�����:f�kGH\ ?e����t���O�y{��T1C��I��Ը��ߣ.��H���u��V��v��a#޺ki�i�N��Zh�b�6��k����PQ'��7d�Y̤q�,�����C���-��ÊSy]���S�(�@��)�#�܄��"|�ύM{ݜ���t���̀�x�YN��0j��J/������P��������~H�4�� �"r�F����\��lf�
"+)���U�"����vA̳:;#�#�3�Y%Vˊ�Bu��t�y�

@KhZ���8H`�{�(��J���ՋE�x������������	��3F7+S�ז/�5s�>�������db�߷���W��l�g���Q��6}f���x��M�-�^�=|�x��Q� 7�r��5�捓о�a���2-�t-�6�T����m`?���k�z���'1;�����)���&?���P=�cba�k���t�c�>j������w�~��ԝ;��I�� ����͹�x��N��F�e0t��U�g掻�ϊԫ�g�����V� �rpT�jÿY�w�|��F����2�'�\�#��OX��2XCt�����ɒ©�s�C(��b8M~o�F�.(W׾� ؕ�m�͎��f1��*��͓��5��D2�]s��,�7)\8�-���"��6W�b'�<j����D�~og���{^�*"��'�ۣ�E���|?�v.����s�����O�m�^]n���3-on�-�z�����p���6
2w�5'� ���:����vT�f|��:�u@��ǚS�+�}�Ɩ@�.��R�%!'�t�
U{G��3�x���{����q��� h���ۯK6 �����rs�UI���"/����Nipy2$��09�K kP���>%�o�2����V��Z�:imx�WSS#k�wĲ���c�j���	`y��F�u����q�,���K˭.f%V�k���2���\�%8M�L���_`�Ec8��C$:F#���Ϭ��;�t655a�R!H'������].��Q �̠^)�zt}���(!�����:���0���O�>����M,*b�c7�Z ����T8 �U)��b1幫��T�Rrr��"XV]��~����L�3n�R�����s��+/9�(���/ߘ99� �//����J�N�J	e �.��i�}����k�0T�������<�g��llJ����~���'��������(.mm�N�`Q�v /��b�j�$c��L����k�= ��������3� �k:��lV H�a���R�p�q�����A~�|�S%CUl����@�`�;\e1����V��ZԚ�~X`�����>����"�h�+y�r-ZN脚f�Q_����?[
�U)x�� ����wɬ�6N���<*q*�i�I^�-Ek�>f��At`�|m%+���vo��F%��O���	�t�;��g���R��gB��ϖ����lruee�؎�Nl��@s��́���5��<33�D&6����
��
{}X
�V��x�7_�����<M,"uQL�!�RSO��Q�H�[�ϸ��*��%[�{��_�_�6{\0B˂@�X܅��:���YN����$#�8T�K9�q���w�	9�з"�ٕҦ�4����Ś�_��6S}��
�ӄRo-��|6�8��l�L��Lm���c��ϡĂ�E%?�V�k��f���������N}��S4�Pn���j�-�����x�΁zoo������Bc}ˮ$�o���A[��WG���o�%Ս�����B�e���;'I��о��B�ؘ!ȍ�B�O��R�5*�ʦB��R��EF�jL�U4��a0�}�ѽ�j9�N��W+�%�I�����j���S����:@�L���eYEE�d���KZq`�[^���Vc��5�^jke)���*
�����&N��ަ}�<�\~,�"(9.������K�@�v�|cc#�Ir�C�̬��/2��g��U�v�޾}l���t��wLh���
�����Bz/a*2V���V��́�7��M�����hY���ǹ�� |u|�T�s� ̘���4����z��U���Jȳ�sJBD�P�z##c����V�����^���:P�dcn���?3244�����%�\�D#����a0[m�> #��t���oȆ�{H�p����k :l{aL�Sb��0��/i�W��V��fzP��~�7�J�#Ԭ�Q�����96)�wTV^��8:2�!��%_E`A%Mq�v�o��!..��f���]_�͡� :��P��@�> �877W�G����3<?��8�E.*��m4Q���HC��:�I��m��hU�y-Z�c�9e39�<���Zw��e\y����ӏ\�K���Uۆ�����^��q��HY�C�Z\x���{Kᇊ�_8:[X��+\��c*s9\��"�u�Ȕ������1� v7z� 3�a��}�U2K��۾@)�3?g���tR̩`,��&|`O�X
�Ըi��P���-������ʾ�H���?5 �&~��h7�������@g��8�E�q@��"!�
�q��x��3<=8��F�;�kB6�n�ȿg�m���Ol����pl|�v���Ä7Z�|�s���)��JO�ؘI��$�H�[�=�g�Ӊ������C$�I���T�@�p�,vt<
�m��;�X$R�����7��Jh�����7E]ʡs:tG<Lr.�x+&��l����s���߶�j���|�GK<���gX���1�ʏt�蕦l�&^z��	��^�$J$�@��J�ˍ�2�E(���Qs��T�/�*�Ni��lT�[A�/��F�\�n򭹷|��\�ױ?s:\��I����Q�U�ԓ'O�=r���8;;7uw�)lN8�P���I�
x���T��&M�>_�Pg��y]g�8��v�d�R*�����aEVB�m"�т��8=t�@�H�K�����7����/����W�[��S��Ù���P�n���%ݪ{ m���ʇW�4
鏭�jaqpp�:EED~x�]?i�4�2
�h��P]�L��
��d���N�gZM��a'P�G�����������+�4��V*؄��t�wt
d����,�|�<Y�S�>e���`�w/2@�- �+�\��I�'q��L��wװ����P��)g;������:�$��&A�>�ŮU�j������JH�۶�ꆯ(H��ê��^�n��y�+��T�W�Z3��{�t��mhP�6.�;{zF��YϺ=t�"&�>�;�y������iD���HHޔ����{6������}�J5�C����I���U@�W��@�����8�_ ܿ�hɄrpp��r��^N�}{���2����G����I�pjZS+҉&��L����MU��d$�j:�圽����vL����d��D:�oV
�)�K��k��fal��%
�W���yۤ$��c8S��&��hJK�wc	�V�"7O�!5\�&�4M���FE0IɎ��l�6�R�������vSb[���r�������S;;30���ǡ�$��{��_x�xF+z�~����l>�s�.DuN���%���62
/#�m�![܍���:�Pp5?7w�h��bHh� ��)��:�A䶛��ҩ���]�͢/LM-�h��<�}������w��6��?�h; �>3�?u���/to
:�788h>E�Y�N-����'����%�I�m���~M<�'�o}k���p�������q�dL�{gg����2 \����U����A�0tIy��4��=
���q�i('���h9�OUUU��%<�[?��a�~���RPP,Z���<3���9;�
���#X������<`�Z0��nq��y:_\�ؕ05�[��&���"L�W�{ Ht(]�C�0�������X����OxU������;�bf�u؂�X��4 ��##?e�|�v�Y��-�	���j��������>��Ʀ$^�ⷔ9e�{j��.p�s�N�}�Z=9	1p�l���o$:��;} �ןJ����k?q�`��_����T^^n{0�]#%%���N���50�U����w9%�u�ᬵ��t�(�X�~Т��Չ�޼���ʵ���iO��;if�#XLwD�mѷ�tdH�-��6*L����i�<z�M���߰�3��B��^Q�'7p�8_��=�y7�.v��R��]l&m�f�V��{���^�-,�R�e|���lhl� $�?j]�"��F����B�.=7���Ą��d)�����{]���!!!�**�33��x����ii����[b^)�ca9t9ЫWn����+I%���t~��Ѵ���ͫPQņR�q�67��99��)�=�*ֺ�?��� B��������U����$Oh�Or�:�'���I� ������jo6�;��^%�Dpiշjjk7��1������M�����^��U�x�w�a�R�P�ʌӍG0�y2��S;;���f�_H�Z?+�^E��U���fyS^�x�����m{S�m��'P��]4�Yn�4;D�xk�ii���-�k_��j͉k�<��4qm���I�qD��斃^'����ց=v�~znN33;�Mwɨ�!$��@�g��iC����oG@:�j
�~�ỿ\U�I��+ݚl�UB_��V�X瞘N )!Ѻ��qX[�Q��y"�p���Q�Ԛ,���ٰ��:@��֔Rzz�+��nĶ��F}�q�Ц2�S�%TQ'j������,*�+�]��5ߘ��]PVY���p�E9i��Аu�R���<�]�=c%���W̻�K��῿/	�-28x��z�khdtg�1.
�?�x�#�f�C��㩗�vJ�S�\8�h��>w�:��j�4ժS�Zʧ"�w�Z!�0$�-�WS����U8�8wYeuE�[I�13�J�xkG����I�5���m�7T��	I������y�
߀A��Y!Cl����A��>�`R��J/���֠�t=�P5+K���aԄOڭuc,���	��V�*	�i{��H��%Nl�D��?\̻,r9���}񠨤Ģ߁�`�������<��A��>b��Rw��("���+���_c%��s�8��75����^q_Q��H�t4ь�)����f)��%��pլĊS\�|aZZn�#J�'R��鮵[�N�
�$r�^�[��l�_ȡ��ֲ��R�=�	~��P8wU5|�@��?�;$��T8��[U�������"�W�� �p�R�CD炫�	뫐�܃��F�kZLL̿��fee�m�~�npc���t͐�UX�Əc��ucB71���V"�m�233u��(� ����N�����A6�K�Lw����lg͢w�A��=��z�Ͻt�M�c�����z����]�I�oh甛r�ˌ�?���6��JJk���F��5�����Ko�Y�X��͑��B ��kM���j�#�'��Į�w*k�y؉>>e���u,�&V~Op�T	m�S��� ����:��xpy��S��ƚ��A5��yt��F?.(k��:�=��]"�K���!����F�/�{�.�ĖS�E7�q�E�)z��ۮ�����$������'47�jT�]%~Xr< ̭?�ĭ%�N��1l�^�[\��!�YH�K4��@�N� ����x��{>���WrI|n�J���n'�5=���w��c%� E���=�v�-(�� ��5:ZX#Ia>E���h����@<:�"���1�{�!+++4�i���kܑ�n웟T�ћ���up`�$�j1D����k�ŕ���g��LL]RL�W���剦��N}șڅ�NNM_:�˟6d�����S6\\�/�U$�:���T�����-v�����*��2}���w����G�C�|�C�=������xg�4���@__: vyyY*`����~q@4#m��s�Ύj:C���Z�% ^�~� ���Nv�������pL��,$��u��˾pXڦ������TT����y��%Ʊ�F�FN�&��H��s5�J)�y�%	�O�66(""�}�DZ�$�#������rG�6��B9 E==����π���q����{ �ٮv>S��Nˤ�����❷w��@�afU��vi���[�FhFeè�ԯ83�\���N�Z���ο#mS:2�藩�S��n��	��ߟ�>��\ �r���H�o��7S�q�،i�:�������H�gfn.tm�0&>����qD���i�8�[�͝�
����.�hXVs�xA|�~D���L�yr�d�3�X��O�C��t�KR)yDX��߿�O�6SW�sRA@7LR�:]�����,m��E����UdN֘��c�����f[�{�_�Ҥ~j�cu�b�U�t�m,���#d���Ag�S*vJ����o[�?���슳���w��p$xv �1��Z�B������C�v2K���>oJ�$B�u����,ոw�����t����B�	�գ��߻�(..P/������	t�����5;���G
Y:�NDnJ+��;�L�wi��i��m��󆀽��u�C.U � ɹ߁� �30-�	('5�Y���A���i��%�K��B:,bUZ�[M�K9�
����N�-O��<��)_��/{D�����S��>��>1.�����|QR9,�6�	�
l�I�w�xy��g�}`�����]�NNQ��h��;w�7d�
�Js��ש*�u�v��]_��������V6�k�-��y�����'�95k?��=��,*.��$ ��3�1��xH�!����7��E[�L���4f�ƾ��Nc�vc۶m�Nnl���{ߟ��}�^{��9g����,���KpqT����Z���F���͹��'����m���:n-�Z�7�o��m��3~�t�mJ�+_����}��v�</�ice��:����v
l8n���K�Q�pI{6l��L{zG��:19�<�'�Ńċ�헻��x��hҒ��QQ���@᫺$����|����)/�>]B1�z����/[^JY]NI\q�O�kl~��U�i�&�ksl�-��/�Ҕ��r�K)6o�L���U��uw|*S/︘ndOU��|�f�?LPd��qa��c��������o�G�m‛�,Hr{n��V���a������[��i��;=ig!�����~U�7��R\��� {����˗�����wM��K4��AEx��a--\qǆ�����XX�s�le!��fu������W4@��iR��ydBz���.����F8U'�r�k�$��+kjF,,(��,X*O�
]C�Ԉ�г�b�'K�-�:?[�?����:��_	���D�$t����@W��]M��ѹ C�� FL�9I�>)�-abR۳S��M���[F}��0IX~��S/K}`%J���;a�қ����t!�tqܹ4u�,U����}�Ě�/��o��n�,KXAI�S��<3_y�rw1Ђ64}��	��{,(��0���a�pq��q��d?�B���·~p��&��5J��y8?Wt(\sp\>��/O��َ��c����	&��Y<��&��kFv7D��g���ٝ������򋚐�Fm�H���]n�.wK"ʁ"����͔��}����[�G,��FW�d��)��~���{�[�
�����Ы���S����j]�"�N�+�@�nד"��'Ke9{�[���6��GpvI�������GG'x�G�A�뎈��4&)���Z��
���/���Y����a��J�M�l5/g��c��!!����'n�z���v��#kK�]���0�B��<Q{ta�g���U��{����sk*�W�=Iߝ�&���ʘAufVՇ�/��t �~����Y���~��V7��ʙ=;�B\��w#+�������X�,e$"��Q-�W�����m��(Ui�]v�b3�����v��i���"��& �>[H�Mj�o���g|�E�˨��JJ��΋�5E~�r�#C��N��Iބ�����ˡ������#�-˕�ａ���vq����Z�C������!geŀ����l�Lq��j� �l '#{�WΈ�����i�{�c�s���V�JWC{v!��!�#�Tg0������U��	�_��:\]�=���_�x+x��Pttu'f�W�<_+w^�y�4PP�t̯�fs�56$���x��@A�b/��f攠c��ݲ�;<<�`����>'����@�JP\U�!���FρZ��(8�U��MOEg��	��:��Eff%����ե$�%58�*ИK�+�k�-y=@-l��ɠ��g�w`�R�i�M�QB%��D�\BI���X��ų�M뀸e�	8n3�D��Zz?�*�7��,�qJ�@Zo�A�i��b-�y���C����R���}y�|8����q�B�p��sy���qFЧ�ˆ��i�<�|w}�_Y.��#�x*v���.'g�|!,�8޶h� VkJ&ǐJM�Ŭ\���sP�M�T���������9k"�����1��v5�v��rv�%3���p'����hG�
��l[����Eʇ�]~�5��Mg��S%s��'��݊�||g�(s���'���˕d��!�]ym^��@{Ym^�3�^��o;���I�m��A�'�@�m��cw���
��E&���$��"�Ы�o����z�����8qF��"�:Ƽ�+_���KLL�׌�}����Gu���5����wk�!Z4A��q;��'������V� �}S6[��uQ�t�˕X�FEG'z��y����%k�{kK�`��0�c�Y�]9���k��͟��"�����2�L����)�m��nii]�6���XN�al�h�&&�hh_Z۞�g�ſ��p�����t�.����������w�"����z�#�zo��Tz���8��<��H����c�B����nv�/9|e7��N=:�\�zarg!�S�M�S%t�����?Qh+��'�?���wQ/�����򞐔�1�	���U~��U𸿽��OC�f�&��JI$nJR�q���k[�1|�yjz��f��A���'�}#��j�ߨ��M�9S����k� $��}�z]���n�ǲ���>%����z���I�Ua����Q���m�p^�m�I�p����y�_+����q�^R�#��(�/���Kd�sуr�xT� :��h2�y���v&44��_�v'�9��8C�
[�' ��;Q�W�z��-?a���P����t"��:��09(�4�]��[���S��˲�Q6�|Ķe��4)P���6rJ���S����Jm�������%=$��|��"_	�$�%qߊ��,��������ُ˫���Ǹ?�I��y-���-�^�����V���Р}�3�v�3"B}Or�y�78��{ܙ�〃G�1�"���i�}M�#�47l� �W�Ҁo�V�)c�C��Ot4��ϟ+^m�u �b�yw)�]n�Ct/e$a�X�a{�azk �u���h�
��Q��_���aYˋ/�m���n�E'$>��x���'��-�#�Y&�������j�c�%�&w7��7H�)w�}�[��Ӫi��s�֘�dI�A�wtɺ�gR�Z������	�6��@�ZN+*1��3��4�� '�u�۵�*M�����g�k��M^6���bH��阉�j��$b�ц�`,e�qDa�I ����5��q���y�i�gh`R�P0��q��[Zヾ����.�����X�&3c��)=4��e,���~�Wel�r��58�O�>�+0�b /��R�� '�}24��Y��4!X�fu�uC�������^*j�S����٣2�X��x���x�rtr��0��" ��y{l�B��6LK�Z#J7^��$79J���nw�%� <�n���'@#M�&
�9�����I���lQqPǑC�}gʃ�C��D����|�{=���$JS��0�R�(�]���ɊA�2͗�%���H2Q�?��E���+�om���g8�~,��*PGM�}}�ɖQ��3H����U��q8[�)_�dQ�x�აUU5uʰ��������^N�N�v���y�����#�ǭw����p�64_xa����������%DDDO$�z!�:�o�Dˋ�s{_���>�4H� �(W���*��������E�G���r�M�*�aX[�T�ܤ�z��-�ݺn�q�����-QDo�@���A�iPϛ?�CݡR�w��,��-�U�r�&��H��=Z���-ˊ!���?_��Z�︑ܐ��Vm�m�S�,��R3�(��/- V��o�آV�dx\�-��_�ߣ}���c�F����ƹp���1F�ƻB���ر�U^������8���PڈK�����k�`��4�[�����ۓ�G|��{���}�q�����L{q�����a�ǫ�Q`�j�1x	�>v^$�j.����'\� R&>l"�gZ�.`��u�v͹==��aGG�y�w�~Ü��W?hy�.�����c��^`�=-������h��y��!&:��Z�I��\���s���8��AC���p=W�������)ѹg��ԣ�]q��=^�%䒐�;`=O��=Ԣ"꿎s��Ɛ���^(����!AjkKk�V��^(���/����/�����`��o�ir{�sd��p���a=x���f-?9�DgG%k~U�L=�$S�ݑ���l>vǙ�a���K:kdd��Al�D�X&(��������L����8�
�aMF�o�bll;Ӯ�BE�.}>�ƿ���T`Y�H{/��ѐ.�Oه_IV���ga
K�ȣD'���GF$����44�3�")W�}���}'���>��08���͒�S��6�,�	�Z�ΕY��ȫ�#�������j���*N�b��5��ĺ�s�:���Q�1��?��gd,�W�F+~+�t*���0��M�!��"X^MX����:�(~�|���o�}��w���z�4V)�C�uuu$,$_6Mu�Ld_P�>�����x.���g�c~�s0t�l��ypv�������}agk���S�����	��(5kyG��fs 3��Y��p�|�V�Q�Z�8����==i�E�s�4Q�+{>\ �Q����w?���	���_$P�@���8��V��Y2�����!8fw8>��8I����Uh�_d��t��c�}¶�7��%�s��+����Dv���l��/ �@�;$6onw��: ���'�m?�е0�X��Ӷ��S����Uhm�/���,�D~2�֋p��V�_L����E�NA1@9�}����(��Dq������k�W.	YM�G9�"~� ��%�OuRkU�bT�,�4�~|��k_{Q��S���9���k	��~��~t%$(�5Kɥ'��������b�U�њti阎�z����)J�K�LU�x�z�w]t��)r��c=��VƯ�/����(�RU�t:"��r��]b��ky�!_/��Ic T��u�e)ϟc�L�h��f�8�BH�P�Re�ĉ�O ��x�����~ka;B�:$�{�v�B�w�C� �E��W~�
X^�P3��=## �>R�����c7�W���]�J��2��?~vGsxLN]��_��p{��j�Y�{k�H:�����	�s-hdՇ��^��Ñ T) ����nD%ϜA�������������6�<���o2���Iܦ�{q���=���T��?�����7��A�S�k�pS��-���æ���q���<��E�~
����O��{�\����?��J �t�!߀�Ԡ~]ԁ�̫��l��a,����z~w�΁&��Ît��e��U��u��vf���L�|~��oDy���K� dI�f�9�zi:٣ت�Ǿ�&'o�_vK"���m26��f�f�;#�Kw��!�k��O�iC�ߊDa�!���4$� �����5V_�i��I��m�c_���;��s��4�HA��	�+	$���r@W?p4ݯ���MI��@���j���$9�Հ
�_���y�+�������|��~�|!@a}�7���fu,��Tp#b|퓥%B�R�<Ug�]X��2���b�K�Q�
	dh��M����\=rL���b�r}�*z*�C�����J���Mm��<��E=zl��]8��|�)�%����\kw\2��@�z-�*��{ɖJ�i�mT��+���:?��9�V9��?:ړ悎&pJ��FO�۳�E5[U<�s݋g�D��Z}��f�8s%��ѠR]�� �*|�ɘ,��`|�N4�?�U�q&dhz
�Kܤ]���֠��ɔK���-��'@o9�>4z��y�S�N	�1���yk�ߠ�����K���|ߘ*��8m�ׇ]?�_� ͏��"U�`��9@�$N�ö�K)�7m{�W0����zr��_�PG����j�M�T�KHo�c��ib�n��X��is�M�����b��h\1�f٫�e��7�凓6���������7Þ�O#`�Il�[d��D�8�,$����o���O6�����0c��!���Hʄ8ˤ�~�
|W��e�pk�(:� /��6'碋��ju{��2l�&޼�x?l�i�hc��(W��u�'ѥ�N/H��J]Cfv����\������km�f���^��V��X���J���ȡ��YW��� �ⳣwK�{4W�Q^�����-C�����P}���)���#f&��cA_��gb���WB/g�;��|��J��@e$��J�Z�x���g1�-�����qgڼ#	(�Jpg�+��CykƂ���`��U���ja��s��MٖV��g9�E��>(Vo��~���}F�ZG�zM4>�ۑt^ ������,�؄#w��:�78,W���~�Π����-I�Cm���~��@�ƌPnuf9�˕Id�Q�����g�@�	��J�ƣ�A�1yԿ���������[�E�Ua��_�̀�h�$��Εk�?�R�AW����dMR�~���3;�rv�~ET��'�"e��� `�0��x( EzF���vA�a��"�����E��c�>�~�z�ћ�<^�>8�x�T&I^0+�r~m����?����a2x��,֙/k�c��o�/�
7~�'�������;1nj1��xR0�^��<17���z� �Ktu[���-����}�����]�N�y5���6��!7�]j���7?���jo_��L{E��~:����x��;����w0O1�Zg$���:��A���r�4\^u\3E�%����+N@�mH��P#p�s�\x�[�B`����2wf��t�C1���S�3����jz3G�K嶮��	}�@8����u��;����˳�E�Ņ��x����������74P�����o���p:j���sD��D�Pb͊��7Y��[S����[��Ԍ8I���y�ے��Ta��=�>��]�^���6��e������@�c��_�1�(6RD|���i�o���	쬳�l���Λ��d��
c�)�A�1_�_�b��3�.תX�GjѠ����C�J�{T��-�,�I�-I��j��y��7���K��"34��l����1���_�`h���-�8X-V�#?�6%�����7�ƻ�,Qw���*B&�A��p���-MO�����Ȋj�Ň�;HK�z��Q,R[l����A!�Uk������Ri�/q����>(���%�IC�:�<�OO�#w�N��Z,t�x,�"�w+� �� �s��.,b	��Cq�����a76?�O&	&��$�#JR�?�F-x�W؊�襧�����w�� k-3bԙJ�F;�����}�����M�^4%{R��/��,+˽P���������j�Bi��[(�,�������KP�xnGLHfF5�*rI/�]��	�w=䚶U�O"�ӎ����z������T�Pu �=���FuI�4W�E,���T�7d^�;���biy;��\g������>�
f�]�֤��:��Z�t��OHߍ��]����w�M�|^� ��/1�[��@#��,F��gE�Zf����3&�LG�eq��֖H�V����_2;�CK��qp�g(��m&�v�d�Hz����N���;��aC�Y�Q�oE�es&�r��(i%���9+�O�㩀A�W�	8�I�lɀ�碷,�$����� �7wroyW��uu�@���*>��atKUe��5wKyˋ�o�����
��d�5�����k�\��,O�}�)*:���b��PO�Y�g�^!�~F`�Ι�vB�/x�W,Xlf(�R�z]*4N��p��=$�d�������1#GǆW����Β��Io����	���;�Xx�'˧�����+��Xc��lF��מ��q/d���4���ut����߿sy�'����G�
@.���є<ڿ�&��B��0�5���yJ���_F�	�E:қ�>�5*�Y#	z�^2M@�P]ͽ���T��������@�B(z�t��{ɍ����Y�|�ІB&��J#
@7K����|�z�\ɛV��VY^��e��]4��Q-�cM��#���FoL�����<ʕ)�i���H�e��?�f/�e�W9�6��R��m-YL�p�s����1,�~]����=���rۙ��T3���CVw�>	r��bL�Y�(��0.�őS(�]�ce#ES#�z�&] r""�kPB��3[_Ih3'��r�e�z3<�k&��+�&'fL�L�Xl�a7�!��fu5�9��$�a��W7��_�k��T4���yG�>�W]ɬ�j��^���x�;t�q{�c!�$�����X<Y���S<��G���ޛ�(�ڷ�������ɫ�`�O��;��	$�p���q"�������MA�wh��,�[�����\};Ma_�� ��F]�2jK�����������rsm;W��;�w����H��a�6�뺐�8�ͅ�L�X����,&Kڎf�Xy���z��Ooo����9i8�H%%������Y%- �<G���oX�
mc�,!���C���:[�f�~�9���0̣�Y.t�7-�l�|�^�U����>�/(W���[t�ʶR�j����L�wK�Rj�yˁ�1�ʇE,��w��δ�&�Ê]��"J}x�Q��*U<�"��G�0��=�$�����@R��4?��(�?��Hv<�>+��Ӻ0�|~$����s���r��>�t*����߁���?�MP�'Rm�JVɖ���$��)����q� ����9�,:q~R��n��p���Q��x�	:�a]��a>Px��E|��Q#|�̑����o����D|@SO�q�/U�~����Yk����p��'X��:M�� E�kK�K��ςٯɰæ��$Kꑳ*�*n\��{tU����o��<aa�ɸ�w�����sd)�R���<.c&
��ň]tp]��RQ�,����0׽8ݝ����_�G���b:
��ƅ��p�����e���Ю��в��z�S��Hc#34T=y6ַ����������\6X0�+�v�77���V��:�;i\�U�ݬ�:1�<{2�q�����A��}�Y;�3�ը^w��g�ǟ��Ϗ�;m?��a�&�"���2�!�k5a��v�R��kfQt�u�+..���?i{]>֜��H���2t�˹��b=W����h����'g2��}h88!5���00�����0!����i����}�1.1��rj�A@���,5Tn�lO$"� �bk����{��U��c�@O'�VƙܔY	���ʟ���(����E��׿�a~�Z\�Ts����0_&� q��f��""=���M����>J��.D�R[,��4��j������AVEa^VZ�!�.�%l��tͭ��	"��r��p[�{-<��M�����/���q��O�@ A�u����P;ma�+!������"��S����"�NL�/^%?�ڮ5��$^�e�:�|�f��n�ҭ9^Jnmm�3i�������K�1��X��p�W�����Mw�"�o����4r����.

��;kQ=��
X�ܛ_7�d(+�,�^� �ZsR3�0婾��s�~����
�ߪ�aV�{F4���������X�GSvZ���A4�%f�#Sh9
�x�����A·Vg��S#�C<<<Q1�q�"T�/���%DӰY�����o�h�����ߟ�p��֭S11M?��	�[,�%;�O՟�8�r��w�
�'
u�6�N05`9�-�K;z~�Ӣ�_v��K:�'���w}y
|8���!��LG�y�*2\�1�R�m��V�<k�๺+_��=d����k�+Ȑ��� I	�;DPٓ�Y�&�8�&�>!�����l�qᕷ�t���a(�� GSI��Q	����W�A�=?����z+��m���N���X�C��.rEs+�2ʖ���z�!�@iHH�X[[+�GH��41�����k+��ݭK����/2�'�F�:g;�Ɍ�׻m�'����U��Z���vԇ�F#K�7ؔ��!��D �_^�)�+=a�����l4�@���qr._w�@7�kd�h���T@�~�fZ�)Ԇ�0�C�G�T_��~����5I��[�d� ��6���,�3�Zp�������cӠ>�����F�ې�f2�Ea����sj��g׍��%
�}Wz��y���Z�0��A�t}�W�&L^w'��ytT�͗A(G!-�(�o��r�(?5���:�zJZ�zi�44���W���2++J*)�m���f�N��9�+��2��{P�g�����ms[g�KZ�_Q����O;o�QNR���r�M�X0&��O oU��b���^����n���� ����q[�O�����K�������9]"���bѭj`��!j�������{���|zI�	�
���U�%ݵ�{s�"e�,�>f5_�+���T2�hEX�&�Í�>x�D9�/��J7ܪ�042B͵���g�c�t���n^.p"%g;�^�UA!�=
�]{x�7	��Id������T_�}�N���B	�������J�l���E{ͻ�IDM1y�z��I�, '��m�3�X[���V����Tva.ʕYo��=�q��6�Ԍ�Wz݄5���\���5WPl��1�v��	.�"Ţ7O2�L��s����{�|Y�� n"�E$L�wσRx�8��/6��A���p�p�R�����G,
�Dk�W �j�������h�=�^�z|�;��y������_�҅#��b�4VӖ��A�樖<꿝o���v�����j�_||�(�ʶʸ{�z�F�m��-O��{*�jΛ�Rl6��r�}�j�Nm������"���'�m���!���g��sp�͑q7�B�&�#!��E��P�419K�C�F=+?%��MO���5g�|�����)[��V�I�%�s`�&1��Ց��3ô{NѲR�f�����nX�6���s�
-)�PŢ�+=��@��-vK�˅e��N��q�U�[��V'V���y!�r�:�� �|&��Y��@��r"f��rfv|�J���r��B�.�P$B��^*���z~��3�ǐnьU/��q�m�̰���0ٝ'�iK���Ѐ'���)a''��������v�M��f���lˇ��l-�n��7z�����2'�ښ�)1Hԟ��~�%�7/��䳧}�P�2E��:kZ��Tq�`c|.��� ,�S?�
Ü�w�nU/��~��t4�q��U17��`%�u����F�E�5�n���ݬP��|O*L�����VeL�	Ȕ)�>��u��������������7��ɭyI[�m��Es�hBc��^F�a��G\l��t5��F���E��R��Bm�vׂ�P)1yأGb/�K�6������sm0��HZ/���`�.��"�h; �r���\k�b��NmZ6Wf/s���У��)�a%	����e��GD_���� �f�V��V+�lG������|Q,��w�U<#!xo��<n�<u55�RR��1�P�킭٭�?/2b�XX�XcB���sj���X�=֤@�=b�Δf��p�����Lج��=t�q�dv��C^sN�C��u����c�t���G�,��ф?��!�����W��l���>�5�Ó����mR֞�TqZ`��>"b��zQ��󞢳�QR���QNP
w��߈N-�_�{hHxx�9�!���UTG�~O���I�������'�&���%��P����z�'әj��[���4�=[�~K.���&2�V����M���!�����mM�31d��,��X�פI���(��3r��n�QQQ+x0��1���s�+���F>��ap��EE�-��T��z�����$e�rFKQR@�e��x��)�0�6�u���3��;@pϷ�!�g�>�Dm
��J����e�"�F��ki�W����$��J}s3�;=[,��NNhٽ3�}i'.��<���pI�D>_K�dHEDlL���/n.Hּ��R�*#3��&���X��m%;;�9A���hx�p-'�ZJ@��Ǧ\��⹓�Rs����p����J��-xͯO��F$M���t�"NB��q	��ƭ���%%*7��O�_���m�lB��Y����xb'������Ce���J����x�!LJm�a s�Onb~�zZT�a�uÊ���s��{�wۓ��(x�"W�
���e��ӬP��S5��b�=��$+l��U?�n��рjsNU:ްio�@^Qq�mUf3ʒ��v��;�u}U,�"Aeb��GO��і��-�m�֖N�|7�sS[�(ǒb�c��#z�.B�9��W�p�OKKq�S&�m�zuz�R�}A�'$���!��I2�
,J�Ҏ���]�::�2�T�Yă�c�:�:8tKf�+ъuܖ�iP'k��I����a�����᧺�7~�=H՝rXߥ}!͕SQYR��H�`2�{��BL.ro�#JH�#�1�XP�GǓ\����*��cj"���Z1�({dDH�VY���km�¼��nk���DKk�h�j֗;ڍ�a�c����uf�]d�%����O�mc�����ͷ��ui�WՖ�t'<�?p������Z Ǿ^=���Y�� B�ͱ��)\��]Fl̢=I���I*�U�A�����Qn�S�VPe�x����b5�H�}j�զ5R孊γZP��J.	rqmi���{�(}���a���D�l+G�Q2~0��DX�d���U5����P��5oq�E�:D��p��!Z�n2Vh?����e���)�g4�Ltت�����b����!���A�`��ft�A��;F��tw����}�|?`�)P{����f���iJ-�bE��5��
�A:t���D��J%2s�QZ Y��{�NQ���{(D���.��u&&&�:ͥ8���&�A5]�`.""�)�D�?���;]j�>�Z���d<\��e��Z�G���6�dH���l�';�ȗl�?��j�J���QOεJ�Hq����֖���ڡNx��߀;O��7�~9��6殶X�0 �Yb"1��D��O��;nu�u���;C>���u#��հr�֨Y��=�`{}����0�H㠌�%���N5�UI�����Zh�ƣ�)"v�J^�����cv��|-���׮�0рZZ��������UE�ĕ��(��H ����ui)�C�P�2cx�ZZ��K	dU^V�����\BFo�q�-��#����Hsg�Yž��E1������A�<����
��@�$��^���ɜ^�<�7�G����� �o�4Q*l�\8����%��B�������U'�Ƈ�J�� � i�>��:֤�c�I�&��Aa�IQ���ӝy�$�����B�
O_E������1�j�����}����<�'��xz��L�-����}bi�o�q��(JQ�(����K8b"�$N�KeMK]��uj�^�q���ܑ}"5C��ѧ��M��Ȏ=��9�9B8g�D��܁�a��"O��P]|�7k���rW��`6A��'F�7)))�ą�$�|�Oų�㊧�n�.��r��)ei��8&�teTKmg���c����B"92D�	�C@?�i7~�{O��fPJ���������
����كs3e.���/W7�8[�:!W���ڔ�?9	�TG緵��~D�VP�����)�������h�!�-�� �8;Xe����:38A�+�m��L�� �)��֘ԕ��#,ͻ˚v�
&0�p�I��O�d�� #��e���;�W`p�'pB﯇q)��^a��^G������+*���]�l���hܦ!/�C.gT���S��[k��R\R���N�Ӥ �fM]n��>eN�$�Ȇ��=�[<�T"�l����m��γ��&����IPT�/����C��H۰�BeÕ+��T�xm�� إ��ɛ�a'j �\�!#5{�8��8ދ�r�;Қ������s���VWS���5;C�+&UK���l��'H'`P�/ w�)���R��K�l/�設����	"�Mz$��8Oy8�	��9�3Q�Y�.o]G{ih{:F��nx�������
�����!����X��:Y�o*��XO�!	���isy�(ꤠF��go=��x0����Q$�xx�&k�0ӗ+�^=�kթ��9xP��k|��淈��-�'�W��4�6�˞�Y����13VY��!�#�z����_�Fi��FhQ� ����-�����>��Zj��]j2������-y��*b�2�d8#�����S��4�E�{T�A�;�n��	���+W�������Fĩ�����L~�&�U��;���m(�M��ϕr�h�F/OC��J��s���ۻ�r�}�#�Ic@}uJ$_oP�ʵg~<��PӞI(�2&V��R�9ᱵE\��m�09�G�#~zf��r`���cu612j�$A�S�O�,*�0��O!�B��{\�G^~V���kB}q�q��1�l!*`��໡���23{k��/$@�Jrr�b�V=���Y�@H��h�\���;R�L�G���]���0�r:�;�zF,AV�<����.Q�5��_�z^�j����稛��{�����g���7{��'M���gu�9�e5ߜ[�^�[��g����5�������mcPj.q�.T>���5B��:��qA`�]j���.\T�wh�轑	R�=R{*��! *%�3�?M,/Z�L�&�J�V�R�#le�l�v��_\?�A�A�$-��?[��a��=����Q�1�A�ł�=xl����~�+O��`^(ݸ��]Z�g��-;��5�xB����k��z�"��Q�&�d����%}����z���R�a��}�_�|̱Cޒy�JM�������L��f�V���r`E���� v���Y=<*����D^PG�	�5�爝�M �����ax6�Ͼ���Ə��ٍb�����9N���6���C;n-L|��3@�ܕ>y�&�WԒI=�,r�}����-~���{ں��(�m�ϟ�,�X��5�"̘�}���� �z���MM�a�b!,�"h��@)c�ӍF�Φ�C�"ż�:�ʫe'� �p}:�V\��5u��U֬��#��f���|I�FDU|_���d�+����V�c���F��Ӣt�~�|�3a�\�ڀ�(-u�Xj���ad�qݸ��_�j�ө]�m��שM�<�}��=������_|��:�:�}a]en���z��E�v�����M�"V�=�~�U�] B!��T����[����*ZK��ٮo����Q6) Ɗ>dVx���U�$��o�^�J_�,#A_���jԿ6��bq���i��,T0#��o)�����z�]*	�%���E�:�<�Ѕ׺X�^3���X
a��8#\PgŐϜ��1To�7���N�!��I��;�'=Q^��u*��Kl|`k#�L�����s~y�	tG52�5-�N-~	S�"Ӥ�5�3��@A�Y�j퉌c\��`��E����~9����q/��=�(X�����Y���a��"Y��A$�d�ܡ��`������:���)M�)J
Ҩ��з���u����Cm���4�4z�LRf;����wƾ8�k���K��ҭ�*~�G\ԉ��7H��B��E����-���v|�����-�<9��幀wJ���H��|$F�(*_�[V�8����0���R̶l@\(,��AS�V�E�=�~�`�� �/!A��X��'�s��ɣHL�$8����a�VJ�F���g� "D�hN
�Zǎ�՘ĕ!�)��أ(�ƴ�Λ��)�`kR��+��o��(@��)F�d+���H�/2�Fy<QDm�d�X���S�R
�6���~�Z��l�r�#�$)�hT˳rF��@��G��Uɤ�9ot��6�l�Af���"$/���RеZ&��ip���r�R�1 �E�ɏ��2A�%���o[G_�<����
Y�� ꊐ�1=���*�E�"���Kj�F�Zz@O��dV󄈔�4�2�����X�O��X�����z����f���fI���V)ʀY���rɳQ�J+�!#�0��V*��a���w�(K"�X`�`s�%s�Ix�X*?���M0A�4�I�^�gA\�pz���O�=Hݰ1��9_��s�?�^ʐln�|!`�ɕi�J���J��ƕ�v��Ç	��6vp�o|Ӊ	n0�lb,�G�I��#
me�.p ^|�&�*b��N)P�D1�ѡ����K��]71C�h��[�bd���9��9�B�#�z/�Z�D~�p�24OI��~U��k����Ph+�j_�|{j��o.�/Y�oH����@��_�����l4k����أKi�2o-g�@3Yb��f���w��z�������If���(�.��/88�%��?��s�T�9{..eQ(Y����v�Y	qq�h����9��u��ܸ�S�!x��j��s�E@xX�_�޹�M8�@�L��Z��E���ΕZ�;�u�q	~�Tl�bY% E��e_H#%oZ0&b�������N�����
ߣ�^�YXX*yX	<�*��Dn?H�E
!É6�&Jb3���]u�0�s�tuu�3)&ʌ?zaS�{��E�ϭ: �|ϱ{�]�m庇f��Z���Xо^c�X�kSwm+�����-cQ�9�r������ta���p��S��L)x��^$[�!��~=@����@Yq'�lU$h]
�SRr�2���f';CȵV�,���hWa�j�Q�J���h���KHI��hf�����J�C�E�Ɛ!��V+���^�Sk�mh��?�v&VQ�E� �q�U����ͦI�~�0C�^( ����W� dg����+��v��K����S���{i���n���n��f�c����|���?;;�[O��f
�$75��B���Ո�輁1�X�f���{�y5LѤWK��ۑ)��|�S�FB�[*.�ՌW��UMs~~�Y �ڄ�Pݜ3I�_�Br�I�����,<H6!�Q�� UL9��~P�j
��Dg!���?�^k���6K����h��p���	r0���Y�Ὼ�r|�IE�`�QƋ�����Qc�~��PYT��ޔF�"��S�����<��B�b�0����(�/��v����|��T2���r�F����R�:�w�RѬx��!�qz���Q����@��,]�:��t� ĕp�Y_�O`$����esk�-����n	]�6��[����;�76�T?�t����P���XL�NS�$�U9s�}-+�;�Lg��M-�����GO4@kgR�KEǠ]w��ύ������n�7l�%�(�?;�����	�-LH��]��8z{'�e�K���yԷ]��'�q��;��
��4��e����2MY܇���<���𮄆�4�vs�������P��%Q��=&ZHH�'II8
Ư�Vjj�-���A�љb4�	����Y���6��UZ<�J
8������nƉ:h�R���(`�3'��K��,˳x'D@�'t<M����)�O�?����z��7�F�����S������+Z�|��B�?_#tlm�U���SUP��M19R��(ҋ���Y�����ԓ%����Z����l�E<��Gn9���Wl�8BY>��3d�������ʅ�KN�������K��d�$��%�Y��K���8�^���ڇ�M���fƌ���������9��} %O����0�-hlej'�[�ٜ�����?d�/έQ*�b�*�*�L/��@,�L���{u�B4�-�;(��d��vYM��������J˗�h��G63���rƖ�@��Nt��?X�1��M!��^D���3?n�56>��9��90���^y�e6Li�&��6���K}�+63g[j${�Si�O/wd

���2�lKl�p:�T4k����R.K��^q�o�����Iܒ򋋑h�l����Ye�[��	R&�Z\�������&��)���ӹ��]]�`K<<<�ߦ�>�L%{�'ZZŠ*��04�¾i�^�G�ِ��G�4W���x�(���]��CB�[����X ���$)i�W�6}������8C�:L��M�=��p^oD:$:��b���#_y�af��Y"&{�5���=�Wg�z��t'�ueccJpM���iB����̈́u���@&�}�##V�;}��^T�+9'�ʒGg�k6��Ӣ�gOP��cʥ6Zq�t�wP�*u�Z��˘���j%�YKK�}�d��ײ�?v,j%i>�T�+u��#��+3Ⱦ.m},��	HuI�{oxS�\\�˟^m\��3E��8Q��Ǐ�4Ю���B��΢�o��AjK!,�u;w���;�.P��k/+o�vF�2�^��*?�L���.y�i��F��J[ہCVb��(���ݽ������zzzF��}��v�t�s�/����7�0Yg3��U�:���:��˫�N�m�K��<�U����C��<.Q.����Vh@�>Kd�.�ۅ��ͫW�)�^��::m��F:�Nk)�ޜe&�o��d�D����6�f��͌q�)��s�]����7�9*(���஘ُ���~���k���R���p~56a��{6T���;�6N�MԬ�,8�sd�)�vd\Ovi��l5���l����)��|	.��t'�����8��eDA��f�vɞ�����~���(M�һ˺�,�5yPR��9&R��H�X��HV�/}���O����R[pƋ�Ykw�o 9�W��CIy�E2�3���L���H�4.�^���[�8;*J���&�)'| *�է����~���g��a|�������n���#�����8�}���y������uK8��~����E	�}Q��N[n[[��P0߃�����3��&�c�����ΎI}SHZ'�mU~ݫ�������w{{���ՏfJqo�|��NE)'���9�أ19����KZ�ݐ��Ϗ�m���������I���C-."����\��q^�5A,\�#�CU"�nr��'{{��{E=��(3��%������k���&�bgP��z)��w>$������ə�76{g)~����e�o|�g��<w��a�	E��3�AG�. ]-c�z�����\�Vc��\�ar�mۼ
q�'������K��'[>QdJ�1`�/I�*��A�H�����*D��l}�ɦ�x������'�"HrZM���#��g�il����+��DB^����h��$5e!�'�8�HY�"߈���
cr�3����Y�������!ȏ��<��|�G��>8����V"�C��m�w��Y0ς��g�P�v���+��,3~�*9�����̩[�M��m,'�W�I}�a���xN��q�_Qݽ�yh'$�Q��%�w��j�!�V������֐�<�Oȳ������iT��ώ�Z*�gx5�+>�()�tZ%��˷��l;L���I!b&����fcc#ˀ��d�Q��#k^Ł�t���3bԓ���6HF��%�L���`:�R.+��A�.Q�n��Ow��(A�C��-���(N �Gcx��f�a�Ҧ����ܪ�t�P��
��N?��NDup�%^z��
:sӠ8t�۰6�����3���~{��b��'N��x�E7��g�K�\&��R��~@�i;Q��yJji{�������a�2��+�=�o���#��t^LW����>~:�¶�:��+���M��r����9����BS�d���iAgϑݿ^�333����6qu,�T��5G6f�}�����<�#��6�WţD�����{�>,�	&������EUe��/�)�+�Eo�����{�'��.ߵ�'��S���#��od��0��AEr��M^�9ff��;\Y�ҭ����P�!�Δ���r�����v9=Ȳu�ֹ�|fI�W���O�Q���0�����dZ;0ԶCW�~�e�p���5��ǹ��6o��}m�y�;�3>(c�I��RA ��D����_�V˫:���������� �H�N7��6�����aߦ�Ƥ|����Ė%�J��0E�_k��:������'�;�Ҝ��y�$�$fL'L����hݮA��#x@��*d�,e��!��v-z�2:]O�k�c^�*0�s��;$U��(���O=��*�]����ia+���䚇�&?��P��J�y��^�'��21+Xȓ�@��Z�:L��΁u��\^N,@c;@;�\��s�`���>2���b�G��i�@SY���v�t-0c8�C�^m���ǼM���u�,�]y~�y"!�2HV�q~�7�����s��du�ė�TDvF���/�g�'�� �n��@9���P�o^3��V�?�>�����;�ȭ6##�D�'��長CXoa�|G�н� ��ܛ��F��L�t�35%^I��S��p,omeg�K�ż����=w<�*j��}��B�
2�H0��}�҆�{@�ަ�����'atd`�@�(�޷gV���x���pn�����/~�Idw��=���W���
���~^�l�wOZ֍"ĉo���>�T �}M��٧b�s��R"�X��4W;�;XXح���ë�G��$���"��N���Og(��)g��7 �?��ӎ��oL�݂>�)7/��5ǒ��{h�C���ƭa���i�y.-~Z�MeJ"n��bc_^^�ʼ��iyц�l����7v�|�_"c0�RUOd�M��c��#�׷]��6�J���6��iY 7 �	!�S���*�$�+����џi�cJ��d������w(�+�e�V��[���uf�S�`���K��}O7?_�}*�H��y`ܶofL`���0��L��8�����
��0i�F������o�5�m��[�A���Iw�&���2R�ե)��z]�e��s5�\�^0��= �CW���j�����)�3�G�l�I�7���s�2��L��9���TW�	8J���;r^MČ]h�5|#��c�����'��镕��כ�5d��ֶ-��(���yQ�ԯ�@��qJ��7�W�����|�����E�Y�E���1����(9�Y1�+2��u_�"��6vVW�ң���s�8�&"%��8_#ެȈ�pp�!���1a5Qv����r�2��� ����ʚ�B���^��iԖ�خ���TUfz��-�_ld?~�y��ધȞU�i .�=�ѾCa�v�J��k/#� �Bd5�����`%zYo>茕���W-����H4�ikG�J��6(R�l�GUd��w�;������nC�+P��=ߎ�q����%���&ɿ��=�VPPRn��.E ڑhy@?���ѱ��$�9�yX䠰�y��v��r��������8��N�`' ���Ԧ�����N�����,"<!�D&Q�l����x�*���#�V��Ľ��
��Y#S=*�ai�R­Kб܏:��V���vj(+�#m�o�P
٫=�r<�,�����������8�.Sx�,i�%Q����*H裳ZՏ7O���k)qw�)�S��܈���RҴ]�G���cC�1��lZj]f◛���:�v=K���w\�3��9��0q�l�7/g!N����.���c9#/�`��Ix>'9������:./�8�����$e�@��EE��}�.�晙��hz���2�s#�h��E��oJJJ��0��
���hX��:�{>�kq�k��2�'��r���g���Q
M�Jp��g��s�i�"�C��c*Csۅ�Yr2~�7��A��3D�6��Gu���)ʃ�q���%rV
�f~��wwl�l��*ۈ�/�޸d�^��/�~��t��rf�E��{��7%|���!��w���Q�Vף���9k�epO�&�[������i/E�����a�	��ab��~ue��6�;�@�d���=NF܆����]s$h�D�o�
;����e��� �r�$��c�]�귦����h�$��#C)������2��պ�D����D#����n$���ׅV)�sD��DI�&�ń�c��[���c������;Z)�3����En� �sމ ���#��oǩ��bG����D:�����r�	��:��{^��hhس�r��]�/��r���s��yA�b�D�o�m��#H�
,r���v{�X��Q1%���1�M������/���!zyˇ�F�f/(ܠ�����T���q��wz���8K��j�)�rv��!��Q�}D���}�}�2�奓�N��%q���Φ��Iw���z�#��?�GNI��"Y�����S���c5m�����5o���fO.�Cg˛�T�zU�FfL~&�]9�)ӃL���d
T��$5=˲��f/@�Fz�vwJ�o���]ϡ�R�cN�_5��{6���+m�8��I����,�O�mɐ���W��(a�Lg�+�4�$�p8��"����Y�:����`0Ky2 ��Lq����fJ��P�7t57���7�.7��%�HK��q.Of�f��W$iq����;:
o����y�>�ϙNxB�	�!�v<��ZZF���͞;�UM�?�Y�?���*b�y5��!ߐ[������hX	QXl/q~���ʹ��0U��<���õ��nkgd\������/�W������.-#3�Z��������C?��H-��y�����84��dī�����W�ń��C)4W���G����&|����S�}16e���s�u��%\_U��_i���W!T�'#��fI�����X�M�FN�d���)mwEj�I:Ӊ�1��-��SQ���ş�8a�`��-x������T+~gA�+G��Bc�T�X):�����}��?�w{x�n�e���o�y{߼�p�ǎ3}\�`c��V?��Ң�@��8"�_�CmC���4�C�f�����[(��r$�:Gi���������Y,I��/&cq�(-z%q̉.�b��E�I�DșY�Zj��2�9�	�;�O#bNMM���ZDv�)������l�탏].n#�۱&��z�uK���D�vE�p�%ox-|N���'�� n{
i�x
� ���>rm�)�^:x�I�{�Nz
��3�	8܍�9& Jv|�Os���U�E���E�ܜ�aSNռ��'�e'�-��8�޳:<ݵ;>;2:�rd�	�>�T��8r�m�8Q��S�d.Q�r�oz�տpr�w�aF����$����� z��ob�ftMLK��p"W�8M�̓1E�Z�\�����[%IG@7�oE�#�,�ܪ�[FNXڅ2���*��Nh�5dD�1`D�ZZ27�QB��K�v��
��kΧ��Ðf��8���[��b �2�7��P*�'�Z��py���98	6R̓��J�`8�B��EAAX�yZ�{w�r���w�r���T�{r��\�f���猖�|�)�U��w�rP�[/�L��hK��|��3J�K�w�m������������.⦵[D�!wĀ�*��9�`̠�I�Y�1����95>���Z�kԐ��T��P��q�nC{��?��{�X���z�}l�Z�PY#��=�JW�F��󣗟�̞L�J���r"�X�c,�������PtL^ų[�{u���˙�t�>�1��O> �����{�R"""5C�t"[x�ۤ��&g!�s��A2i��̮�?�<��d�3������Z@��r����Kl�(}�����[3�3]Z`��sɖ�h��B0�v�%<,b�:����oHH��8��RF��z[�I���?lQ_g=(sX֕p������_�Z��r���!�/��~0�u)�����qQ���`��b2�1?����R_^�w�ɞ���&���L��.�#Q��?O��i�g�4��e#��U�S����=D���9�KR�G�-~��0��׺p��֥����&�؃^�ǧR�s��ۍ1����������tJ)������"�׽�iO�U�WId���.�n�A�\���++r�l�e�}����2Q�=�^��5n]���Ӫtke0��M�{ǧ�������	:z11�ukp9�mK��0&��~ʔ�`˟�J���@C?[h�������ʷ��k;�ϩeťC�9��g ��j[~!�jk�^��OM�tHU��*�	�j-�����)p�Zs����Ru����UQ.$;%�X
Q�i����20U����z_����Y����<վc�~E��V56�=����O�d�@�v�\կ��&�HsԐr���B��$[�����f�`zN�]�:B%�����]�*nA�D�󨬩�mѢ���T44`e]���[q����͐XG�S�[��4��/bb��UO�$�NUk���t	n��8��J���Oͭ��� �i�r�{E�:E����@�J���(üU
����̑��-׮㊑oϪtT@F�>��>�b�\U��� k��eT*�����F�.�-MM�K� ��1:O��[k�� �6�������r�ꗽ/����]]�P�KL����a\-�䴼߷�39��Q���}��o�2��E�h�=g�[O�I��F��k鮿�r��䎕��l
;�� ��6e��@����6��G�ݹ)�j,�^B1|kN�Jm�������!7�j�����B::�7׺+���I�%_���(�U�a~Fs�۹����ݡ���#V�����e�w�������2�hz4u���c�tw�<���n,�E�^|կK�N���q��:_Z�
�0B�}A�O��������,����5������w����3O��Y!�B,���^��B
l[�xk���# b�C�5{�柽 ��a�����FDƒ��m�=z#E}�ܝK���Y9V4��j*ѧm�S�D�]�ss�kY9�)���yy������F����Z�ݿ]8��Q)a`��p��)L��L�h�H���l'"&�/-�N�	��L�%L������vo(*��9"dgggY��}��sō�?NX��^̩e&���>��}�P!V+�%@#��;*�:)*Y��F򘬃�p��-�Iq9�t�K�d�ht�b��#Y�,;�"�vZ�oQO�k��a�~Qr�B"�=UJ���<��b �nk�thzfe�BH˓haa����2�����w��?��vZ��9[���ɡ��إwE9�r/��1%������?er�&ZѺ
��9�/��AΌQ����3��T�k�f��f��Ӎ��'��Y�}K6�\I/��g1��]�=<=�LI'_དྷ	��f�ۆ��R�j°s��Ώ�M�p����P�Ad�f!8:���Yo����̈́{���7�V���.�2'ӭ������~�F��N_Z����� ��8�Az���ôS���0���R�����br��΅��E}���g��/R���5�CS+6�6 5B��@�z��������Xx+�����*����j�zoD���F���� ��'鷱����H_\i}p����]&Cnnn���1��D%E�҂��1��E�d�SԳdr�Q�-X�j�=��G��<i�:����U�"�1�E�)�l�K���{;���S++~l����!��
��\�%����J[���!X�

�kjj��L A�e�Y�sl�%6)b��y������'ꂆ����]���/`B��9�s����"�fCD�)%���>P�rD` L��8�6��R�e��Bs�.���rJd�
����E
WW�W������d|N�#�X��
�@���X�����v�G��Z�嵐j�TC�_��^�qK��x�g�mՔv��D��@�'�#�	��d���\�� ʻ�I%�Յ7K��ʩ|[�-@!q/W�X�Z���G/�:
�HR��z�K�xҒ�K�?<�m���������\߁.gN�h�,6�ե��9-U��[O%�2_�z�Ck�32Vb�?��mZ���\]y�aչ�>W~���d�im��S���J߁�1V`�V6^6W:|�D�g�织9�������y�,԰[�F�YB�~L4s�3�"�N�[���?Al3 �����E����cx �PCԾ��l��e*#9_���J�jQ��i�V�H����g��D&ܰY�A�hR{2��,׆��b��r[)P�a:;����f�<_��+�X���ޕ��ή�k��&��X9�@�ܨ���ZX���7�B^Aܶ�$���!]/��U��v���N�dj]��ir���H�OA�����g��Fhg{���1,�������c�C�@:�n����o�b[��%�3�]��������|��2�]|[��*ȇU���6���"zwO,���y�|��}��� :K=�E�5D��z�v<>nkcHZ9����4�����;��}�����M�����n	�����a�<�h.�܆�6�3���^�1'p���׹+��˧�`�c%|�L`�&	�R��������y�&�Ş�z�w(5/�|����{�U�����жucÄ����^�#��8���ٽ"�*��!驩�bK�ze0`G���Á�l�&PX4\�|kl�j�;$}'XƼ~j}��ኹ�x����������yLҢ�O��㡺�Z�zl�`
 ����+�8�%�猽=�o��|K��uE��
Aӯ��SL!�az�VA��331�[��9� �ޚ�"��#|�T:�Z2'���'���o �	�*�/r��j�;��"o�`�Ժ��T�!D���|���������0AF���-�u �H���r��=���ؔ����xN/݆��y����Q��v�3��a�P���t�H$���_��7,��tzVaF�%�;F��"�������9?���>���g_��BδȬ��2i2���eB�tS�m��w���e�s�7777U��	�����<�'8Ρ��]�S$��7��e����R;����K�QB�{��شt7�]_O�^���1��Rm:IT_�_�KC����]@�u�^,S��d+��s=�n�'.8�����p��_�ǿC�W�����vfh�NwI��^׫G��LlJ�<@�����B�*K�I���Lܭ����y���r�$�Y�Y^u�8��6Ϲ�ܿ�fo��-"����Ƃ裘�>`>^w�ˀ��ǿ��F/V�
���%��Ψ̨[��Y9��_H�y8��,�3��A�?���f��5R�|�!���7p��KM�g_��8RO2U ���g���[d�h�E��jw�
�6�JCfI�[:&�c�Pw����9!��0�,	o|��YuE{��ϷI
�b�M�JN�w�xK�\?,�P�q7�SSr��c��q����v�.%z�o��{����;`-��A����T���q�К'�&B*jK,�R!�۵F������j#%���q�Ԋ���"����(bټ��Z � y?�	�1�<�KN�YYu��uE�`߼�C.�D�r�_�´�ý<,���Dݜ�z�\�k��[A�K�4�q���~��$��[?!�7^z7�4)D�����ǰQPP��4�Raױiyc�(3��^��/�j���/�	��FIb��Ze20��mJ�hY��i��.�*���E*�E֙ˎj 7�	���b6 �c';E�ޕq�����dR���'Q}	@5o��JӪ7g�"|����nv�z���"pB��bhc4��@FA�\덏��.vVff\|����	�|�w�&���ɭ����_����^hh=?�<RT}ȹ�Ps�r��®
(p��Wg���,���A�Yt�HH�m>�¼��4�Rs�B���������^eSЉa]}���d0I�������?�U?X���ak�dŐ��wz0X�3����j�X���z��f�*ذN�oN���� `��ݦ\���U�Y�-����c�B�D�g�o9��(�����ۋs�t,���:�O�%MUQ��3)�����s���Gn�;騣�vc'^�\O�P��0/��FJP%ҭ����	���Uv�z�M~I�c�̲�S��B~���ۑ�L�O�`q!����0��N ���fg���.@:*�`�'�!�,�h�p�r���f	��1~ck5�͜��C�>��,����}#TECt���(�䖫T�u��|�ᦺ�G!B�7��Y���[-Zw���W6'�����>����c��x�k�K��Q�O�
^���X��˘���6y��6��)Њ<��&j�=?���QRS�����Ɛ���	Q���јD��0���M,���2�V���8A��ʞ�@hgA%	݊{� ��W*{�������"6�d����o����Q�сFx�
����r�8��ۮ��s��1��R�3�s>:�WS���@D������u>�b�w��{}�sxWg����_�D�K��pxT�iE�
m�Ne9�3Af�̨͖��K��ya�)�R�۴M�2�CZ?US�@�f$3��M�ĵ`�M�U�D�miiqYn�	���خ\��:�v*�~)��}>;~�|��9��=�u��
Q4-.�9�~��>=���dgfF�{V����5q`��c�M(,K��[�@�0M��������R~a�����ɉ"�@yY�Gي��B�h�'%�7�f��Hp�(��N/xV�]��6�
�٫Y��dO�r5R�KË�L<��rs5�4��|��z����:p��s�A0��?,b�����gOpҡ~|��ǜ�|4rk�@�����k��Gsy@�/��W���<�}�Ank���=N����!�7g볼�t20�= ϛ�F�աwH"z�<�\�<_���{����--����Nxܞw�bE�V��ap~1>�<�C*D�;�j���:�<��3=����ʤ�������sr�3y�.�#�̳����;)����Db�"՝>�c��&�!>1��B�o�þK���.�����Ϟ�h�|�zw&DU�ϴ�u��6����}�����VP�@����$;L����7����5^�b��	
%nыJ�kO�y�t��6S�$q���J��]-�����@�>8�wq\�o��<{x�e����:&�_���T�����Elqԃ'Y�f�����5��yl�L��f�apR(�Y�l��[㗬�� k�+8��)q;{���TYٽ�� s?檂��#��Y�>�����R�$�}3K�6�$��fXb Ҿh`��k��P�'B���\~tjnaA%$D��-�	����k�C̥48wr�1㭓(�r0��ጌ��De�mw����&YG�6�	�(}�Sq�@��G`X�I*r�L��c�Q�a��N��%&-RQ��Π����ȀA����D�Ҫ&�2�ZYi�˷��v���dAfa���ּ���Pga!BOOOqIɡ[��2F��f��k��aR3�A���0B����@��\�*|ٖ��EP���C�j��R�Q,)�q�]���wQ�O	7�L?}��D��!�wO�o�@�}/�e����.��$:p� ���{u��Ye.C]HaR�
rJo��V�>�v�oUGM��=f���n�q^>��b,�x(���,��`��O�:�0<:�����uHS������y��W�!=���[�S
6%��g�F���">��`�l!5r,
��HT��]]�s�=��W%*9���O�4�G�_9$��[��(�>|�+�0i���s� �i�M2��yO���{h>�G��fM�lk����	�F@�CU���6:�
�N	?��5����B/Q��f뼅u�zj�P���$;�0Had���d+&n~h�[�ݟ���W�I-��$Oc�W�8����>R:���P��_P�39{�:�%8d��O. ��栦����Lu�Y���VBI	��#؇U�5�<hM
�� m���W^�4qI�8rr�Y�l���f�$��nB�].�S,WV���_UW�~��������~)**J�����������WqiE��!N��#B�qT������X��d.���
�w����g�r��(�q\�GN�����?�,�������0������\{���~1�������$�E��?h�}��I��ZA� ?��JB��{��塞�+8���m�P#Qs!��=z%�ɣ64��l��e��Ĝ�[�Z���($ia���a����� #��2^�D�u������RF���"������B%�_&|o=[ܤ����ll3;Z|�4�L9;��,�����%Ajͻ��o3ۊ[���<�:�^��}�dd�ϙK�G�6a�%b���rg�(7p��j��'�	x�/��KΓ��!�s�`���-P�ѯ�oo���l�w�qB��������+��w�֣>�B��Z���`����_��iLf	��Đ	*ۄ`I Q/�����B^��&'�=�e����:��w�n6��nJ�*�)5����� �{��*BvC�ʾ�;��M�.�Ce:�d�_h��E=<<��5񷹜+Q}���F%MG�ܭ�nj��=���$��$bk���F�<	ɞ�C_�P�~�������ț��đ)��|�������ѽ�+g�����������^b�PB�A �l�)��82���*P�$�G���4Ρ���������-�'(8��`�w���\x@KS��[��sr�����FQ�2�J���*)�sU��d��2f��!�wL��M����<�Y�c�x����f����f�y^i���o���L>���	)������:"wtt�h��u��� Ỵ8s���ֳo�[-�Z.����G���Y�=-�N����DP�	��̭}��4��>�Mf�nl��:yu������*��A^���9m��i�F�o�����-Oݦ�3ך)��2�X�m>Of�r4Y�J{���H��A����c��Uà�y���n��Acr�+@�l��L���㋡����K`'�7���vv�#5Oo�[�ߚ=/�^u&�]�C�y8{N�\�(�����
ǆ��r�7т7���&���9�s3R���0�;]���63���C9^7��A:G�Z1����#��o�&g�;8(�~ދ�il������-T�g�����F+�1]dE��ٹ^��`�?^���o}��l��<����ײ�P#!~��ܧ��I(((�)������:7�\g�WS���/F��2R���l%�����ۧ��6��.������idc��C�[�ǳ�h��'�P�W�C<����0��Ѵ�a�`�E�o��*�h��8\�|���E�f639y�����-so__|JJ������7��8�:|R�#�����C�GQ�J����JK��R��g�}�M��Wr������3�+�Q�]�
��MO́�n��?�X<� RXUdN���tk�����hRàuf4#���GE�����q���7<s��eƊ?1rw��J�bU�^�}o����9��-HoZ�?~��+L����Orl�d@�����Bkx}�I)����z�"��A�����_�N���w�-�7���!��N?b^���y1���ݓ�*�.��-34�`���Y]�N���7��;�f��y%���R3"�j�%r����~ծr^����~N�J{FFF��h�x���+��w�{���!����9-HOO���4*ԙ� I�fC��{��Dtu��k~�60�wW��Ӊ���4�7K�|2 ���:�_S���م�R�(TS@�g�ki�tx綴h�C���/��0)3�]�֡����>�w;���T4�^�F"s��n��4��wcp_��.O�Wr��U����bӨ�/�b� ��!jѦ �y�hjjjLf�XcH�+{��!��T	��z!��#$����*��]~���*P{iYw�H>�+Q��w������Z��;�U���,�E���^�O���0�MH����Q
����������>7g=���硖�顀�;N��$�����Y[[W75Y�o�|����"5���u�C���_)ykEui�u��S��X�^3>n�Bma�[FW�
3s�3D�	�gz�4��f(�b(�����rMMM�7�A	�����p�P�4��_�8@�6�.������Ɛ����6�����I��s+1�Cq�PZ�+���j��NM�w=���{Zv�&~�J,J�����HnCJ���t�P`�A�(��������aѠ��tU{]��0�����vo��o�5�3��s�`�\���$pM���Q��ܼRX���kڐ�6�,4�2PX1�>����~������������p�wxx�	T$�o���R!߼|B�bd`���ٙ�Ċ\~y�f��~�'��-�]a����	TE�h]�����6<:<dץ�.d��]P�q�5}��jr��X�4�~�q>H�������u�8Z���F�Ĕ��j�<��Pb!�m���(K>~ԙ�OEĉ@FFF<t��ݚRT[�7��c���w����S򅞎�Pw�3��R�}���s��P����^MCmV��?�����126�9�;^���8�����X�/���ֽq��{ 	x|~��k�eM1}�� �v���I��cԊ��J嫺���z���qUՐݬ�Zx�͆]����.�fA֤��Ջ,L]L�]��J�b��O�,:�H�����͗Հ �����dl����w	��'ݭ���1X���s��\�Mè?JY#E�O��:���?GU�ry��Q-@�g>��ͭY������ca��qus�rq�����-,�ȈL-�P0C��󌾥X������O��K����a�3��9����D���7�̳|�8ޮ�z���0St�x�j�V���g'"V���V.�/��c��+Z���n<�tdY^���|]�_������P|�c�P1Xg=����G:�xS\��Tw�~�u�1~$TB�v�o f`)c�*��3�����������T�sҋ��k�V���݁��V��P|�j�sfZ��"]��j��]]9�����f�����Ì�&��+���	���G��w��6Q&)h�����?������>n߸nYM:H�-�762G*�R44ֿ�lS�^<��h�˚�䀰�++���[Xّ���hY��Q�]݌�����}�`;;;'����|�<���/tFe<�
�����0��a�O㦡����`���q��M�Ʌ'E�Ou�ג9�
ֲ
ۘ�p�՗�++�M~�:D!���6952�mX�QpIW�_V�0����s\�~ү�E�o6|�M����Ags���~[�z\x\ە�x0'(��7]/��>-ܜnt��.�OL(�Fwe��$<�]�&)D�(mMo��##�1;A�!���;�=^,���o����R"%4��#л<��l黆�A�$���j٠�����%ñ�2 �9-'������^�����������~����n(���1�(�Zu��Q�>Λ�Z�����3?3�<��to܍�u'>�tuB�&���:먪���@P���n�VRBZ@�AB�Sii����N	�~׾�߽��c��sv�5�3?ϊ��2��6C�$*�����u�����	Ɖ��^tC���̚~i>ס�i~ƽ�����9y�ZB�zC�J��,z:��<�yT�� I��)]��z_,�����k�!Hb��3F��Sut~��4߶����ׁ8Jܜ�:�yTΓ-L��+�6Gk�.U5BM%9>eZ,���g��1H3|ښ	����<$G;��%-��f��k��<�#�j?,��.��ǟ�5R������Z:R�ۻj`�"Ow�k�˝�t{Uz����9�A=SM����q��B�l�g��gs����		���y��,���цTTU=���<-���IR��ʙ��>������$���J]V�����)/�^��۝�V�x�72�����06G< {h_�M�T'5��8@���\T�˹�Ë�ó�s:������83���"c<���V���B�ߨ\	����&
�#
�W^�i2fj8S�W�	����\��> �p����"c!��'�HhbV��'��lH�\�����-��;�	�����C�CT�E����Գܵ\β�*c�)mmckk�7X�
���U�������a��ء��_^?WAqT�MQ=�*���+��r��O���u�kH�dd�z���Y���7���]��9��'Ő�&��#=Á��I�F��;n�z�]�PZ\��C��u�7]�˿\<m���e�[�����VCf^U�=�!y�L�Iaoimݵ�����.
�ߐ�`������GPV�ON9�)G؛*P��5�^=&�ᓏǕ��Rb,��:��P��]� y��jB�U�{�t^ۺ�!��&�ǰ󍆣A�F���880 l�އ.��'��%����������X~��q�:��E@�m2�b-�k�b
d���e��[Ͼ�i�x;��/�b��;�����n��Ul���X�m�;��7�%zQ1���^�bC���K}h�gT`jx}k8U\B��_�Bj���^�z����F.�6u�/'�v>Q�֨@��Z^^�T�Y��  .!ij��S^\LV����!�bY�����Qc(e���m�\�B���wq�T�7BD��q�g+$���n��������
��b.q��Q����R��ȅ���Q�?�7���������()� ^QQ?EěX<ݔ���TFq9�p�����<y��\+ß�_�m,��*��B��o�ޘ�M�9��(�A�d�v#)o,���
�Fb��6��/_�toF^�N�ĢÐ0�?��j���M�܇�d�[����旒��"q�z�x�73?�ihh�Vo�9~zNV�&r~���ʻ�7�Q�?^� i��yy{�����3e������w]�=�7���Wo���qƣ<�TL�����D ��C#�I�YQSӃ���B�GI�f�J�绲����\r�b$���@�RΤG|vφ��
��VTT������*ES�W	�$'/Q��š˨��u=�����t{Nf�������h�cb�˒����#K�݉���<5Ff�5�Dj�>��G~�d�I9����6��� ��w�h�b`J��A�*T��q����쾛O��$奵=C�����X�a�u���ln���%*�ibbb�!��fI����:u~+���-Ш�ZO�L�{��c����f�&�j�?��"���S2!0��'2��І�0�SEnS&��=�����3Ly\���'t��Z]52155<���|2S���m����H��ϟU�#Cl�R�X�7bF%V?�^CK� @]e�^�~�������)2�`4T��Ȟ�1/�D���s-VD��s)���V�;j�Z��ֈ���D	�842ۘ�YC��Do��	�" ������,����IFV�ڔ*�zw�4��'��QYbT[N�������Nvvzq�\<v�NКi��W���S���o^7�R���(Va�}�I
�O���MYi6���I���~��l���%���F�ʪp���c.]{�
�ί��t���;�� $����2�Uu�9A��؟�������J�;<"���t�r;B#(7Be����E�.�S��1%�����'{����lz�'&�LLL,ȖF�ۆ���ҥ��߽b7t���PlkϜ&$�����3�[��k����|�<�࿸A-nh �.��͐7�0|��M�rx5��(�?q�+(����(�	��l��q�����!A��&Ǒ.s1�foE�����J��� HL�ӳQ�b�=����#S ��0��=@���Bv؞���P�A;����
"���IK3j�L����eU�hL;2c*������?��<����ZWT��&{h��`�ܯqj����Vd)cbb��V�B$��.�%%A��ٯ>��Ҫ�,-��ЎZ��Ec�0�U�����r�G'kbk�,�Fty���{���8��=��ޞs���'̫C�@U�A�}��E��c�k.111L�~�*��'�UW��C�����-��K�w*������,�p��R���pFIK�0v�%��E�5��5�����e����F��V�P!��os������m,�V/������R����g��~�W�����)���0�ז<�B]PP0���1�yEE;>��;Rk�"��
p2(<ap�d��Zn��� ���#em�M�OLM�h�{1O G �9�.�U�U&Wx�G1�Kln�������%;:i��<��]�w���i�'D�3�r��IJ"��ĳq��O!�oEH=�L5���i�#���W�h�D��\�}�N���Z_7 V��|=L���ӕ��m��-'5z�f�尌��I�j�:*2,��%�f������3ƸYT��i7�Npͻ*�Ϳ|$�;����u����w�v0��齓t��'�휨K�'B�MB�s9�Hv�'DD�A�\�h.~�h�x�$1��4�� �>�Mw��x/������W���V�������̴����>)����\��s�g��z��f��?G�	V����Yf�&���`
���A�!w�Ro��U��p� $�ICS�K��&"�]k�?0u꼤}�ccq\�g>FSK/p���Ac%�7�$խ�Z`e2%���Y��������g���y�Ch�$refRKE���H�ip�)��{�]�s"R"�(��Kǧ�o2Q.#�Q�ЩX��;^�ct�B�e���Uh�#����u ���?�P�s0�wtvBu�toz$o���,M��a$hM��o6�+v�^E�`ٷXՖMH�1�?�iZ��Ê#)�9�ﴪ,>�?�H��l� ���-G t�P8(4���9��7)IX�3�q2�˼����^�v�=O��;r�|
��(Fp�H��~�*
��;$%Ɯ�+k�����9���A�G��N��FR	�}��e�1��9�hm[�xjl�Э��2{�|� ]tG��-�BD��	ֈ��H���,.�y|�ѱox�w�!P��SZ��e/�/�Yu�.�,N	ie-�����@��VECP�_[F��ճ���x@6T@�7��� l�~��Ȼ����
��QN�7�9}��t�y�sxz� z'yrr�h/��0��й<P��c���T�c���AN��K )��p*JDOY�0�tO�����P��Z�O &��=�KPJG��]�6"2��p���[����z�����@|�{]�<���i�m<%9�DX���ϡ�u��n�kN&p���# ��XY��5��vt6CJL��#ŏ�%�J)8W�Q\T����'K�xz�& ��$n����yM���"аq�??�f�����j+���F+44I5��S5���d��c�]V:S]�0�Զ����=}z���j(�W�P�����b��!�T�kQVV֣���d���'
ޢ�����T8�ZA����r4��bR
8�eФ9o�;&'�����W��TT�K�[#A�����5��}�y�rÚ��Z]c3S��&�}�K�|_�󼭻�;��\(�Z��	�#��c/���X9��d����8�z��O��yc����J�O����Zܱ�O�>mB�%:�p��6	�O�l ������(�<ք>�W�yj9�M��f��RR�M�ͩh�5�5��*d�LL��~��9�W������}ZJ�Ûjnn���rt2�1>����p����R�Cc@O��Y������Նgb���g�n��7�k���Ez�ZVsM�'G��MG�"�\T��Yh�^����L��HZiu��\����T���Y�m�j�|�roo�H��0Q��(|o)߿QWW'�wxM�HEUn�C��CI�H���oݛ�{H��ttt.�(�����4���Zm	_���ȧ
����tC��V���B��\öN͑=��.���R7���h�5�I6�Q��\�t1�e{�0VR>>-2k	~���s4Ɨ�/D�5�����K�A�;%1��JG(ѩ�^��|�~��L'��fQ�&��k��3݆{�*�<�O:��g�ڇ\HHH=z�yp���:׃A3�hrll죥�{�/��M߅=wuޖ{߸��b4Ƀ�����Az���E }Q-k��ɠ���F�E7�)p
L<��4���e3A�#�͂��v�]Oɨ�`a)+,4>�V��Վd�C��͆�I��s�[�GH-O̾��ռ��?m�	��~5Bޫ_F喦<�"**�S)œ?�Ц���(r%q`���oŠRW��G0�{�D2QR����o�s���8����+<Q��61/���6��E��sxrq0Ps$�H���ąT��a�;����Iw���FW[�V2N�A�˨�VA�s��Ç���n�=S��0R�9v�7w�u�r�̤{��]�D��DP�N�1qq�}���x? �˧;�y��-��j�*����3u���#�����׺Bq@����ځG',L�}}mb9I&���~y:��,�u�B6M}��Gy���i�����Է��D�6K�/X>�Q�V������(���2AM�̌������7�'��?��:kV����k�˸~��mm�����m�Zh�h�jl�J}�P888���vW��=X��ېtN�\N&$��4:���E�=�a��h���l��sgH�� �5�H U�����G��խ�q��{O���CNn��FYY����!	�!��;+�>Ћ������!Y�֕9n)�F��;L�wD��a�C$�&-����TΔ�XjN��[og������E�1�������
���|����4�MbO���~�ooϔSCTU�ո���_v�����'��v�DTT/�gʍ!�H�`�4��A0����h|,P{�.t�K��\~y"�5h���aK��'�"��d�}xxx��v�%o�19ܙq6��H`��������8/�L��XX� ��QL���/�}La	<1d��#J��S>{���E�:y���e��c���j����BB�T@ Q�5�]� i�����'Q!R>-��0�OL=f�)��9�W�y�ٍ{P��Ut����IB��?���ڻ�e��c�0�åZ�?�	��l��f�6Ow���X�m�3���a�k��y/���
��E�=��?��i681���
��ְY^'��<L�@�9��t^��+]��be��g
Q�=���@ĩR�(��Ϩ��  �V;l�������؈����k|u�WJ���#p�]_T?_�};�z��=�-��Jid�XkJz������#���Q�k�u�#�7:&������4�6��@�o�1��S^;K�G;�uM2Z�o������
hR�~+���h���m�˛h`�v����8_q�bZ���#�g�q�>���ߑ��R��wގ���߿�)�O���N|�r'��n.�=W�g+c>K�X���a�.�;N\K�T��7}�ح���{� �%O��gum-������12�����.p��{_�@�h'\dD�����W'ǳ�iDBS�w��/$�1�Y�k���	ΈA�e����g��#�Hٴ8�����{d&�?�rz@|Y���V�T�V$$T�ԋ�k�g?e�}���z��ǫ��5��i#���Z���j�^��4l4\�>�āv�~X��sK1�ާ't�]�	�TF��Ǩ���a���,ED�m��:k��qg�	*���O��.��T ^󘙘<o��e�^lz����e��U2�{tp��d� �@Z�}�;�
�h�5��{�H������=SE��c��ot=�4:�2C5ZH�̌�g�v�7�A�z�fh����C�#� �9�}\l�+�����+����<�h�:��7�<[��@A�"sX�;�L���9�֡�k=�N�"p�����kQH�'�m��O�R��|n�2l!
͕�*&������|���ϟ?;�n@�B��c8tHW&�Љ��B��?��},���#
ߋ����-�<������(�́{��A�v�CC���qI���p��1���~����K�*�O�O7ہ�g�Y��'�ז>����T����$B���t
^~rn���
��0�fO��kۛxˑ�ZQQ��Z�W�¾���h'7����uGh޶�8 �_�����zep@�J���^��]
[�.�tpx��QR��v6O9����P��+D2P��@K���Z6��E���V\����S�ZA���ؔ�0�-����$sϝ����Z:r�7>	I���.����Y`:�.67���gT�[.�oi��LM������J�T��
Ƅלd-i$���4"�S\<!�p�303�]X�����<U��/����P�Q o��q2v�80��P���J@-�DTHH�9�� ���-��KR��L�
��R]rhw8�`3��D������V� ��SEL�B{�L�� O�оae9���qL�]!X	"�YUm�br���2�����VV������|P-��ι���\�R�TD��ӧO��Un��})X���.�:��D�.�P��t�AS��ub@�U5�
������[q����t�ETs$~LՀT��y���$.s���������!p{�K��" _����m�V�^�3ӐA��'�C�e�M1�+�
%�LU�lബ�;}7�bheu�7��6�m-�k�w�84\QL~�Z&'�J0[%T���p,K&Fob����\����^��@�m͍f�9�g@�	�Y\\��X�&!�$`E�4q�t��A[�G��i�9I�?t-��x�vdTS�mGV8�s���&%�c��O��.3��ڦ� � �¾�q���OJʌ�ge����^���21��_Q+GZ'���S����U'%��F+�	����;KϟQ=���I��̊\���xz�����(Λ�YtX�F)����`
?����˻�3��ٹ9j꺍.,,'8��j�qzs���3�A��Ǆ��i�)��=��m꧓�$��L8gk��X���Ȉ4(��C ��b�s��͹aMLqy�J>�Ӷ���J0�6h�Y��R�b����|�LWs�D��);�*�)����L2F���R���∸EN����s���Ǹ�1���4����bƾ$[-����ﳛ�az]��j����JX���ܣx�)|��HX�X��L6-���t�>�旴46@��~p��L�����""����q"�W�s��e�;���UUT`# �b����e�&ll9 �?Za*7���c��`����\���d��"����kX�h��՛�;r���P�G���贴R�MPF�D9͇'�:{{����:�vC[㶼��?���X�(p���]�㲜x�V��V-O)}f�uF97r}���Ɔe��f<'�h�|��d퇅���[_`DS@����0$b��������S��V
ؼ�j�~Q<d�seƹ9�3M=�
�����<5��y�k�O�>Ixx4��e``0���/����G��L���i]t�����l��Cש01ȅ0���:��o�g(�K ��&$de�f}�vvv�ӱ�"$�8��;*g�>quu�쩨�%HLL�Z
ڭ.�@s����NqrsO���ؙ��<�NQ�����ػ<��uޝi�n܏� 9@�d��ɖ�"�bd�ݺ�T���,�=W[ZVQsw���]p�����?���ÇKKT(m���j0�����t 7p���b�1ŀ���A2���!_�^,�-$4��Ƹ�f�G���f����),�i�0??(u�=Ĝf��5)��>��$e�|06��*�A�xp�X�]�?�5gLl��p>�� ��d�����v�V�q��GC��������������57�[@�z��������'%����8��N�Kt�h��3i�~��wN�%Q��XևJ��Vt�u?	任#E2�U����(p��ֳ؞^l��\�o��4��*Ju�&4{#�Ɖ���z=�G�"�a+kk��9����9����mV��0�;�rs��
��TQ�mq���ؘS䟝��� �NvTj���B:������%�A�����?D���f od�9��
�I��U����T��m��'��<`́�t��� ��|��g7�Bo�u<�Y�5�k�Ĩ^D�U��%G!�H��}ɹ>-mX�q��5HP��gH��� ��+��x���ж<f�۱Qj9��gz" ��m�Svtt�]kQ���J#�u��8�r� ��U*�X��g?���җ2�,��}����4F�k�q�8�r3��Tk/�9��0TT||�]���3Ɖ@ͦJt�W�O�aY����>��ҙ��������0jv옟��06N�� �w�ޭ�Dy����ս�V|�H��D���YYYO��R�w0���2�����R���G��	����p��ƈ���ϟ'����M��W�lY�TŮ&y	� ��DB>�2o�3��#����8�O�+"�u��a�z-���$d�*	��Ј�Z��H����
����hdl,wˁ#"�yN�U��
�O8���N��C;��.�$L�j�otu[��t���@�}��)	ʕ���ܾ�

�r��h��9Ȉr�~l��#��_���|���rw����Mӊd蔩�(��T5�NB@�{��b�'P�qHН����2�T�z;� rlc��`�������ت9�n�e��r�E�gA������txL글�.8w/��^prv;�4�/�=g��B�m����z��֖���C6����1=w��7{��� �X�=J��h���Ǽ��W��L�c��#}��%r��v��NM-�ond%%%v��PѨ��Z_FK�4::����***��>�A���%���It||0�.�"�ll�8䚚%z\;�O���)))�k���@�'���Ne���0��9�����Xx♣~W_�`C����_�]�ݮ��5��rpPRmz*f�}��mg,�rK�!�Z��*�u�[��qX�I��fCI���^�ǽЀ3)��b+h	�����zȩ��M�7��de=�����b<U��dD� ��d~W[Ż���������_������ݽ2�)-��m~^g4
�8r�,����e��J�J�*�"'z�9v'����h.�8<�Ɛ�������ue��D1`��I�{�8� �:��0���m�:����*ϊ����ׯ1��M��?�,���/���N���Ӻ���%z�Y_
���CHH�/�����T� �:N����?e��o���WA#�����cU�y��"{��]w����X���L�D���������Cz��ϟ�,7�-x�4���M��Ō^R��n��+��WˏI�z�|�ƪ���FB8r_�3�u�#��ᝉ	5Cc�o(�����|  Q4>�X"��&,Ek���sk薥ӕB@����	]��߃���� �Y��{wZ&�%;:2f��w�*G�c�L[G`����}ɶ-bbb&i*o���P�h=-�p3����Tcd�`�sF���Cq Ȉ^�Y�D�4���{�y������B9�������l�'N�7�gq��"�`ۧ�L�'+l�*�
�>�� �YYY���8u{���E��"6�]xey�@@�@l_��.�A'z� R��(��y2��,&V������$�V�=���X88Ԯ2�W'[�\(��s�t��o�����f�])%L���R�<�r��-/?�$c*ѩ��H�3��j�F&8����`��T�-4��ڥucX-�	���O����M�UH]����@e�f%����`TA�4=qD�L���������xn��ۘ���ѻ� �ZZZ���P����-�:���C���jJ�<-?:��Vp�|1�F��ˁ�����?��3��wtz*�xRC߾\HXRR�h 4"����"
�2�s�xI	l���ˍx�����9;E�����V��ݞ��*2���r[~~[����Y��DV)�f�R4b�6�4o$ʀ�<dD�����7�����1�j�3MW/�2+�	����s;z��N���� !����`R-�zgbjJ���#���Ֆ�К3���*>���Ԇ�n��	�>��ۚl愋h1]��Ya
H1�&bH�����!^�+]u�<���;�E��n�s�sc�b�]~|LSǝ;�,���Aye qsGȮAwWۙQN��@�mm���\��f:ހ,Lʮ�Jڶ笭�f|���y��}\���U�-��K-@7��bC����%L�a)�n���kז�/�T�G�����055��K�øu���x���`F�Y���L9�-�f�x�f�nt���]mU�F��$��9��o�����Qb��Hhر�o����}��L Ĝ��&⭵���&��n"_���͸�h�FK����.��vveи����ߚ������H�6?8(�zzvo[��멿1������͎�ۢT&�;B�JL������d�%;�R
8?P��;�| !p����11����E�1���˂+c����[�Od@��!~*˒z���Ǟ�A��B��$�'���')km$�[nK�����ڳ���m������szfg���⁞�{��&hP"�A������3�N���JeB��@�͔���w���'����_a/dy��a.p�(m�S��c��?z2 b������	l��d^SS���z`Ʃ�'ZQQ
@�����>�lz��Y� H.��P~����GZ�D�i�W�x�y��O$��V���
���'ٽ�����l��ydٷ���%�^��`�@�Z>��D������pM���ё�N�ޛd�����0=�G�blG_4�r�b�����HXX���Q�7��O����*�ith�td���e��%����S��z��ɳ��F!�,����l���
Q?3�'�Әz�~a�k\CC�'((L�f���д��8���^�~���r�: ��*�jj��DD�L%τ�HA=wqq	��0� �-�g�����$x�j/AW��k���4�&���횓������.����$R���$*jT��m ��6���.#�V�N$fͲ�Vs�������ih�$eUz��z#!��(!%E��6�FpJGA����N��	��sa��K(�����Ѡ��xx�s���TT�=���]ًp�En�)��>!�mņ�G���G(��%=��	����L�@��^�梃f:�mU
����0jh7+)))�%b�' rMMM J�@�@2)N�>R��DNA������sJ���>�ҙ��_�(�F�aűj�NY��Z�'	@	�p���Ɔ�B���W�Д����ȽQ�ē���{>����KQ ���$83~c�g��I��uY�4����H�4��]$���*�zr��&���d� |�o�_/	��x{{�A{;U�]ݢ�S]cc&��<�L$�����O��r;���^櫉e���XN� �v}� {��O������׎EYl����$�[})���A���U�:�8�i�l#r �x�ݰx�Ro�IQv�;���1ɩs`�����7�����O���8?��WW��^`K('�wڈ�bm�T�����;`�3+�_*
,--�9;�_�����l���ࠗ�#��MC~=V�@p�3�rk��,����>,����ɞ�d�%YM��ь��ڈ��8+�7Ō�KLL����z5M��5��:��6�|N5l�5��7HHH����把��</>@�Yjr�P��{|��3��N&v ���M_W����!ъ�J�n���R�10�z1�s?���u�6��i!��25_^^�!�LKQȥ�����bTlO� ��g{�����%�k@�XPa:??��8�
q����;c4�i�����CX�{P�VϦ���H��͏�"GHer*��}ߞ����k��i���=��_&�0q%������%$��/�(���-�7�����z5������vL���a5�\/G��
\�h��/��@n�����ch�j�`���㵐�pq11��B�����j�Zx |�JKټ��~��;EF��!r��p+ZE|�����1:�ɆveA+1kl���Ek�����#"ЀQ��n5]����)�[ZH���[��V�G���!n˥�k`�B���c{)��2��(�la	-m�X�9�~0ܔ>�V�^�:�X���F��S��=�!ͭ���l��ё�!o��9��X��c`V�F8����C��ߎ�x�/���-�l}k+�~�gGW\Y�N�{dD�<Oƛ'F��Sxx���5;����w�Mh�k���?�Q��P�кA���Q�����t��|qJpF�fA�Аp���]�q�x *U��\M��I��3	I�tϋ�'��1&B�r8ΐG�P^j��MJe�Y)��C�?B����
	�f���o ��Z��]쒜u�&7,�bQ3����OQr�D�
����>P��~s��+49�`'3n����'���1�NP�c�s��s2R�ez0��z|�W)�w�NO^��`�$/��@��.���V�׳�Y 4���x��<W/�ɯ�3_�ȶ`�����j��S�"	�3����g����(ݤ��G�{.b��
D��W i����]��Nw?ٴst�W��D��*�)֮�;�V�m�GL	utrr8������퍇-�h���GG{{z�7hh{5��T$i�H���r�`�Ϟ:��zh@H���i��O(������@�B�nY���71	p��d��ON��_V^�T�Ғqum-:>�N�����������?F-���q��QL���������1�?�})����b�C}|�#����F�"8v��)��JmA�w�40
�Tnq��;Ծ���a-�\j��+
��O~����Y�8���!��vq�q�"��lE��� �Oo����Ky��×����tt�º7�2(A%���V���g�"��1�|a�@[L�HLP��D�-�Z�~|j���e�XX2�H~��	�w�M�J�:�X��aHpyt��M���/#C�8��iJDr�<��#D��2X�ߩ�_#�	�j�g0^��򫑃������v�����%���`��e���D�S4鬰%��6�E���;�����������iL���w��&q�)�Gp}���� ��͍�#,�!��˛6~���$����~�Y<����{���1�a�q�r�F���YI��B�MF�%�[�Ǘ~��l0��{&��ˌ~L0VћCX�:s�v)������CR���d/S���%��=���ˉJ	��7��Tc8$j�jR�֚i��OFN~W��'4�����N7`�ںa�����v�p`�C�ۄ�s�a9���X3ק���!��`�ĽVy��ؙ-fRm���CFRA�D����PK   �EX?��O�o  �o  /   images/ffe61187-e64a-4024-8cee-95dd034d2257.png -@ҿ�PNG

   IHDR   d   �   ��z   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  opIDATx��}`���ݽ&�ԛe˽�;lӻ�5���P�$$��z�!�)�1��ƽɲlKV�~����۽��tw�-������v�yS߼y��:���?����V���O�q�J=~��g
~F��1:8l�p�	�1�A~.��"8�� ��W��b�l���@���s3h������az?zz� �S�?���r��=�|��@e=֑#��!� 7/��j�����3���7�,zz�-���	�+pЫ��p���Ҥ�~�c�͢�ഡ���g�dE��I�7�~?�=���
�dQ���i�9�XY��o����&g���QD&@~푱���(�`�$&�.��긌�O%4<����ϴ���2]���/��h���0�=�Ֆ�ȴl�}=CI�cJ�3��6�	+������ޫ+����~W����YPS�"6�5�pwց�*�F��S��t��e|���VI ����XY|^�������g�}hh��>��|,�
��}0 IAB�P�$BN�vR�JP�]P��Q��>K*`�M`
-Ha��Gp�"r�2ɪ�}3�p�7�O�A��{�;.��,��(2km䢸`���b�	���Q" �o���Or�@�ߤ����z>�i�g��B}36�"!\��@��U#-T�15��%�CH��N��&�q4�wkJ����~s�#1���§W5¨,�M���@�f㳼��e^8�7\�0lLU��5�T���F8g���V����E�L��ϧ�a�����SjC,�ק���1VUd�&�{��	ɦ*�M*{^|N�>���=5.�}��T��Ќ�B�.���VH����7@�dO�P�n5�]�Y���9cݰPl�s�I�N�^	�y��3d�� ����ۀU&���<��� f��ŵb���\����b�"_�T�}���p�>A��gnY~ %&+��=���³V��ML|Ρ��}�GU�c��j%�=|T6�BiU)>�ϝc���-�@�;�ꏽ($QPg�)�7�>�^��Qn�g��Z�o����\p�;�6��(�� }�k~����� *��2�e��������Z�ʄØ+	�����g���{��E��c�2�c*��)�-W��A�}p�0�2HC�7@�/��&���f:T�>H,��Ud���c�
<6���}�^�d�FG/d�	����W$�~|�����Zdܺ*}i}�Ow�p|��/&\�����[���D5̝��������lcO��x�Y�>ϭ*wa���h#�q�@�e��<>��Y#��$*��[�����'�破Q�X<��2TRˑk��
�[�HV`j�~�5A��Ӳ=�G�z� h���ށ��;�f|��	2�6ݩ���u" �pq�l)4��! ��OH}Ы�{q��ע)3��H½���Y~P�gB"9.d���^D���4a��Q��u���U%PPsI)��a������AZ�(�I���EC 9F%��ټ�E�g$ꞟ��zGX1pS�8Be�^e8���w#{�!�l�a�7^��D���a��� \�%�J7�w�]�$c�_m�Fl�����ή2	����>w\i}5���'�Ҹg�܀>B�ۡ�c>��d7ͭM�&b�F1@�O��ᶩN4�;Ψ:��-m��V@�(pKN�����
�K{?��F�	B����27�B�lwGO��r�A�������&:�������bl�%C2=[m݄�g��'�ɲ���@vU$�Pw�N3M�U4��F~��$��Qj�CjV?~�'�h�&�/w��MBX+KDMi4���ê5(� #F�뮹|(*e��#�R�$���s��;���9�g�Yg�����~L/5�;+ެ�E=Q�).�O?\��hdX�o����_^i�����h����L����a_���)��K�n���ݑsF�/E�/lB��S;h�7��T�;p>*����o;"i�mP��+*�j���B��|عs/2"�8x�b,fHMM�:�[�&ޯ��������?*Z��0|�`N�����a���J��>En���N��6�U��0�G{���<�ѻ�/_W��Cv( {���wyF(A���� )k���dp%'ˋe����jQ����n�'$Ҋ<�TH�����RB���_��u�Lbl��*(�?���|d����Ñ��Px����W�����X������U�a���p�ݷ���'�ۊCF8�&@�	���*s���'���4����Em��^����:��Ҽ�V�A�`�­�֡�V.���Y������K��)\�%����kVc�-��<��o6^>�w�q�x��8-����$''�����M��$Z��=�E��y�^M�5t�4��H\ѳ�+�����Oq0g��sI5D���W�wz7�b��@��#�c9N"�W�8[S� �D&�cU��CB��P�Wz\ቂ�����&�=�ڹCE�'g	��n*JZ��EV�Fl��^�.��<HII�%K~��*��\�������l>]�5���~p�/Eb����s-�8A�P}2���N�S�i
��b_��8��
�\��;,���V�%h�]o�o�F3ģ���?�X��E��2F0>�ǫ*F4{��2@;�l"R���_��o㠰G�<�&�ڈ�3��f��,��d�F�4�l���#�N�1��b��Ǖ�r����l<[������0W���C�9hP8���8����k���A.:�<$z}���Dp5*���m��}t��w���j�#�����&QE����hxB���+S�`rl}G�þP$��N��;��I�GUP�A�x�����l�/cQ]L:͐WQ�GG��/���E{�p�8�A�O<:V����"|�r�k$��.D FP�D"+>�
7\G�ǟ~&$Tn�����⪶��#8TlQ4��=���87T�H�K.>���p���g��A	���D����n8k���H&py��
�p��)0{�P�);�M�����ol.���	���a�K�o����u>����U���<D�k�WUoC�����Xm��mHe?�>UpbL��?7�C��獛	ŵ��5Qƴ�����?
�`j	���&M8z,�"�qDY���e"��'Z� �VyME-�K��MLM��@;�*�=R��=QA�e���M?�,�^6��>�l��XZ����s)�"2�A��sƞ���?�qО9�$�j�r@���q�$5'
;e��:�D�I�d!9�tq`��U���r���D3���K�Ez%X~�]8�,���]��ӝMI�������x���� ��MK�M�ε ����½P�WFNqCg�D�煿@��F
���o�&?>�Z�4KJ�N�4Ձ�h'�FI28�/Ě,��#H8�$9�1ML:����&v"�dW�D+aA1z�B"�\�R�ϐj����\���b���_	K���x5�H�A@ܠ2�a�Ep���Pଆ)	bM�Y��|l����$�� r���@��?]�1S720(��?��5�s��i{�������i��}�=��Ͽo?���I>:����?��&�i��2$����%�����R1��	�6%|`��M�q6�P<ƍ�ښ�t��d����O��专�_�_@��J�H!DBD4d(m�uL Hڧ+�v"��d����=��^wh'�S|YW)�a�ps�f� V�UBo���־���J�'���A�4�N��~���bI�^�!XYm:G-^�np+�����E� ��&�G��,Q�4�e�dM>/<_Q#�q1ɒa@ب�1f�K;e����nuX��,��#�0��0'��`�bH����&�E��
���u��(0���h��c�Ǘ���	>��򬲁d�ǲ:�/���5�Ϛϐ�D�+v�{�Wv5�~������!;�C�֭ �,pY(߁����,����`��<d{�.�!�s+�B�dUg�`B�o�_�$N=c�[Pz���A%�A`a�E��Ų:p�p�D��!�aGI�2R3��q���-w��S����H>l:���L��	:��0؎��4hlD%������tn��.��N��&g�,͇�Ź�x^�#
�#�U5H��lF�*�\�:_��h�����#`_y��GɌO���x(#��5,=�[sGL��yy}uk���@�%��	��a���p"�ݸ������+�y������G����	���t�QĐ�J"F��&]b0���t�F=��Qn�=t�I>��g���Z�4��[���{�&�C")5���˺��"to��� �>��{�WM=���xrВb��	O���ѳ��蠜,~�9Pd+�e����s�Hx��[�
^�?o�g"R�1Brq��火���n]�mr�}Ӡ��:Lv����J(�)�8b�YӠ�����	�)i)P-�x���0Mh~S��qEzdp� 蓀m���6�hn��%@Ecm��P߲�)P[Yퟦ��48�����T�p܎��w��A�?��O+=��[��Ы�k��^��Eވ���'�?M�w6|�G)!����/�DF3,ݻ��hq{�QC7�9���)4;������χ��۠��+�u��O�������Q�ז��h��Q\��_�X��h �;��б�6x|��;��p ��?ݷ�G��#�U����$�Sƻ�|�I����&N���S�(2�q2� @QeQ^]D�k�E} ����	�W��2ma���nW��	�G�n�'�~?�Ǳs����<џ�7��O�B3)2��N	�5A�qb_j|�.R��c&�gA�)z,���&�R�+[��>.8e�'�(%�#��Q�M^��#4�@��_�z��S"pU����t��t���A�D�������N�3�_�8xV�7YJ�=�s�ֱ�d���w4�?,�5�r�1r�[}�����	e\$:�9��ף�36.
Q��q�4y�Y��	I�+����/C����H�;�k�����D�	*��&I�����=���*F������v��^��j��R00�������n��<��pEl3)!NA��F�;њs���ʒ�/���p.��Ɨ�C\�\v�Y�c'�>�%�+)s3�;Y��gE���î�"FWھ?��,��cgK*q�r�'#O����������F�W�k���
��.a�Z<���;$�Q�Jf�WEٽ*�h�]d��^�>p,<2�rش�4�|������9W�}?�;Kr[���dr-
54Ei玉�O/�{ecu�}$���wa,��N�mMu�:��Ip�Q���_��o�a�*��/ �?&��z3T���?��t�Ȳ�S�Z�r����ϛiB�/@Ѹ(��h�#� te,+(��AY!|.��Kђc;"��נ���׆�߹�R�{��t��#+�8X��c�YjS��׌��9���:��5.�G���y�0��}��1B8<�s�(����҈�C�_8p�;Cen��fZ�k��&�n��*u�fԣ�-L�V�8�rZ�\KI��j�����ֽC��8Ś���j_�!�^�J���63��GH��b$q��ə�@����G~�>���"��zb: �ÿ����x��f(�v��xTB��>�� P:�Q���;��楂ݨ��Jl;Ú��M5\iw�H�PTl)���4qNo������'��&ua"������O�1�4����W�R�{$��z3��Zc{$��;UByC����_�Z�^�!R��HKi���a�8}Ѽg��isS�O�=�;�����\�fw���+5c!\w�F��,chىh3��Ɵ$��+���#��V��N�9Yt3рh!�k��R��� bг���Y�qM��M���[K<.�'m�BZ:���>�`D� >2��H�[V�Mլ��	Q!�]gE$^W���V����7W}И&�#A���T!��צE�5 �8�m9�pF�K7�nm�}?�U�T�Y"k��0Ev���V��;P�Oy�xl�=~�'I�eW6�E+�@�kp��� 5�<�?��"q�~�/�p��LY�8���a�y��!^ji�!����>q����D!�T�P-Cz��Hד�¾=y�1���;�.�`��e4�ğ�A��gZk����M��K��oM�(<i�U�( pJ��[�<r=��$QeCu �Ac��\�W8��i�{jjj���D�L���Q!.6���H)�~���6bq��E���\,|�#�!��ґ�F�^F��j*p`���L�M�N��J����!�|�U>��G�?Z,�u@t�?{�,(���ꗘ��w��&����
Y	��i�O3���������<n���s�����Cae+Az�l'r���(�qDuW�eQ��N<���f�~޿E?��Wь���Zp��0b��V+��1 )%���������Z]��.�eI�|�2XlX��߇�Qt�x���8Y�� dG���DN("J����l�R���@�VE豬H���+F{��� ����{K��,)-��q�h�V+477C^^^��s��U4-���a����F=������?ڣ�;k�IPX[c�PLaM���lHg��&���u�_C
B6�$3w:�?�i����3�����B�dG%���V7ќ|t+kr�̡ཌྷ��$
���%d1���@G�������>��l4h�X�!�}��v0�D33v3c��h�����w�DäkR�R>�q5e#F�A����r�r��-#^����so�/����I�j�@R*�3hLmST�z|�s������O��p)�.� ���;��]�u_�n0�$&|��0ۚ� E}#Nɢ"�h�|�)/���\}���x�RRt�f������x��F����������zgL�X�>���&A�,y����~� Uop0�`�-o�����d�7O���)����lE�"�u��>�t�zm�pO����d�}��B�+K,��D%�qg�;�D��Mu0/>ŇX<:A�DJV�2�᪖}��^`�GUO�������6�5�o(���dUD����o�:@i?$��EVO���T�S�6=��RA�{���	�f�ϩ��XO�m@8#ܥ�7Tz���.���(16'p=��~]_��eɦ�+caV���ld���Z$ưZ�w��m~�,/ k\X�P��6��hK�v	)U�
a��תD$�~� 3TGsj;�/8v����e!���vl�/
�Lټ����|ދ��7���J[7$	��|�e�G]P�_�	�e&��M 7^C��g[n��GS�,���>Z�#2���N�C�(F��U[��W���ZE�ar��U�b����͋�J���HEJ��[�#������K!r�,�yG31{8��n1���w�_�+49��9b.��	q�����z:�Z$����q�i��,�Ӻp3�9�)fO<�꒮�\��]��P�0|mVu�^V(�(9 ��\�����C���-������BjzZ�*>�@�F��s���|"'���
�����́�hi@���jeti,e�}��������FmC_����				PYYɿG
�P�dРA`Z�+](z� tQ��ZH��B3�59�}��>əPUUŉ����z�����п^d��-��� *��2��D�$��P�O:�<7�-�x���ƗF���CEy�; i(���%P���zp����^qL���o��C#�2�%
Z,��g�^f�5��kFD�Dv���]����lXͨ�o>�T�q\�qr�$��|�!�u�PU_ó��$�Y�x�7>S@ԇ�Q!_�y��L�d䎚,�Ů�@�.h�H3�$�tN����fbY}T�����w`G��4X������4i�9�&����9:Q�>)u�9��7�������!Ȱ&��P7����q��[�-ű(���v:[p �]XW�m�
*Ø�*_����;�*�Ѕ\��9ݚ7�e�;���,-'kfp34&��F����NEYo��g:#z��e��XQ��E`��	i��lk���)���~ˢ�N����D"�\v��&p�+�Ԗv]a~�=�Ó�K��#�]U��<9qG8|Y���ͮ��
�V|;��B�,��jɥŲȃ�eڶG{�H�x5�����:� �/�E�Úo��Q}��~Z�W���W&	��"o�~Q8�^I�j�N3תŲ֑>N�4���%{A'�h@sOR6�)� b��Q�aM�7���_��^���*��m<� @1u��i����}�"g��|K��g�h�ꄻT��ʛ������M��j���)-� ?��$��.���,H�#d[�l��ۯ�s*�i��W�kmŚ�g�@�����@������p��h���߼�M�����L�3�h��벪^ *�E�(^����*�A_$��H�5�uPJK���~4S�\	�8��i_)W{����A��9R�3*T}a��y���N<�V�Lk�d�0��1��bF�z�|��׭�VkyY��e1p�]�t9[^���C �n:�B�ڗ��d�d���z��a ��x���3`|�`ȩ9���m��x�Oܔ�	��CA��@����I��ՠ�܁��cP����Tmo��6~�	$)C�)Lh�P��
V�W�>�����Bx?�#�,��ƒ�~@K���>o���d�WR�6��b!"��8z����êO���
�A�� �͝��S,Z&uW�PP�jk��Y/kӱ4ge@�M��6�^qj�� S�|Jն���B[{h�!"�o��NZ'��a��O�Ao������9B��Y�p��&kV$c��)0ޔ��*��F�z��i�X�t���\���W ����Z�G;A��'_I�X��ʏy ~��F�RSz�i������:8'C��I�,0����c�an|J��5�����ʄg��r=�3	i����x|�(K�%oT�T������Ñ� �	�(�k}���"a�8r��_`�޵�0KQu)U�����N�M�ߥ�� |�?w��~)���DK�L�.%���T��&A�.p�����c�*�7�LL�q'rIg�$�$�^��Ce�<�VD4n*&��s���(���-|ݛ(T��}�r��w���1�ť���k���A��$����x�E�F*W父�-*�Д�Yj�v蕀��֛R�W���z��\�hrۏ��Ҷ]M��iP�d03��ZE�,7XkUH�5vTR�HH�O�eMs�J6,K��}5��3-K�]�\���@��'=�9��53�����ǧ T����Z,�p�b0^�,��͞=�[��ZZA:�9#N�����o�ȿ<=�&R,k�K��!�����%:<ͫ��d�Ɍ,/�����?��Hj�[pI�S>r�}߾ڪ
�?t�Q^��
n3�o���f���x��"�����3�rU���v������F}���(� kNIfM�
W#�x�G^�&%"©ԑ=Q�#Í=�)���#��"�P������3P|��/iu/t���'�$}�u�9E�<~��c�C"�ߵ��l���M����*_b� nKg�w�=�{����1m�I:��yYv-�xQRD�to��B+��w�e9Ƕ�� ��{�lWڼ��f{��6ӱ#xd�}�,A�4���	�S�	^(˷N���s.u��@e��1p��S��� /�,��Ei�� ���?�	��H��B��'H��Y���A~B�{CM>l�/�y��c�]z'4fD	"�͂o�Bz��C\`0�32�Y���s��k1�!R߯)W�)*��[Y����Q$RRb�u�� N��T!lUR����2�=f����,	itU�x�X�ɼFth�H�H���qԠr�7�B�h 2,G\�A�t��oEX"��Y�Id�z�"/51aa�m�ԫ*sЉ)��M�?���G��&"
-��_L����O�D�*�����z�%��mܪ�[�(}&5Se߇Ĳ6"�J)�\}���u� H�Q(�e��z��i������/ ��"¥�q9S��_B�����FtJ%��ԙ�:ѩ(Ih���\XN;���tgI�r�"z ��k�����8D\~�G{�L�p���kaF� �H��f&�6D��Dq�r!ʻQ�]!�>@"WUW�ּ���A��/����v�c�h۾N�O�nF�Dفz�r�!t3��mޖ�T����Ak����s��q����`dЬ�H+!;	�@��R��!9��������Q>�8�HY7Wi<<T?b:���o���	DI�V%o�_?�8Ύx\�$��W��	gզ�(z@Z�u�T�M���
�m����>}औL�gn(�-�(V%(���9t���D\vJϤ��n2 Gg�j[=ז���!<����%X�`d� ȯ*��Gg_�7~n�w��$�����u��Ⱥ/�E���$��u$�b�ŭ?���90{�$8��D(���K����F��XT�֗�[<Ӊ�E�Y;p3\cתQu%� Jg o��0A]V
�I=ȸ�`�cR�Hi�ym�������[�����Ǟߕ����'�m��!����M0�2�Z8,Ԁ�t��g�����J0���Y��/JCi��,�� `4@������pZ�KƉ<Qc�_�Ѯ@�P�&z��I�Y��!ǰ7]�t��U�C�-f/�ߞ���}�{�W�@����7->���xE�5kւ���9�p��>ْUc��22	<診���.�h�����0Y0�$NKN��x�阗��hթy"���I�]�$�'�En��X*�JLL�~������#�_�Q�((/��c�B�lB� RS`��q��Tղ��I!�n���7(o�^JC�A/�Fb/����Sx4BU�>�<6%ů�lN��\�r{�0Xok���r���i���57�s��I�����[��g���E��L+��XW�~�2b:T֖�Z�ڈAbHF�6	u�����;i�}�x(u��K�?�ha�5�B��
_�o��5y����f�p^������ږ��bY���k�렬����(�H!�DE�/�����4+
����m��B��6T���^�R�޶j!';%,L�����p.O�얍�X�r��ؖ�rm��(aSs!��Vr�A��2�U����lv�� ��L�~�$-�����,�4D�e��g`GCs�+�˰#��%N~����!
�|~�����L8�/�u^.�d����#�7����]h��(�=D��Vm�V�����ے�Z��/?E�`�!�X�#c m.��GLц`��#�<,��(��r~�⻑r�ZNB�OU��{��0Û}uAR�Ϻ
�>G�GK��Hɑ�v�� a�	D!iۑ�7�qG�X�Ze�E7�e�U!1�F�6��Q�ۓ%�[R"����xP�d-#ٚn���(C2^���8��Sa���P�TFd�ԸDx����2x5k�l�0	׽@r�r��Ғ qG�ŏ�K�N+��<䒵��b�����������H*5�JzB�쳠A� � lF3��6�_�S�L�g�}e�� �o9�:�o(�L�P��@���A���� Q֘�o���;�ċ��C��@����#�q���8q�y"ݎ���ZZ��m0�"�k	#D��{���1��� ���� �1	��-�q��m��������Й��%�����{�RM�"7%��<���j^�!9!ds|����8��&Z�3�BU���"�0f�Z@�ά#��nH�w�҈~�6I2\�o:*��h�#���dS���ǡ��C��ʦ�2���!l)ʁD45�>���3zee_�Z4��A�dn�c�C^�=�&<9���
Vs`�V���P�:ѧ�&���h��k!��z{���a��Ŀ�O�.5��bY�k�S>j��S�(>�j��6��^\W/Ք���8Mj]˝̞�%��AN�z�<�+�PS[
Yæ�6~�5��n� ^h@o�5�7�ldK�:@�`oh�)�?�ᆑ_F��T�m��q�HJ�!
�����*�[S ���:�d��![=8z�o��R�{�ύ��5�Gx��N[�{�#�$Р��Z,+j�\4��t���a���Є>�+�I����~�s7�p��S�Jk���À����~�=%��t{�.4Kr���qr8_�z�8L�0�d3�䘬�����!�h��g_��/�i�
Б�SQb���k!=d
��K�8%_rֲә�
���I�|$�%���B4wq�k0���q�`���6-���7]y`;��%@ay!<���S�����j��w[I.l����-�F�N��p���!�[vt���$��#�?f$I"~$^}�ǡ��:>��N3���~m���jQaoDT�*���b��q�p��Oj��Ъ;�
�X��0Ā񂨥��j'������,Y�����H1az\��զ��e�+&��@-H�k��a���/xp�Lk��W�+q;���%�ǲ�	d���q	�d;q�_T�.��4�(����a�@bd�b���TL� �� :�$�j�-��EJ���}��ы|.�|=������9$&�`Z|Qr��i�)�a4�<���|�"�em*���wah�{��&x�/!^�	B@=�N��Ę���0⎈���� 9ā��d��� ���GU�l�{^*B�������fz�q|��Fƶ��:�d�*��2��k�� 	�[f_�'^���[g-�7�-��##��h��(��[�vt��嗾�1:s]�3�Ųތ%���0S�V��J��j�ݭ�����f�h/x@�Z�АB�SDb�(H����zO��Y�i�����+�Q}r%�]�L���\nXbL�@>�_��8Fp:ܜPԖ8�KA�1�W� �3�]
�#.2Y����b�SI�3%�6��#QD����_
��C�,l|�jt��촃�__�\ҹpŤ�|:uKQ.�;���'�@�N:ÇD�XL\d:bb����8�d6p}C���AXp�{��S�g��3n�?��g��kR��+2�c ld��uv�:u4����~O����~��
-L��D��ZXE���(tJk�់_�,+U��u����P4��C<��'� ��8�5� 11������>�lX��b��\|>����'��p��"�_�8#��������D�e!�@��-}�q�<o)L�w:@�捶O@�G�[�����T\���!��;�9T��g�l���-&�^�kDh��
&h<0�ɆX0�{�G��5|*���Q�X�o����E*w}z�l4�I�'��R4��g� ��	eu�]n`LdC�E�)K�����ne����22Y�o���(̐�f.�U�oc��@I�r!Jc��ѫE-`�ʺu�\�����ҽ�!3!�ω�uQ�@����!���"�n�:1j��脢�ta��e� 2Qg1͂��p@���w�$i��z��R�A�%^\�Mp��+`����ܲO�ˁ��("H\9Њ"L�m���r����p�BD"�ߥa���~�h�����G��}�Jhvt����ˊV�'R2 M�o][6^Z�	��[�T���Q�YQ4�)hH[b�@���(�z��1����J�p�t�zq4;q  �/�9*�7B3�fbќa5�+��yY�$#;=I�*iP"~'Χ:[�`�[4*���zVc��W�+�v��N
�������oF.p3�]MF)PƜ�	�}u�?T�lW^ }�B����E�:_�}�C7`rl$�_ş��z�c1>�&��^��>&��\��4�=7>%�bY�WX�h�ѧ�3D0y�>c7c�Ez�r""��ڿL���������4����@M�l�^=�
�?_d��}�0�y,���\��(�Zx��$H�����.���E�c��6*�6�ٗ��hY|qr�Wå�#���}I�6��yy��Ě>hL1[�������s���ُ2�K�w�<\t�xLK���%�H\Lu����ט�δq�����τRڟMD��p}��{A�(ՠ+q*:���8���v��o?"=�q�̋*���mS�K,70a��Z�ƫ*��7ZfX��~�lcm����-@��������ִ�#���ΊK�2�a��Q����ƴ'ӱ��G(y�Ũ��*\�wm�[�͂��}	e���a��X@F'�?U�F��pj��2_�˝o�U-���y���i3P�� j!dMB���"$B�E��� b���x���6@bR:\5�t����)���(��n�_�׋Re)��N	b'���*D�{M�4�^w�/���c��'�����̈o��f[C���o�����#Qƃ��S��ޕ{Yk���~�:��ǎ���(G⨟�o:6��Ecu�xM�����D&�}A�K��t��8��9UO��+m��f����RF�Yl�Y�Q�p�Zp��������w���w�D!��.K�s?>�JdnC�ވo?%��	i���Gh���k�o�߸����?��o�<WK{� �O5����l��@Z�;�yH�G )k�ь��B�Z����uB�d��9���m������F����;�$W��v���U�`M*7��u�1p4>�pg`,�k�s��a�Ixx1_cx����e�f��ݎH#o�<o��^:��K�{oYTR��c�Q�{]���_�A$�9�E0����@h������-�v��c�>��,A����
b[r�1����	R��J�/�^��?�9���RT�F��E�J�J'&�����c>9 ^���H�u�|�&�d_k.��<o�Q����)ZҠ�����h�����X�� "@�4���hL�lg��I��*�O�\��i�;�s���\w��n M���^��>?.�s�V�+�':�_m����I�(��;�?C��ޞ����9��`,���a�Q�G.)m>��X ����u��Vŷ�Z�l}��ߙ�M���H����F�(�5U2�	im�R�e�q6�[���x�
p��O��e��,�4�K����i���mus�,(~�/�B����]�o�&t�Z"�e1zc"H����Br��anCS�yxa�B�#�b����ke�E���d}�q*���[[��uK�c-���M\��K&tw���l0­�`�)��Y��tm���
�R��;��(���{�ιdU�򶌁_�RY4h�9v���}&�QY���8�2��yW��%h�ъ*w$��@m��	B�-G )�1w�Vb4@��pg��[p[ڀ�׫�/D��&�F��<s�n���%�����+���[دeFA����B��_���l�y�M,�@��Ef���9ẹW�)C���:�yR��������p��#�?�8.|���r�����2�����]�R��1�.	QWkN���ݺ.͠�hr8%���@U	�?n&Kφ�YC`���G7A�_���U��8$\J����F��Z$�#�Dj%l{�A`�ă��'7˾�D-�u�Ą���@a;r��MPgo���WV����ˢ{ g���2D�V��@�E�����YPe�)+�_��"���w��Ef+m���C�x�;
��=g��ν�9@��,��<-.�}#�Q��͖̀��j��\��J7�4��_UAk�@�b /z�1&�ڏy��т�R���w-�ڛ�8^@bka������B�/m%��ɤ
4ދ��D4�<������'_ k�w@>rȩcO���P�uG:i+PU> �d��+�r���~�!������F��
�z��?O��fW%�Nw*����h��'͇��)0w�xo�w�|!�	2V�E�s$.��R���8����K8���.�e��C&�9cN���#��m�awI���#d!".�	5�\dUWBIsJ�.X9���R;`{��i��wۗk� 9n0����	�����"�҃��>�S��x� M��O�/I�OCGp�_c8N�X�59���@[�@���B��t--C�KH	L�c;�q�<�Ar�s�󠲹�+��hr��7C��w��N~ބ�$*F��.h�1�<�X+��Maa"Dx��MA=cn�� �iC�%���Π$����G�ʗW}%�e��0�3%�Y���q8eb{\��`b"\�:-�>��]أZ�]߶Q;�bM�R�"��e���tދs�SU>51aRw!��#�<_xю���*��=@H��z���[v�y(e.w�J�E�@C�?x���F}���yP�aB-��Fֺ����(/�(��(���]�����o�}!ħ2��mR/~EJ�p(�E�� 	@;�I��M�V�P+�{�Y�螙�c-/�1*O(�>|"��z8D��n���A����I*��?n�g� �!�T�֊b�L�FN�f��F#w<A�r�`�KQ���:NUكa�N�53/��5h�ȋ+?���C]��������}��~B�$AJB"�x�\x}��=�� �������Y�t:N��WQ�̌�d�⤭����C@���8m �O��J|R��0w�d�Xǁ�z�YY�&��!�g��I]��A˥c�4�<��}$U��6䭚C��m�5�b�[*���cY-��`f���R�����rz�8�*=9M�!i}ᥕ�w���BYC,C3�vD�?wX|�.�q\������U� ��v�m,_[�.I*Vdu�˦/hߵo��^�U�6��,�Ԭ�=O�xϫU/���J;�
,���.�@���cm�%D��-x�@�W��?D���'!�~t������B�e���xQD�Kʀ?Ͻb���H���x8^�e�sf|
�m楰�� ޤ��y�2b�,=�B��a��̱	-��[���a/���1�u�ׇ��
H�����cf��"���>�����ᲃ��Z��?��jri�h��D^�=Yз`)f�ΖL!�L�;5�RJ��hf�֔�3̎��q�|���?�)���P�[��p�:��FnR���'�5�[�D4�Q�]����XU� ��|bؖ���l�2ڨ�'�9�,����dUy����S��GN�I͑��
3�N�kBN5�#����Y�k��'>�5*p�����	 e���>��x!�f�a�C����>��uhH=A����gNY~ �,V�S�{D&��g��=��{Ρ�N�xT��11�W)�U�S�y�K��a�A��,���O�����o O����p����'	��11�9���ʹ]+�H�{L�P����6�A�Q���<�B&)��`�d���iQ�n�K��)9�w�}��A�^6�S�y�O/��&-��`�[U������F&<�㰵M���H��#�@yS-�P�p�e�������[����K�B�%�p7?!�A�*�E��C�^�"k^P�x	��NE~P�2!����&��؋����/���� ~E���7*��N>�d�z�����_�Ob�u�E �VB�v`�z��Tz���
��$�%J��1���F�5��n����ūPd�/}�sǕ�Ws�7AH��DzU#'��bCR��;����#`���P�h������l�y_(O���J1*�l��ʋ�Ж�Q%���1Q2$��t�&w��'��~�
(L�@�(�gr+�xEk����z�̻^]MS�AV�����@�����e��M�/��;��6t�px�^7����ᮀ�jDvU��ǲ�ر<G��������B�,���x~r�6��/i���}���#��_c�$���C�Ĳ�
1��*[�k��p�у���AD����!�X�ǲ�"S̱�� ��	Mְe����2M��e%H ]h0),c�Ж;�>�xUŸ��ז�t����'��+J:��U�Y0)6�������[���RՉ������rE��m���ώOyݦ�_Ҵl(� �)��X������Nsga��L�o+�:���%_��s�K�3v���=�O� �a�K�o��.t'~���_��ɪ��WQ����p��&0q/�SU��-���L�>ź������mˍ#��'g��SN��J�P���M[�r"�/�cL<O��~�+Bs��T6T����z��oB*_�e����>E8�r*��C5}'�n$�����2M�c����NE��O�ͻ`���m���$�Ped ��TcV[O���z�D[3���`#�~{�y��Ew@.��w{~��w��x�:�"�©g��*i�b�5	b���
�3��;Uᦝߞ[�	,ܶ|nW�؟y�O��.���>����L��+Oy�7�BaM_���.���!���ֲ�3v�<��y5��j楬X���M�c���($�ϵEYh�0� ����p�	'���x*�k�+��w���|J;"	��Ms.���^'d���|��G���AA�H����0 %������]p\�������|�g�h��w���C����6��=�`g��-/#"�Wډt��SyA�/�:�:xc�bx�珺ŷ!��fYS��V|��3H�.G"��w����!)U��CPF����#i9�fˢ���OD ��?�TZ�$j{��Zu�#�,$g�#F�W��W�)g��z�z�rD���v��[�~(ή�r���`�swp]t��I����^r���c�jT!������"�Q��|�F�n�]�d5���"�(o�M��[-�i�ϓ^�"@�e�FJ��T&�҄|��VN�O���������IK*y��a2C�3Y���N+���j��&��\�*$!����`=��i�N�1�\�E����1���$��КuUi���gH\���^�������W�Hs�%Y2�k���i�']�)��<�� �ƒ�XV�����B�Q������3�JQ2�,��!�HE��>��g��5���qk�hi�#���Ӈ��W���s���-�0�^����
3FNF}d���gU�"1�y��Ho�)w� �u4A�(*��*,�.����Ew�D����������@���4��S�5$pYV��h�U�٣g���KQ7,߻>�m_�Pq���;u�/-���]2�,���^����Z�D^k�V�&}��F3t+D�e�]��\��ˋ|��yT�E�G�����[�t�<x�y)�<�C���z�O�ˡ]�ӯA�̓�-yʩ@M��LB�Y����Q�]ۑ#��-p:�5��=�`T'r(�7��P�	VJr ���X���4�5��\�B���Z�#�0��K�L&�\<�TxEQ z�+f��E����K��_�����8N?a�̓g\�hg���̼���EXG˳I�g�#G�Zᦓ/������F���kMJ��lF�n�Bi3�m��(
��֏+^�?�uԲ�q��8�� �CD���Cq�
Q�?��_(����YȈo��&�����J��W�2��F�y�{2�4x,���]�uh�]�������*��bY�3�RTtj���-�4�R��d�)�n��q�����[�;��hӠ�ڇ>í?	�]� ,��_p���hկy�v�p	m�l�D���,�"/���F���'΅Oo�'<��˰6ok��r���⒨���C!�pg�~WO���b(��<�y+VO<;1�Y��$~���C6@ef�s�:�?��m9�}��085�l}�=���GaS�^��ZX	>a�xx�ڿ��p@�x��?s�7�IL��~�%�w��E}|����_T�@8')��W���;��h��������H���(�oM-��*a�7$���j�ϝ>Pҧ�%<�Ccuۈ/W���ڷ��W��c+:L�=���ܯx����۟����MK���ԁ'��Ac��+a'�_NT�}Rx���YP,��r7ö��!���O���'.���Q�8�� #�O���X���wd^}�xW��K�ߝDm�N���Vb� W�اz7h)�TCEg(�hf\�QY�k��bR߂���_T���+Kx1�Dt�N5��R��́Ǵ(���u_���7��~N2�;�3P?�MpB� �=�ħr�po�!�D�c�R�]�3��mU�qڤ�A5A͜D"�T,{��D��ص�v�X���������?F0�]�r�ɓŇLBP� 
�Q��1/iC�OGGp��@Jl<�û���/��/w�`��5�����1��j�ZL�&{3,ݾ����͏qn����?�b�a�'/��=�	�����]�����p�aH�۩xW���?��i;Ol�JF�q��憇�Q�1���!��`������8A�*p;����B�1n&����cH�@z�kP�uGy&*�/n~�����h!�㹾�4~s��p���ܸ=uK�B�)���=��/��+�;?~l�f�i�jX���A1Hf��G����'J7� ��t�i�@�e�a���"�� �����S�R.�������9��Q`lL��]8�]����u�F��g����}l=�(��+��~{���1�#0[hO
���7����mPX~���a����mSmRJ��
��;�\U���S������}>�%m7����%>��>����IN��ɑR��g����U�Z\�XD����/�/����ޏ���H��ar�h���g�o���\�f�>	>�韐���N��@�_=��S�l�28�⌔5%�e'e��S��J�^��"(o�bb׿�4�[�\�>rEy��dhv6w��3���:o����j{Ĳ�z#���^��p,�ԩ�lB2LɄ[�� ?��]�^r7G,ͯ�����f&����p�+y�.�[䗐)�p�28�廡���-?n<�|��\���`;ꘕ�qB�Cn�E���ґ��]�Xӈ�W?�{�UGNM�6��p�ؙp"�QS�H�{	� �w�{��C�����w������z+�%y����[��(�6��6�m��@\�-3��]	/95�վiH2z>��Q!�d�62+��AK$..=��3��BQ�}�r/l"#��x�r�r����w��S��O4�z�eHL��"=��n܃&�.��3�6�h�k�aK�渓ٛ���P��a&�h�hg���hL;��;E��+����&;i^�#��kBD��J_�Z���;x=m��}��aS.�f�$z(t?��0���A�0���ݶ۬��&������y�f�ݯ¬gn�]��SE
�GL����f�.7Z��5")#��x))� �HDL
�������l��0x��?�D��X����8�H왣�����k���`h��B�Q�`��o��䓭?���M0������Ϲ�bw��89��L�K�ZA�����l|H��o!E'_�������\�W_���磈I��`ְy�E;Wv�jANJG%~'*g�����yP}ڼ<-k D��Ϫ�khS��
�VN�ہ��<j��v4 6 Qhn�4����}(�:ܵ��t:�C��oػ��b܈g�	n��w��xDB1�ȭ(�fA؊��PD��zG��׾\���[�mbgX���������QP�=��{A�uaH��#����2d<M?�l��e�����$���r�=7dHE"��9��'�K�>�K(r�g�P���rm>��2��f� ���B���d�;*B񔬪O���;��X�J遑���z3��Zc{$
"nK(o��K"���"���s"�����d|�ˏ������&+	I���"�Z���襡��qIP�w��%�0^���r��� E~���&K�����	¯Q����Fm�Ҁ�L8����pf�fR��S�-��F�{��B:�?8�o"_c�'g��_� {�c%�m%g�u�xM�A��$�����bU� �"	Ǡ(�܇�^�9�����%.�K@�k���<!.���_a.�:���hj��uɈp���Y�a�n��.pS�|�fW��%�JPD�L�5˾�uh(�Y�C½ ���zLZ���4[����ٞ$�y,+�$��i4yI�>��]�1�i��X��D��e8�U�ó�s����n�J�_��[t|5/ZWWͺ^��^4���24w)��vg���M�ͧo�ؾ�o@s�S�����9g�Dx��x���$�܀.W�*Ų�!�`:%�hډ?�������:��*���{o����WX$	VIT$VE��V0��kx�OYWAE�
��	3�r�!͐&�t�����힞��a�}�������U�:��9UNm�zmq��!Z��מ��W�X�V�y}w��-���J�%����҈n���?�ǧU5Ț�CۃZ��@����4�ۃwr��'�H��j5�.V�����J˙=��mRB
���X�p�i�p����HCs�x�-Ըn#y�?���r�e��"�y����#t�+�Q-�����7�X���k�|� �V�˪��s���^Щ�}��J<���\�/?�"���\��Ѵ�&I
~ⶡT��q59n|��/n�ﻼ��Ԑ���;
����^���gz�)(_�1�u���Nۥ?���/̥6��ҭo�55<�*�r��ך�s����8%�@�i���h��B�o��nq �sҖнzJ�ǱW�l�N�r� �-L��ǵs~����osdcQVֶ�s��zQC�5n�A6�:�e�Ay[��2_]L��;�3K�[��h%_�D�"��J��P�_��x�$�5[�5-Yf�K�!`!L�SW&=���^_>CM/~�� �_Á	�.N�<�z��u$;�3�)���,�a�l<�G����6�Fӂ��Z%#ːZ`llqHV��^�,l�r�Fy>�|���@V��n ���	�6q�<+1O#�F8�9l�&2B-~ ��c�ð�RU�-D�/+o�1��#]�̂دUahP7kV[��a7����-.�-`a�>��9A�@��j��()Р�ff���Ec��:_ۆo�6�x �j2D��*3�PEv���e��4�BG�[�@c��6�!䊥:F�������$C�L��U��t�DJ�X|U��;F��+�Y\���B�q#�Ζ�LJ�@ʒm��m�=�޺/�8#-R  <���c�*5vN�����X1�V䆊K�4$��̫ߣ�A��r�S���0�}��o�>>� 7 !�*�6�A;A��@L�+Qްc�\FSM�}G�h@�[H��ւ����$;个%�ޠ�s�J ��Z �0����KӇM�m��#R*��ߓw�� ������0/���[�<��T���HL�_hO(Y������*��NE��,��;�z݃���^��b�
�����P-�����`�{N�7W}
u����h�����s ���A��ؐ�<�#y��[�C���=���@�&&jE�0�P�_��(�3s
�^~�I�w��U�g��#�8=���缞eum�_��vVp0¡(�5���ڏ��Z��V���m��)�b[�O�0�xi���a��פ.;���e3�YjC)��=�MX�O�|t��[���������kgJ�����Dȣ<+5"6.���;��>p<��g��5BFWuO�#�� !��q�.v�6FFv}����0Ya����n�L���z��{0��;~ܡg|�m��^g�����$��-;J��U�y_LY���I()�1>�7�yz��8il�<G���`�rF.�zpcV�d�:�;8��٤��]�77m'���&�O�PF�'�f���L��8~x��bԂ�ߨ9%c�r}��]�n�*��CF���z��*�&�	�#�l�V���1ӵ"ݿ6VQ����)?��T���ke�f9�2��*�������~W�>������
ĳШ82��z�V��p�|�J=�5*a�(s��X����h͎t�E���<���r�s��+��Yf�v;UGu[,��B@ۨ���h,��*�=�vE�N�L�f�]ɺ涬��N��{��W����Vf�P�����c�x�ڕψ�]�Z�3xx�d����˺z5�1��J��F��D�u ��oL���� ���%\CR0��[���ƶƤ%�h��4SI��0Z�:Y�Fe[�?F�Ι�ZK�Le�Xx)pt�^�V�ӣ�=E��=�^��_f"�U�K��y�����LD�W� %�,h���?|����m��h���s��s������N�7�%���5_�|v7gu]��5��OӰ[��彄'�@B%�ʍ9-b�]�q(LC�ܯ��%�a!�*�/Cj��^o��^�0|��Y`W�資�&eրv��c��KcO{	�w�-m�~b�[P�KL�J��ʠ7�`�*�T����/�#U��������Nҭ�:˿�r��:����٠�;��8��6���ޘ��/n�*���}���I�J��5��^ӂ��&)^/=е�<}�Q���<g�s������W~J3ҿ��CE� F�	�|�!?�v���h��҂`�XT��	�ٍr���v����/�A�����+˔��هaD�C�fH��D�C{T��ٜ҆�S��Uf�|cU� Զ�]م�*"E�� [�����]c�]T��{+!��6 �c\2�#5^0+/���T� -^��f�3 � l�t��z6��9cǨ���aH�7�|2,3�~�e��O�qX��F�Jb68Q��|�5�̎lH�����^��?;�o���	����/t�"�(��.�#1��ͅ�ޯ�݅��k���p�����4`��KQ��-�n:�����Z��Q����V���@{)/����6���N����rK�/�(S�ŊQs!.�B�"���8�=��T�<�Zպr�S vL�X'�� $Ef7Ya�3���ѹP�A�.�h���z�ə4g�c���y���(3���q:����	:����K*�;��-L��2`�2�U�~6'�j�<k�+2؁ca�E@0,��:�Qv��J��뗝�Ȉ�	����&�~���S��\WA�b"&��f�Z6���?3g��o��f�5!����T�'��p���E�����v�]���f+�N�5{�����0�x�&v-��K�������F�o���[bH>VG��6n)�����;�X<t�2�������F!��d�;AC:���k���Ky��A�t�L��^Gϟ��|�M�m̭�4��j]�Gv��.�����v'MM����2"�`ưkhw���#B�kF/�qh7M����P>���(��1��eq�{�,�mzi��<jU�'w	��g�ejj��K3�z�+7=�0�rEX�c���p��u3d禯�k��f'Sؠ�s4
�ز[����[�V\���M�k����.r�_PY����?4���u��)X�{m-?�Ы�__J��'�ve�*"���%�4�t&u�O霢�:�T��9��?H[�u��7�2�2�$����7#s�1&����_q��x1~�Bԯ���yt��I�V�9 'K���cE�#V^z�pХ���=O��Ri�Ayv͗��g3�<�I�M�q��8����S���Q�6n�˭������s83`�z��C����d:��V$6̉	�swV�EV��"�F���^�~�Ըv2t�������.|bS�T�1|S^X��n�Х���хo+q��|���~xGl���۳Q�:�dp6˄�K�$r�� ��{6��-n���l<~>[:��Ә~����+�	=��\� �2�����4�ګ)F[�n
^��`ˍS���K��j���G�������C0i�Dƒy1C�P��#�t��+V�ڌ5x^�ݟo.���c(�DD�# �g��-�4�T��r��,�eF�/�n���g��A� 9��3���^U��:�p�MŦ�H����cl�)ݚ2^Y�w;V�s�{�8�a�����K[��MA_������40¾-<���;���'�sx{hԆ����]]h]N�8��/6���6o��S�F^Z��Y��0 �29��#Y%�*�MeH���#��N�y��JN�� �^���v���a3z��I�ɖ���ed�&��Hw|dd��|�m]�T��&ޥ��=������ϳ�7����Ұ�Oq"����>Z�7�K��RO�ߑ'���썪�ǐ�R}&�9x�)Z�	,���-cos���T7��������[	�H���*��M8�e�9E�5M#V��W��˒�s�?�����S�����N'=ک����8�,c%0�B��r�x�9��(��s�`��5�q��Iu�� p��>"��_�5/���;�&Q���%���a�U��,�O2�\�h}�v�kNu㥥��I�͈���b�3�V��P9QW'��P�
{�(쒔�>|�:����c��<��q�*Q6�3J�-nw(�[x��M�v�L��#K�6�w�w�������3PG�6��qIg��1_%���{�m�W��Y(py���,�}	H�ß9c4�$���X0�20�ݝ\��ŷy�9]�؜�̀�i�M�\�|_?�i�gY���%���qΩ��X���]���p�ЙB�<��P�ImL6EYv��3ߴ����"9�#�1�T���8%���2ݺ~>ˉ1S�f�I�3f{Q~�g�t�F��b�[P����C ���|�ka'p�R�y|���J�S
��,�t�X�nO�]	X�����J zG���Y�9�V�Y)��yt}$���B6`į*Dޛ5�c���,��V(�wx�Z ޾���r��ssc�vU*֦O`-O`]F��������3��xԆc��(��a8��e�	`�!�`�}���ƪ�w�� R:&x>�}�dp�oʊ$U�a�A_x�w���0���J3`_��$���%���댦���;	�� '�E�=蠽g��gp�'�feyK7�x��G!c�S(�d�n��z*,��4Q����EQq�˰H\�J��K>����,<��>ʷ�Ernk�ة/�&� W1w����<��usc�_��$�J�D�k����I��aR�a�׮&q�4+�\"���F�AB$��A<h. ����
�euvz}V�RT;a�L�r�,�8 /^^㢙C�I�R0%A�-��u��z��SCo� ��QI�B/�t��:��L�x�$U�ߦ
���E�7����f�M�>@�����g�d�+�ۅx�R��gV�Q�ۋ�\ԣ�G�:�.���;7��-��8}�Xt�)��$�ky������W�/���4�@��K����>��3{I���S�� Sc�SQ����F6���B�YmK����������C����!�O;�'�#t@}��0ni<m=f�f�@�B|�9���'�gz�*�-s&�q%��FQZ� /NM�?��,� ���b�[���[�@s��Ν	K���V��o�uIXTP��o �qu���N���.� �q�q����e��bwiEߊ��x��\l�u�tG*�l�}zy���_o/�ډ�媦2U� ���o���ݎ�-t3l<U����e�礱?U�ˠy�b��*�v�jq��%�HV�х<�^�1���[n��Ɖ��P߁��#�Vo��ޖ�
o����-��'ص��fsU��$�]��{�4�m)��WN~l�̋*�p�NK�8��H�
�5�ɀ�-{H�CE��֧��'>�`V�ٿ��a5��{�;�zP7���CMS8e���UZ�i�E���uA�|]����*~˸�"�A/����H��dЪr�U��K�^Ko�c���h|������G�3�����K����Рz���F�\��>���n"��`*��}N�|��*�
����|�%`���9D��Qe�F'����l�oV1�Ӣ�+R�G��e7�Q�]8}�9ߙ��0�x����nu�1�>�
��Jgs��g��<UV@՟Մz'�B�+2�+~��z�0�RQ��7١��U�&;{?QP��F0.�ժDM�[^��G9,�]�ll�k�(�ԥs!�+]XШ�����x���!���!     IEND�B`�PK   �EXϋ�+�  �J     jsons/user_defined.json�[ko7�+�>��^>�M���q���l�EPpf8� ���� (�ߗ#i�43����-1�@��s�:�\�w~�??���x�r˟KW�sW�/ƿ��^��4��Ym�棫��~kyc��N��舑�K7�w�ni�����W����r��ѕ�g�Cv�>,��=�xR�j������6L�M���l�.Ƶ9V��r�4Ae�T�H-�[)��ı�S�*���z�����օ�=� hE)@�DkK��ii���f���{���z^-Ɨ��盇i�z���W�����h��?u|�v�y��G��f^���-�_�w�e����6X�ꦡ7����Q��*^�_!��ԫɼ��X�o�/�ˍ���]���������X7�1��?:a?�m�����������料��3q�[��m�l\��nM`n`	�.xN4�*�ל�
�h*�5�\�Ž��Dسg�k�_;F<<��٦�u3����z������j��xhn���ի�!H����e�m�vқA
E��Me��p�/¶�]��M���7Ïeῲ����]�̏���^/<�w������[|t�	��d�6yu��Kɰ�r�j�P����^?�ь�YZ?�(tE�6�PԊHf*���ҙ����\���B�KE��	eN@���P�F3�����.`2����	�ќ������8��ҙ �O2��*I(Zx&2�ة�O'	B���.8g��l������^�(;��V�#Bс�{x�Oh����=>Ə����{|:?2���'��Р�_l�ր>�|b`��̨�O���C�>��q��9f=V���ɨRp��,�2K�xŌ�@aK/���giY*�����	fɅ����nykW��[.?����_���o�b���^.f3߫�/V�ЎҜT�Ή�J�
���Y�J��j�S˥�W���0�#�:g�T�I��
YN-��R�~��,7�|q�����qד�e��ڒ��f�̛�V��Sb�Q	�N>�˨��q���#���� �	�:�b^��A�#�0�A��>�)m"�=F��6D��#�}Ԁ2�I�p߇SN�DP)^z� 	3��T�vOe.KX�&�N��Il_YK~(���C�jau��-���5Ӛ������eoC�y�z�݆����CB���z�݆)sf6�v��C���lC���z�݆���s����)s&7��{b�|�0�Y��	SarC���arC��ꬁ��iw٭Κo���Vg-[���Vg���.��Y"a�C���,-�0šKqu��C����:˙ Lr�\�e��9�h��(`��%zJ��a�c��IiF2�Փ�Osc\OJ�1Lv��=i/�a�c��I[�ctOۙ���1�'m01Lx�~�M��ϻ�Gv���0�y����a��.��]���:k;���m��??8��p�yN̎g�U�$cZ'�%�'�p�Q�y	 ����9/���^�0l����q4���_�[;��F��C����k���	�SX��2� R���H�(T�YU䃯�K^I!� �(�y�I^ICJ�k��܊�����w���+m�2�Fq�7%]r�^�����]�A��ï2b��]{��MR�UL�V|���\��8�_�J�~s�p��(�3&��~Ϥ3��z�U^װ��˄��N�-��˪��y&�`�2���^V�8W���d^�
�qi?����H�^*){���m�i��'/ۢ"�%���d���O^��.�z�RZ��^sy*C�\��c��h�WX��vgv� 4"��8�s`�e��P�K�souh��� n&?q-F������}�G����{8���+Q�ޔ��4+UiS���Jv8��iPT0b������A]1�].A���8��	��yJuH��ʧ� �T�O�*u[��Sq�zm����T��JO�L	�TBH�#�=�{J� ���w	��çT��t��:�� J������p�G�l�˄��JB��ѻiCSR�o����^R��]Qz���ѫIT�\�c����EUZPm* +4���\M҅�
KI�d���E�N]IE-��h���y��F<�@b�
Hɰ\ќ�ɚ�sS���4	x��3���P/ %��g_�t�I[h�a��OQ�C���ZC���3([|�i��\^|3�of�ͬ����ʬ߼�~��֌�B�R�xI�|/O�j�s�(ͮf�yݚ6���Q��p��K�Å�����ꈒR�9�TyZ��mX�5M���\)�4�O���9�5�	nM�~
O��ޣ�6�r��wkzt���t�<b�
��_��LFw�z���s���ޘ�[K�,,)���ҼrJ�r��9��d�(����m*�Q7I��O92ᓅ��x<��_��s�υ�"M�2�Z��=z�d��q�1��7)�y���9Y������/`�N�Q>�����U�~�|@WV�"a�Q�����w(WQ'Me����]��*�Go��)��4G� o��8����SRVY�S=Ts�(�"�5��z�c���1�|Z�_�n]^�w�)F��5�7��ة�O.���lS�����8�� ��}q��Bo��0�ۗw/��H=�l->�OK��0pt����� �����zk��@�p�P7�n��@�p�P�Z����åB��[Ď���������j�0M��4R���@�Nc�a�$蔱7?�]�ԥ�!����������O�pB>�W��*��|��"�y��� =U�E�^��=U�'�rޞ�LR�x�H�y�$U�'����Ky)�y�$Q�'����J�DU�DJ�#�H�I��k�vy:"�ف��ܾ�GJy�L�f|��c�2����>���h��N��/7�7��/��mJ��1�؋]RȞ�����3)n�YRjW��+���e%E�9O�ncĽ1��0b�4��%U������A�BU�D�� ���h%�yd]a���N�}����PK
   �EX�&:  �n                  cirkitFile.jsonPK
   �EX ���  �  /             1:  images/23edf803-1010-42bc-b391-ef0e69fabd63.pngPK
   �EXR+`�p �y /             $K  images/29dd1623-773d-459f-838c-8b03343154c4.pngPK
   �EXo�>��q  �q  /             �� images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK
   LYEXG��<�~ H~ /             �- images/31827051-9966-4dbe-80e9-38f1832eb628.pngPK
   �EX5&�ܐ    /             �� images/3b95452a-4474-454b-80ff-b9153f229806.pngPK
   �EX+_-�$  �$  /             �� images/674f1970-5ad9-47d9-a0dc-0530c1f88674.pngPK
   �`EX4�Z�ȅ  �  /             �� images/7751e6dc-0a88-457d-995b-e2164771e840.pngPK
   �`EXv�Y�:�  �  /             �g	 images/80b57f79-5f7b-47b9-b633-c76636766127.pngPK
   �EX�ʩ��*  �*  /             3�	 images/83339b9e-8b21-457a-a82f-74d48bbc839f.pngPK
   (YEX}[֤�n  �o  /             F
 images/8a867033-535c-43c3-abf2-d13f5470b1ca.pngPK
   (YEX'�T~|  r}  /             l�
 images/8c7873d6-161f-426c-8be5-8f6703290c9a.pngPK
   �EXN�v4	� m� /             7
 images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK
   LYEX�cX�� 3� /             �� images/9e507620-50e3-4aa7-a16c-7d7ceba17d8d.pngPK
   �EXr�>�� � /             �� images/b24f041f-17b3-48b1-9f28-cb1f31b050cc.pngPK
   �EX���ɀ  �Z /             ��  images/ba250f07-c285-4988-88a0-9b0d9a82567a.pngPK
   �EX,��2ϙ �� /             �! images/d4f65665-9cd5-4bc8-bf69-d8b87beba5de.pngPK
   �EX-t:X ~r /             Þ# images/e121b57f-ec89-4d70-aa13-01e52b785a2d.pngPK
   �EX?��O�o  �o  /             J�% images/ffe61187-e64a-4024-8cee-95dd034d2257.pngPK
   �EXϋ�+�  �J               �g& jsons/user_defined.jsonPK        zs&   